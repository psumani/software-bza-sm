-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 1 2024 11:48:32

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "zimaux" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of zimaux
entity zimaux is
port (
    M_CS1 : out std_logic;
    ICE_SYSCLK : in std_logic;
    M_MOSI1 : out std_logic;
    M_DRDY1 : in std_logic;
    M_CLK2 : out std_logic;
    M_SCLK1 : out std_logic;
    M_FLT0 : out std_logic;
    M_CS3 : out std_logic;
    ICE_CHKCABLE : in std_logic;
    M_OSR1 : out std_logic;
    ICE_GPMO_1 : in std_logic;
    EIS_SYNCCLK : in std_logic;
    M_SCLK3 : out std_logic;
    M_OSR0 : out std_logic;
    M_MISO4 : in std_logic;
    M_DRDY4 : in std_logic;
    ICE_SPI_MOSI : in std_logic;
    ICE_GPMO_0 : in std_logic;
    DDS_MOSI1 : out std_logic;
    M_SCLK4 : out std_logic;
    M_MISO3 : in std_logic;
    M_CS4 : out std_logic;
    ICE_SPI_SCLK : in std_logic;
    M_MOSI4 : out std_logic;
    M_MISO2 : in std_logic;
    M_DRDY2 : in std_logic;
    M_CLK1 : out std_logic;
    ICE_SPI_MISO : out std_logic;
    ICE_GPMO_2 : in std_logic;
    ICE_GPMI_0 : out std_logic;
    TEST_LED : out std_logic;
    M_POW : out std_logic;
    M_MOSI3 : out std_logic;
    M_MISO1 : in std_logic;
    M_DRDY3 : in std_logic;
    M_DCSEL : out std_logic;
    M_START : out std_logic;
    M_MOSI2 : out std_logic;
    M_CLK3 : out std_logic;
    DDS_CS1 : out std_logic;
    M_FLT1 : out std_logic;
    DISP_COMM : out std_logic;
    DDS_MCLK1 : out std_logic;
    ICE_SPI_CE0 : in std_logic;
    M_SCLK2 : out std_logic;
    M_CS2 : out std_logic;
    M_CLK4 : out std_logic;
    DDS_SCK1 : out std_logic);
end zimaux;

-- Architecture of zimaux
-- View name is \INTERFACE\
architecture \INTERFACE\ of zimaux is

signal \N__54255\ : std_logic;
signal \N__54254\ : std_logic;
signal \N__54253\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54237\ : std_logic;
signal \N__54236\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54228\ : std_logic;
signal \N__54227\ : std_logic;
signal \N__54226\ : std_logic;
signal \N__54219\ : std_logic;
signal \N__54218\ : std_logic;
signal \N__54217\ : std_logic;
signal \N__54210\ : std_logic;
signal \N__54209\ : std_logic;
signal \N__54208\ : std_logic;
signal \N__54201\ : std_logic;
signal \N__54200\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54192\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54190\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54182\ : std_logic;
signal \N__54181\ : std_logic;
signal \N__54174\ : std_logic;
signal \N__54173\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54164\ : std_logic;
signal \N__54163\ : std_logic;
signal \N__54156\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54154\ : std_logic;
signal \N__54147\ : std_logic;
signal \N__54146\ : std_logic;
signal \N__54145\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54137\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54129\ : std_logic;
signal \N__54128\ : std_logic;
signal \N__54127\ : std_logic;
signal \N__54120\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54118\ : std_logic;
signal \N__54111\ : std_logic;
signal \N__54110\ : std_logic;
signal \N__54109\ : std_logic;
signal \N__54102\ : std_logic;
signal \N__54101\ : std_logic;
signal \N__54100\ : std_logic;
signal \N__54093\ : std_logic;
signal \N__54092\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54084\ : std_logic;
signal \N__54083\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54075\ : std_logic;
signal \N__54074\ : std_logic;
signal \N__54073\ : std_logic;
signal \N__54066\ : std_logic;
signal \N__54065\ : std_logic;
signal \N__54064\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54056\ : std_logic;
signal \N__54055\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54047\ : std_logic;
signal \N__54046\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54038\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54030\ : std_logic;
signal \N__54029\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54020\ : std_logic;
signal \N__54019\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54011\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54003\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53992\ : std_logic;
signal \N__53985\ : std_logic;
signal \N__53984\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53975\ : std_logic;
signal \N__53974\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53949\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53930\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53921\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53913\ : std_logic;
signal \N__53912\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53904\ : std_logic;
signal \N__53903\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53893\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53877\ : std_logic;
signal \N__53876\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53867\ : std_logic;
signal \N__53866\ : std_logic;
signal \N__53859\ : std_logic;
signal \N__53858\ : std_logic;
signal \N__53857\ : std_logic;
signal \N__53850\ : std_logic;
signal \N__53849\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53841\ : std_logic;
signal \N__53840\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53831\ : std_logic;
signal \N__53830\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53812\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53809\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53803\ : std_logic;
signal \N__53800\ : std_logic;
signal \N__53799\ : std_logic;
signal \N__53798\ : std_logic;
signal \N__53795\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53775\ : std_logic;
signal \N__53774\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53761\ : std_logic;
signal \N__53758\ : std_logic;
signal \N__53755\ : std_logic;
signal \N__53754\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53752\ : std_logic;
signal \N__53751\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53734\ : std_logic;
signal \N__53733\ : std_logic;
signal \N__53730\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53722\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53716\ : std_logic;
signal \N__53713\ : std_logic;
signal \N__53710\ : std_logic;
signal \N__53705\ : std_logic;
signal \N__53704\ : std_logic;
signal \N__53703\ : std_logic;
signal \N__53702\ : std_logic;
signal \N__53699\ : std_logic;
signal \N__53698\ : std_logic;
signal \N__53697\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53692\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53678\ : std_logic;
signal \N__53675\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53664\ : std_logic;
signal \N__53661\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53653\ : std_logic;
signal \N__53650\ : std_logic;
signal \N__53647\ : std_logic;
signal \N__53642\ : std_logic;
signal \N__53639\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53626\ : std_logic;
signal \N__53619\ : std_logic;
signal \N__53616\ : std_logic;
signal \N__53609\ : std_logic;
signal \N__53606\ : std_logic;
signal \N__53605\ : std_logic;
signal \N__53602\ : std_logic;
signal \N__53599\ : std_logic;
signal \N__53596\ : std_logic;
signal \N__53593\ : std_logic;
signal \N__53592\ : std_logic;
signal \N__53589\ : std_logic;
signal \N__53586\ : std_logic;
signal \N__53583\ : std_logic;
signal \N__53576\ : std_logic;
signal \N__53575\ : std_logic;
signal \N__53574\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53572\ : std_logic;
signal \N__53571\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53569\ : std_logic;
signal \N__53566\ : std_logic;
signal \N__53561\ : std_logic;
signal \N__53552\ : std_logic;
signal \N__53549\ : std_logic;
signal \N__53546\ : std_logic;
signal \N__53543\ : std_logic;
signal \N__53540\ : std_logic;
signal \N__53539\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53537\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53535\ : std_logic;
signal \N__53534\ : std_logic;
signal \N__53533\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53528\ : std_logic;
signal \N__53527\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53525\ : std_logic;
signal \N__53524\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53522\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53519\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53516\ : std_logic;
signal \N__53515\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53492\ : std_logic;
signal \N__53489\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53483\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53481\ : std_logic;
signal \N__53478\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53471\ : std_logic;
signal \N__53468\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53446\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53434\ : std_logic;
signal \N__53433\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53427\ : std_logic;
signal \N__53422\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53409\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53407\ : std_logic;
signal \N__53406\ : std_logic;
signal \N__53405\ : std_logic;
signal \N__53404\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53402\ : std_logic;
signal \N__53399\ : std_logic;
signal \N__53394\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53391\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53385\ : std_logic;
signal \N__53382\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53367\ : std_logic;
signal \N__53362\ : std_logic;
signal \N__53357\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53355\ : std_logic;
signal \N__53354\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53336\ : std_logic;
signal \N__53335\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53326\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53307\ : std_logic;
signal \N__53304\ : std_logic;
signal \N__53301\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53295\ : std_logic;
signal \N__53294\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53290\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53279\ : std_logic;
signal \N__53278\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53276\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53269\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53261\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53248\ : std_logic;
signal \N__53243\ : std_logic;
signal \N__53240\ : std_logic;
signal \N__53237\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53224\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53221\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53216\ : std_logic;
signal \N__53213\ : std_logic;
signal \N__53210\ : std_logic;
signal \N__53207\ : std_logic;
signal \N__53204\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53165\ : std_logic;
signal \N__53144\ : std_logic;
signal \N__53143\ : std_logic;
signal \N__53140\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53134\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53123\ : std_logic;
signal \N__53118\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53115\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53107\ : std_logic;
signal \N__53102\ : std_logic;
signal \N__53101\ : std_logic;
signal \N__53098\ : std_logic;
signal \N__53095\ : std_logic;
signal \N__53092\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53086\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53078\ : std_logic;
signal \N__53077\ : std_logic;
signal \N__53076\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53072\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53060\ : std_logic;
signal \N__53057\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53049\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52981\ : std_logic;
signal \N__52978\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52956\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52944\ : std_logic;
signal \N__52941\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52921\ : std_logic;
signal \N__52918\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52898\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52896\ : std_logic;
signal \N__52895\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52893\ : std_logic;
signal \N__52892\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52889\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52884\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52876\ : std_logic;
signal \N__52875\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52871\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52853\ : std_logic;
signal \N__52852\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52850\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52848\ : std_logic;
signal \N__52847\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52845\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52841\ : std_logic;
signal \N__52838\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52834\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52814\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52809\ : std_logic;
signal \N__52806\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52796\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52790\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52778\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52774\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52714\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52699\ : std_logic;
signal \N__52696\ : std_logic;
signal \N__52693\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52680\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52678\ : std_logic;
signal \N__52677\ : std_logic;
signal \N__52676\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52673\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52671\ : std_logic;
signal \N__52670\ : std_logic;
signal \N__52667\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52659\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52645\ : std_logic;
signal \N__52636\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52620\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52618\ : std_logic;
signal \N__52617\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52607\ : std_logic;
signal \N__52606\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52604\ : std_logic;
signal \N__52603\ : std_logic;
signal \N__52598\ : std_logic;
signal \N__52595\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52552\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52540\ : std_logic;
signal \N__52537\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52505\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52501\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52480\ : std_logic;
signal \N__52477\ : std_logic;
signal \N__52474\ : std_logic;
signal \N__52469\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52467\ : std_logic;
signal \N__52466\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52461\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52459\ : std_logic;
signal \N__52458\ : std_logic;
signal \N__52457\ : std_logic;
signal \N__52456\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52454\ : std_logic;
signal \N__52453\ : std_logic;
signal \N__52452\ : std_logic;
signal \N__52451\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52442\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52436\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52431\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52424\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52418\ : std_logic;
signal \N__52415\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52403\ : std_logic;
signal \N__52402\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52390\ : std_logic;
signal \N__52387\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52384\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52360\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52356\ : std_logic;
signal \N__52351\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52346\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52342\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52332\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52322\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52314\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52312\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52310\ : std_logic;
signal \N__52309\ : std_logic;
signal \N__52306\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52302\ : std_logic;
signal \N__52301\ : std_logic;
signal \N__52300\ : std_logic;
signal \N__52297\ : std_logic;
signal \N__52280\ : std_logic;
signal \N__52265\ : std_logic;
signal \N__52262\ : std_logic;
signal \N__52259\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52247\ : std_logic;
signal \N__52244\ : std_logic;
signal \N__52241\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52238\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52230\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52219\ : std_logic;
signal \N__52218\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52202\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52184\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52172\ : std_logic;
signal \N__52169\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52165\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52156\ : std_logic;
signal \N__52149\ : std_logic;
signal \N__52146\ : std_logic;
signal \N__52143\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52133\ : std_logic;
signal \N__52126\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52086\ : std_logic;
signal \N__52083\ : std_logic;
signal \N__52082\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52074\ : std_logic;
signal \N__52073\ : std_logic;
signal \N__52070\ : std_logic;
signal \N__52067\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52061\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52046\ : std_logic;
signal \N__52039\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52025\ : std_logic;
signal \N__52022\ : std_logic;
signal \N__52019\ : std_logic;
signal \N__52016\ : std_logic;
signal \N__52013\ : std_logic;
signal \N__52010\ : std_logic;
signal \N__52007\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__51996\ : std_logic;
signal \N__51991\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51964\ : std_logic;
signal \N__51953\ : std_logic;
signal \N__51932\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51922\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51917\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51913\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51898\ : std_logic;
signal \N__51897\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51884\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51879\ : std_logic;
signal \N__51876\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51869\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51863\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51854\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51851\ : std_logic;
signal \N__51848\ : std_logic;
signal \N__51845\ : std_logic;
signal \N__51844\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51841\ : std_logic;
signal \N__51838\ : std_logic;
signal \N__51835\ : std_logic;
signal \N__51830\ : std_logic;
signal \N__51829\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51822\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51808\ : std_logic;
signal \N__51805\ : std_logic;
signal \N__51802\ : std_logic;
signal \N__51797\ : std_logic;
signal \N__51794\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51779\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51771\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51769\ : std_logic;
signal \N__51768\ : std_logic;
signal \N__51767\ : std_logic;
signal \N__51766\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51749\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51739\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51737\ : std_logic;
signal \N__51734\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51719\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51683\ : std_logic;
signal \N__51680\ : std_logic;
signal \N__51679\ : std_logic;
signal \N__51676\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51664\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51658\ : std_logic;
signal \N__51655\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51625\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51599\ : std_logic;
signal \N__51594\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51569\ : std_logic;
signal \N__51566\ : std_logic;
signal \N__51561\ : std_logic;
signal \N__51558\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51512\ : std_logic;
signal \N__51509\ : std_logic;
signal \N__51508\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51485\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51461\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51436\ : std_logic;
signal \N__51433\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51404\ : std_logic;
signal \N__51401\ : std_logic;
signal \N__51398\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51390\ : std_logic;
signal \N__51385\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51379\ : std_logic;
signal \N__51376\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51359\ : std_logic;
signal \N__51354\ : std_logic;
signal \N__51351\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51340\ : std_logic;
signal \N__51335\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51319\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51316\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51314\ : std_logic;
signal \N__51313\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51311\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51308\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51305\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51302\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51292\ : std_logic;
signal \N__51291\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51289\ : std_logic;
signal \N__51288\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51280\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51278\ : std_logic;
signal \N__51277\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51275\ : std_logic;
signal \N__51274\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51271\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51266\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51263\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51260\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51256\ : std_logic;
signal \N__51255\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51253\ : std_logic;
signal \N__51252\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51250\ : std_logic;
signal \N__51249\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51247\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51243\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51240\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51237\ : std_logic;
signal \N__51236\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51234\ : std_logic;
signal \N__51233\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51230\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51223\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51215\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51209\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51202\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51199\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51196\ : std_logic;
signal \N__51195\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51192\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51189\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51182\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51173\ : std_logic;
signal \N__51172\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51170\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51167\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51165\ : std_logic;
signal \N__51164\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51162\ : std_logic;
signal \N__51161\ : std_logic;
signal \N__51160\ : std_logic;
signal \N__51159\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51157\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51147\ : std_logic;
signal \N__51146\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51144\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51141\ : std_logic;
signal \N__51140\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51138\ : std_logic;
signal \N__51137\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51135\ : std_logic;
signal \N__51134\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51132\ : std_logic;
signal \N__51131\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51128\ : std_logic;
signal \N__51127\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51124\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51117\ : std_logic;
signal \N__51116\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51114\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51109\ : std_logic;
signal \N__51108\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50672\ : std_logic;
signal \N__50669\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50656\ : std_logic;
signal \N__50653\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50644\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50633\ : std_logic;
signal \N__50630\ : std_logic;
signal \N__50627\ : std_logic;
signal \N__50624\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50609\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50604\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50601\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50599\ : std_logic;
signal \N__50598\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50596\ : std_logic;
signal \N__50595\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50593\ : std_logic;
signal \N__50590\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50570\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50560\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50554\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50550\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50511\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50508\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50504\ : std_logic;
signal \N__50503\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50477\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50468\ : std_logic;
signal \N__50465\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50413\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50384\ : std_logic;
signal \N__50377\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50340\ : std_logic;
signal \N__50339\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50337\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50331\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50328\ : std_logic;
signal \N__50327\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50317\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50314\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50311\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50303\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50300\ : std_logic;
signal \N__50297\ : std_logic;
signal \N__50294\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50287\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50284\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50281\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50275\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50272\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50270\ : std_logic;
signal \N__50269\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50267\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50264\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50259\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50253\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50212\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50203\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50200\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50152\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50144\ : std_logic;
signal \N__50143\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50135\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50127\ : std_logic;
signal \N__50124\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50115\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50111\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50093\ : std_logic;
signal \N__50092\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50090\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50057\ : std_logic;
signal \N__50054\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50048\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50018\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50005\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49996\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49966\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49763\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49753\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49734\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49716\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49695\ : std_logic;
signal \N__49688\ : std_logic;
signal \N__49685\ : std_logic;
signal \N__49682\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49631\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49550\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49547\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49544\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49528\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49508\ : std_logic;
signal \N__49507\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49504\ : std_logic;
signal \N__49499\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49485\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49472\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49469\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49266\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49263\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49257\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49228\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49222\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49201\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49199\ : std_logic;
signal \N__49198\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49196\ : std_logic;
signal \N__49195\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49178\ : std_logic;
signal \N__49175\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49158\ : std_logic;
signal \N__49155\ : std_logic;
signal \N__49150\ : std_logic;
signal \N__49145\ : std_logic;
signal \N__49142\ : std_logic;
signal \N__49139\ : std_logic;
signal \N__49136\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49130\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49118\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49079\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49049\ : std_logic;
signal \N__49046\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49040\ : std_logic;
signal \N__49037\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49024\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49012\ : std_logic;
signal \N__49011\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49007\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48978\ : std_logic;
signal \N__48977\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48947\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48930\ : std_logic;
signal \N__48927\ : std_logic;
signal \N__48924\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48900\ : std_logic;
signal \N__48889\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48679\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48658\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48544\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48539\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48497\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48387\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48382\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48380\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48364\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48246\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48070\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48067\ : std_logic;
signal \N__48064\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48046\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48023\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48007\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48005\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__48001\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47977\ : std_logic;
signal \N__47974\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47963\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47941\ : std_logic;
signal \N__47938\ : std_logic;
signal \N__47935\ : std_logic;
signal \N__47930\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47888\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47804\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47719\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47687\ : std_logic;
signal \N__47684\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47603\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47599\ : std_logic;
signal \N__47596\ : std_logic;
signal \N__47595\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47405\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47371\ : std_logic;
signal \N__47368\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47359\ : std_logic;
signal \N__47356\ : std_logic;
signal \N__47353\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47338\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47326\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47323\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47320\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47315\ : std_logic;
signal \N__47312\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47309\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47291\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47285\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47248\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47239\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47236\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47230\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47188\ : std_logic;
signal \N__47185\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47183\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47142\ : std_logic;
signal \N__47141\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46952\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46905\ : std_logic;
signal \N__46902\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46870\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46858\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46820\ : std_logic;
signal \N__46819\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46758\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46748\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46718\ : std_logic;
signal \N__46715\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46649\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46630\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46621\ : std_logic;
signal \N__46618\ : std_logic;
signal \N__46615\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46609\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46603\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46600\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46579\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46574\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46562\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46495\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46442\ : std_logic;
signal \N__46437\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46431\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46396\ : std_logic;
signal \N__46393\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46368\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46358\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46341\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46321\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46313\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46181\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46164\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46150\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46141\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46126\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46118\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46011\ : std_logic;
signal \N__46008\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__46003\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__46001\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45928\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45881\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45777\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45754\ : std_logic;
signal \N__45751\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45703\ : std_logic;
signal \N__45700\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45689\ : std_logic;
signal \N__45686\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45680\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45607\ : std_logic;
signal \N__45606\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45598\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45589\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45583\ : std_logic;
signal \N__45580\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45539\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45437\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45413\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45308\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45297\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45278\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45261\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45230\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45217\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45109\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44960\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44954\ : std_logic;
signal \N__44951\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44945\ : std_logic;
signal \N__44942\ : std_logic;
signal \N__44939\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44918\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44888\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44860\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44813\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44786\ : std_logic;
signal \N__44783\ : std_logic;
signal \N__44780\ : std_logic;
signal \N__44777\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44765\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44711\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44705\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44681\ : std_logic;
signal \N__44678\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44523\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44468\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44464\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44426\ : std_logic;
signal \N__44423\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44399\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44361\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44345\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44303\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44294\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44180\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44136\ : std_logic;
signal \N__44133\ : std_logic;
signal \N__44130\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44074\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44041\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44012\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43996\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43906\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43863\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43801\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43774\ : std_logic;
signal \N__43771\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43731\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43688\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43681\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43637\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43611\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43605\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43567\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43558\ : std_logic;
signal \N__43555\ : std_logic;
signal \N__43552\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43543\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43489\ : std_logic;
signal \N__43486\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43439\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43402\ : std_logic;
signal \N__43399\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43393\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43380\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43297\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43282\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43259\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43238\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43138\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43127\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43117\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43109\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43090\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43051\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43045\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43037\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42992\ : std_logic;
signal \N__42989\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42968\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42962\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42935\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42890\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42878\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42872\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42862\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42763\ : std_logic;
signal \N__42760\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42703\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42649\ : std_logic;
signal \N__42646\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42610\ : std_logic;
signal \N__42607\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42571\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42560\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42548\ : std_logic;
signal \N__42545\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42533\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42523\ : std_logic;
signal \N__42520\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42496\ : std_logic;
signal \N__42493\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42441\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42299\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42280\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42228\ : std_logic;
signal \N__42225\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42197\ : std_logic;
signal \N__42194\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42161\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42088\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42059\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42028\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42022\ : std_logic;
signal \N__42017\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41860\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41849\ : std_logic;
signal \N__41846\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41801\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41789\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41674\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41618\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41612\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41600\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41578\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41524\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41479\ : std_logic;
signal \N__41476\ : std_logic;
signal \N__41473\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41467\ : std_logic;
signal \N__41464\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41429\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41404\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41380\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41362\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41340\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41323\ : std_logic;
signal \N__41320\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41314\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41288\ : std_logic;
signal \N__41285\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41257\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41210\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41204\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41155\ : std_logic;
signal \N__41152\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41114\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41089\ : std_logic;
signal \N__41086\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41068\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41039\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40969\ : std_logic;
signal \N__40966\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40944\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40903\ : std_logic;
signal \N__40900\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40880\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40834\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40783\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40753\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40730\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40706\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40546\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40534\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40460\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40457\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40346\ : std_logic;
signal \N__40345\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40304\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40294\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40258\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40252\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40241\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40123\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40117\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39766\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39746\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39728\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39700\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39629\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39556\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39440\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39275\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39256\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39167\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39149\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39068\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38971\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38965\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38908\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38875\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38837\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38834\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38735\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38704\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38683\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38669\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38642\ : std_logic;
signal \N__38639\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38444\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38381\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38306\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38108\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38090\ : std_logic;
signal \N__38087\ : std_logic;
signal \N__38084\ : std_logic;
signal \N__38081\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38048\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37976\ : std_logic;
signal \N__37967\ : std_logic;
signal \N__37964\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37949\ : std_logic;
signal \N__37946\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37889\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37778\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37755\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37670\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37553\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37481\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37441\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37387\ : std_logic;
signal \N__37384\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37370\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37349\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37345\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37315\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37136\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37070\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36725\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36577\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36323\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36310\ : std_logic;
signal \N__36307\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36229\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35908\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35825\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35765\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35753\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35650\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35554\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35339\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35190\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34538\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34520\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34493\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34118\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34010\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33638\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33328\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33157\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32624\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32444\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31394\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31379\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31292\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31174\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30839\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30518\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30497\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29078\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28493\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27674\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26657\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24299\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \ICE_GPMO_2\ : std_logic;
signal \M_CLK4\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN_net\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN_net\ : std_logic;
signal \ICE_SYSCLK\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN_net\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN_net\ : std_logic;
signal \n25_cascade_\ : std_logic;
signal n27_adj_1173 : std_logic;
signal \n14114_cascade_\ : std_logic;
signal \n10522_cascade_\ : std_logic;
signal \TEST_LED\ : std_logic;
signal n28 : std_logic;
signal n26_adj_1180 : std_logic;
signal n10 : std_logic;
signal \DDS_MCLK1\ : std_logic;
signal secclk_cnt_0 : std_logic;
signal \bfn_3_7_0_\ : std_logic;
signal secclk_cnt_1 : std_logic;
signal n14009 : std_logic;
signal secclk_cnt_2 : std_logic;
signal n14010 : std_logic;
signal secclk_cnt_3 : std_logic;
signal n14011 : std_logic;
signal secclk_cnt_4 : std_logic;
signal n14012 : std_logic;
signal secclk_cnt_5 : std_logic;
signal n14013 : std_logic;
signal secclk_cnt_6 : std_logic;
signal n14014 : std_logic;
signal secclk_cnt_7 : std_logic;
signal n14015 : std_logic;
signal n14016 : std_logic;
signal secclk_cnt_8 : std_logic;
signal \bfn_3_8_0_\ : std_logic;
signal secclk_cnt_9 : std_logic;
signal n14017 : std_logic;
signal secclk_cnt_10 : std_logic;
signal n14018 : std_logic;
signal secclk_cnt_11 : std_logic;
signal n14019 : std_logic;
signal n14020 : std_logic;
signal secclk_cnt_13 : std_logic;
signal n14021 : std_logic;
signal secclk_cnt_14 : std_logic;
signal n14022 : std_logic;
signal secclk_cnt_15 : std_logic;
signal n14023 : std_logic;
signal n14024 : std_logic;
signal secclk_cnt_16 : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal secclk_cnt_17 : std_logic;
signal n14025 : std_logic;
signal secclk_cnt_18 : std_logic;
signal n14026 : std_logic;
signal n14027 : std_logic;
signal secclk_cnt_20 : std_logic;
signal n14028 : std_logic;
signal n14029 : std_logic;
signal n14030 : std_logic;
signal \clk_16MHz\ : std_logic;
signal n10522 : std_logic;
signal buf_adcdata2_0 : std_logic;
signal cmd_rdadctmp_8_adj_1068 : std_logic;
signal cmd_rdadctmp_7_adj_1069 : std_logic;
signal cmd_rdadctmp_6_adj_1070 : std_logic;
signal cmd_rdadctmp_5_adj_1071 : std_logic;
signal cmd_rdadctmp_3_adj_1073 : std_logic;
signal cmd_rdadctmp_4_adj_1072 : std_logic;
signal \n14_adj_1035_cascade_\ : std_logic;
signal \M_CS2\ : std_logic;
signal n15165 : std_logic;
signal \M_MISO2\ : std_logic;
signal \n8302_cascade_\ : std_logic;
signal cmd_rdadctmp_2_adj_1074 : std_logic;
signal cmd_rdadctmp_0_adj_1076 : std_logic;
signal cmd_rdadctmp_1_adj_1075 : std_logic;
signal buf_data2_6 : std_logic;
signal buf_adcdata4_7 : std_logic;
signal buf_data2_7 : std_logic;
signal buf_data2_4 : std_logic;
signal \n4304_cascade_\ : std_logic;
signal buf_data2_5 : std_logic;
signal \n4303_cascade_\ : std_logic;
signal n4302 : std_logic;
signal n4301 : std_logic;
signal buf_data2_0 : std_logic;
signal buf_data2_1 : std_logic;
signal buf_data2_2 : std_logic;
signal n4307 : std_logic;
signal n4306 : std_logic;
signal n4308 : std_logic;
signal buf_adcdata2_5 : std_logic;
signal buf_adcdata2_6 : std_logic;
signal buf_adcdata2_7 : std_logic;
signal cmd_rdadctmp_15_adj_1061 : std_logic;
signal buf_adcdata2_3 : std_logic;
signal buf_adcdata2_4 : std_logic;
signal cmd_rdadctmp_13_adj_1063 : std_logic;
signal cmd_rdadctmp_14_adj_1062 : std_logic;
signal cmd_rdadctmp_11_adj_1065 : std_logic;
signal cmd_rdadctmp_12_adj_1064 : std_logic;
signal buf_adcdata1_5 : std_logic;
signal buf_adcdata1_7 : std_logic;
signal buf_adcdata4_5 : std_logic;
signal cmd_rdadctmp_13_adj_1136 : std_logic;
signal cmd_rdadctmp_14_adj_1135 : std_logic;
signal buf_adcdata4_6 : std_logic;
signal cmd_rdadctmp_15_adj_1134 : std_logic;
signal buf_adcdata4_0 : std_logic;
signal buf_adcdata4_1 : std_logic;
signal cmd_rdadctmp_9_adj_1140 : std_logic;
signal cmd_rdadctmp_10_adj_1139 : std_logic;
signal buf_adcdata4_2 : std_logic;
signal cmd_rdadctmp_7_adj_1142 : std_logic;
signal cmd_rdadctmp_8_adj_1141 : std_logic;
signal cmd_rdadctmp_5_adj_1144 : std_logic;
signal cmd_rdadctmp_6_adj_1143 : std_logic;
signal cmd_rdadctmp_11_adj_1138 : std_logic;
signal cmd_rdadctmp_4_adj_1145 : std_logic;
signal cmd_rdadctmp_3_adj_1146 : std_logic;
signal cmd_rdadctmp_2_adj_1147 : std_logic;
signal cmd_rdadctmp_12_adj_1137 : std_logic;
signal buf_adcdata4_4 : std_logic;
signal buf_data1_6 : std_logic;
signal n4146 : std_logic;
signal buf_data1_0 : std_logic;
signal buf_data1_7 : std_logic;
signal n4145 : std_logic;
signal n4152 : std_logic;
signal \n15131_cascade_\ : std_logic;
signal \n8738_cascade_\ : std_logic;
signal n8847 : std_logic;
signal \n8847_cascade_\ : std_logic;
signal n10611 : std_logic;
signal \n8787_cascade_\ : std_logic;
signal buf_data1_2 : std_logic;
signal \n4150_cascade_\ : std_logic;
signal buf_data1_4 : std_logic;
signal \n4148_cascade_\ : std_logic;
signal buf_data1_5 : std_logic;
signal \n4147_cascade_\ : std_logic;
signal n8738 : std_logic;
signal n10590 : std_logic;
signal secclk_cnt_21 : std_logic;
signal secclk_cnt_19 : std_logic;
signal secclk_cnt_12 : std_logic;
signal secclk_cnt_22 : std_logic;
signal n14_adj_1163 : std_logic;
signal buf_data2_10 : std_logic;
signal \n4062_cascade_\ : std_logic;
signal buf_adcdata3_2 : std_logic;
signal cmd_rdadctmp_11_adj_1101 : std_logic;
signal buf_adcdata1_3 : std_logic;
signal buf_adcdata3_4 : std_logic;
signal cmd_rdadctmp_1 : std_logic;
signal buf_adcdata3_7 : std_logic;
signal \M_MISO1\ : std_logic;
signal cmd_rdadctmp_0 : std_logic;
signal cmd_rdadctmp_12_adj_1100 : std_logic;
signal buf_adcdata1_4 : std_logic;
signal cmd_rdadctmp_2 : std_logic;
signal cmd_rdadctmp_7 : std_logic;
signal cmd_rdadctmp_6 : std_logic;
signal cmd_rdadctmp_5 : std_logic;
signal cmd_rdadctmp_3 : std_logic;
signal cmd_rdadctmp_4 : std_logic;
signal n15168 : std_logic;
signal \n15168_cascade_\ : std_logic;
signal \M_CS1\ : std_logic;
signal n14_adj_1039 : std_logic;
signal \M_SCLK1\ : std_logic;
signal \ADC_VAC1.n9312_cascade_\ : std_logic;
signal \ADC_VAC1.n15338_cascade_\ : std_logic;
signal \ADC_VAC1.n15360_cascade_\ : std_logic;
signal \ADC_VAC1.bit_cnt_0\ : std_logic;
signal \bfn_6_16_0_\ : std_logic;
signal \ADC_VAC1.bit_cnt_1\ : std_logic;
signal \ADC_VAC1.n13981\ : std_logic;
signal \ADC_VAC1.bit_cnt_2\ : std_logic;
signal \ADC_VAC1.n13982\ : std_logic;
signal \ADC_VAC1.bit_cnt_3\ : std_logic;
signal \ADC_VAC1.n13983\ : std_logic;
signal \ADC_VAC1.bit_cnt_4\ : std_logic;
signal \ADC_VAC1.n13984\ : std_logic;
signal \ADC_VAC1.bit_cnt_5\ : std_logic;
signal \ADC_VAC1.n13985\ : std_logic;
signal \ADC_VAC1.bit_cnt_6\ : std_logic;
signal \ADC_VAC1.n13986\ : std_logic;
signal \ADC_VAC1.n13987\ : std_logic;
signal \ADC_VAC1.bit_cnt_7\ : std_logic;
signal \ADC_VAC1.n9312\ : std_logic;
signal \ADC_VAC1.n10667\ : std_logic;
signal \n16470_cascade_\ : std_logic;
signal comm_buf_5_5 : std_logic;
signal comm_buf_2_5 : std_logic;
signal \n16416_cascade_\ : std_logic;
signal n16473 : std_logic;
signal \n16419_cascade_\ : std_logic;
signal \n7_adj_1238_cascade_\ : std_logic;
signal buf_data2_21 : std_logic;
signal \n4103_cascade_\ : std_logic;
signal comm_buf_3_5 : std_logic;
signal buf_data2_17 : std_logic;
signal \n4107_cascade_\ : std_logic;
signal buf_data2_18 : std_logic;
signal n8787 : std_logic;
signal n10599 : std_logic;
signal comm_buf_2_2 : std_logic;
signal \n15388_cascade_\ : std_logic;
signal \n16389_cascade_\ : std_logic;
signal comm_buf_4_2 : std_logic;
signal comm_buf_5_2 : std_logic;
signal n15448 : std_logic;
signal \n15447_cascade_\ : std_logic;
signal n16386 : std_logic;
signal buf_adcdata4_18 : std_logic;
signal comm_buf_2_3 : std_logic;
signal comm_buf_4_3 : std_logic;
signal comm_buf_5_3 : std_logic;
signal \n16440_cascade_\ : std_logic;
signal n15423 : std_logic;
signal n15397 : std_logic;
signal \n16392_cascade_\ : std_logic;
signal n16443 : std_logic;
signal \n16395_cascade_\ : std_logic;
signal \M_SCLK2\ : std_logic;
signal buf_adcdata3_5 : std_logic;
signal buf_adcdata3_6 : std_logic;
signal cmd_rdadctmp_12 : std_logic;
signal cmd_rdadctmp_10_adj_1102 : std_logic;
signal cmd_rdadctmp_16_adj_1133 : std_logic;
signal cmd_rdadctmp_17_adj_1132 : std_logic;
signal cmd_rdadctmp_18_adj_1131 : std_logic;
signal buf_adcdata4_10 : std_logic;
signal \ADC_VAC1.n15263_cascade_\ : std_logic;
signal \ADC_VAC1.n15553\ : std_logic;
signal \ADC_VAC1.n15264\ : std_logic;
signal \M_DRDY1\ : std_logic;
signal \ADC_VAC1.n17_cascade_\ : std_logic;
signal \ADC_VAC1.n12\ : std_logic;
signal cmd_rdadctmp_13 : std_logic;
signal cmd_rdadctmp_1_adj_1148 : std_logic;
signal \M_MISO4\ : std_logic;
signal cmd_rdadctmp_0_adj_1149 : std_logic;
signal cmd_rdadctmp_15 : std_logic;
signal \M_START\ : std_logic;
signal comm_buf_3_0 : std_logic;
signal comm_buf_2_0 : std_logic;
signal \n16413_cascade_\ : std_logic;
signal comm_buf_5_6 : std_logic;
signal \n16518_cascade_\ : std_logic;
signal n13493 : std_logic;
signal \n16521_cascade_\ : std_logic;
signal comm_buf_2_6 : std_logic;
signal comm_buf_3_6 : std_logic;
signal n16410 : std_logic;
signal n16491 : std_logic;
signal comm_buf_2_1 : std_logic;
signal comm_buf_3_1 : std_logic;
signal \n16404_cascade_\ : std_logic;
signal \n16407_cascade_\ : std_logic;
signal comm_buf_5_1 : std_logic;
signal comm_buf_4_1 : std_logic;
signal n16515 : std_logic;
signal n16512 : std_logic;
signal n7_adj_1240 : std_logic;
signal \n16425_cascade_\ : std_logic;
signal buf_data2_12 : std_logic;
signal \n4060_cascade_\ : std_logic;
signal comm_buf_4_5 : std_logic;
signal comm_buf_4_6 : std_logic;
signal buf_data2_15 : std_logic;
signal \n4057_cascade_\ : std_logic;
signal n10604 : std_logic;
signal buf_adcdata1_17 : std_logic;
signal buf_adcdata1_18 : std_logic;
signal cmd_rdadctmp_26 : std_logic;
signal cmd_rdadctmp_27 : std_logic;
signal buf_adcdata1_19 : std_logic;
signal cmd_rdadctmp_25 : std_logic;
signal buf_adcdata1_20 : std_logic;
signal \n84_cascade_\ : std_logic;
signal \n15593_cascade_\ : std_logic;
signal \n8045_cascade_\ : std_logic;
signal n15573 : std_logic;
signal cmd_rdadctmp_11 : std_logic;
signal buf_adcdata4_12 : std_logic;
signal cmd_rdadctmp_16_adj_1060 : std_logic;
signal buf_adcdata2_8 : std_logic;
signal cmd_rdadctmp_9_adj_1103 : std_logic;
signal cmd_rdadctmp_28 : std_logic;
signal buf_adcdata2_17 : std_logic;
signal cmd_rdadctmp_13_adj_1099 : std_logic;
signal cmd_rdadctmp_14_adj_1098 : std_logic;
signal buf_data2_14 : std_logic;
signal n4058 : std_logic;
signal \n14_adj_1031_cascade_\ : std_logic;
signal \M_CS3\ : std_logic;
signal \M_SCLK3\ : std_logic;
signal cmd_rdadctmp_4_adj_1108 : std_logic;
signal \DTRIG_N_957\ : std_logic;
signal adc_state_1 : std_logic;
signal \M_MISO3\ : std_logic;
signal cmd_rdadctmp_0_adj_1112 : std_logic;
signal cmd_rdadctmp_1_adj_1111 : std_logic;
signal \ADC_VAC3.n12\ : std_logic;
signal n15162 : std_logic;
signal \n15162_cascade_\ : std_logic;
signal \comm_spi.n16911\ : std_logic;
signal \comm_spi.n10433\ : std_logic;
signal \comm_spi.n16911_cascade_\ : std_logic;
signal \comm_spi.data_tx_7__N_811\ : std_logic;
signal \comm_spi.data_tx_7__N_831\ : std_logic;
signal \comm_spi.data_tx_7__N_812\ : std_logic;
signal comm_tx_buf_1 : std_logic;
signal n15411 : std_logic;
signal \n16446_cascade_\ : std_logic;
signal n15391 : std_logic;
signal n16449 : std_logic;
signal buf_data2_3 : std_logic;
signal buf_adcdata4_3 : std_logic;
signal n4305 : std_logic;
signal n16431 : std_logic;
signal comm_buf_4_0 : std_logic;
signal \n16506_cascade_\ : std_logic;
signal comm_buf_5_0 : std_logic;
signal n16509 : std_logic;
signal n15424 : std_logic;
signal n15412 : std_logic;
signal comm_buf_5_7 : std_logic;
signal comm_buf_4_7 : std_logic;
signal \n16482_cascade_\ : std_logic;
signal n16485 : std_logic;
signal \INVcomm_spi.imiso_83_7340_7341_resetC_net\ : std_logic;
signal \comm_buf_3_7_N_501_2\ : std_logic;
signal comm_buf_3_2 : std_logic;
signal comm_buf_3_3 : std_logic;
signal buf_data4_19 : std_logic;
signal comm_buf_9_3 : std_logic;
signal buf_data4_20 : std_logic;
signal \n66_adj_1153_cascade_\ : std_logic;
signal \DDS_SCK1\ : std_logic;
signal \DDS_MOSI1\ : std_logic;
signal n15522 : std_logic;
signal n15523 : std_logic;
signal \n16398_cascade_\ : std_logic;
signal \n16401_cascade_\ : std_logic;
signal \n109_adj_1155_cascade_\ : std_logic;
signal \n8048_cascade_\ : std_logic;
signal n15578 : std_logic;
signal buf_adcdata1_21 : std_logic;
signal buf_adcdata1_22 : std_logic;
signal cmd_rdadctmp_24_adj_1052 : std_logic;
signal buf_adcdata2_16 : std_logic;
signal cmd_rdadctmp_29 : std_logic;
signal cmd_rdadctmp_30 : std_logic;
signal buf_adcdata1_1 : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \ADC_VAC2.n13988\ : std_logic;
signal \ADC_VAC2.n13989\ : std_logic;
signal \ADC_VAC2.n13990\ : std_logic;
signal \ADC_VAC2.n13991\ : std_logic;
signal \ADC_VAC2.n13992\ : std_logic;
signal \ADC_VAC2.n13993\ : std_logic;
signal \ADC_VAC2.n13994\ : std_logic;
signal \ADC_VAC2.bit_cnt_1\ : std_logic;
signal \ADC_VAC2.bit_cnt_7\ : std_logic;
signal \ADC_VAC2.n15261_cascade_\ : std_logic;
signal \ADC_VAC2.n15595\ : std_logic;
signal \ADC_VAC2.n15262\ : std_logic;
signal \ADC_VAC2.bit_cnt_6\ : std_logic;
signal \ADC_VAC2.bit_cnt_0\ : std_logic;
signal \ADC_VAC2.n16\ : std_logic;
signal \ADC_VAC2.n17_cascade_\ : std_logic;
signal cmd_rdadctmp_2_adj_1110 : std_logic;
signal cmd_rdadctmp_3_adj_1109 : std_logic;
signal acadc_dtrig2 : std_logic;
signal acadc_dtrig1 : std_logic;
signal acadc_dtrig4 : std_logic;
signal acadc_dtrig3 : std_logic;
signal cmd_rdadctmp_14 : std_logic;
signal buf_adcdata1_6 : std_logic;
signal cmd_rdadctmp_15_adj_1097 : std_logic;
signal \M_SCLK4\ : std_logic;
signal \comm_spi.n10434\ : std_logic;
signal comm_tx_buf_0 : std_logic;
signal \comm_spi.data_tx_7__N_834\ : std_logic;
signal n16428 : std_logic;
signal buf_data2_20 : std_logic;
signal n4104 : std_logic;
signal comm_buf_3_7 : std_logic;
signal comm_buf_2_7 : std_logic;
signal \n15382_cascade_\ : std_logic;
signal \n16383_cascade_\ : std_logic;
signal \n16494_cascade_\ : std_logic;
signal n16497 : std_logic;
signal n15450 : std_logic;
signal \n15451_cascade_\ : std_logic;
signal n16380 : std_logic;
signal buf_data4_1 : std_logic;
signal buf_data4_2 : std_logic;
signal comm_buf_11_2 : std_logic;
signal buf_data4_3 : std_logic;
signal comm_buf_11_3 : std_logic;
signal buf_data4_4 : std_logic;
signal buf_data4_5 : std_logic;
signal comm_buf_11_5 : std_logic;
signal buf_data4_6 : std_logic;
signal buf_data4_7 : std_logic;
signal comm_buf_11_7 : std_logic;
signal buf_data4_0 : std_logic;
signal comm_buf_11_0 : std_logic;
signal buf_data3_15 : std_logic;
signal comm_buf_7_7 : std_logic;
signal buf_data3_8 : std_logic;
signal comm_buf_7_0 : std_logic;
signal buf_data3_14 : std_logic;
signal comm_buf_7_6 : std_logic;
signal buf_data3_13 : std_logic;
signal comm_buf_7_5 : std_logic;
signal buf_data3_12 : std_logic;
signal buf_data3_11 : std_logic;
signal comm_buf_7_3 : std_logic;
signal buf_data3_10 : std_logic;
signal comm_buf_7_2 : std_logic;
signal buf_data3_9 : std_logic;
signal comm_buf_7_1 : std_logic;
signal comm_buf_3_4 : std_logic;
signal comm_buf_2_4 : std_logic;
signal \n15403_cascade_\ : std_logic;
signal \n16479_cascade_\ : std_logic;
signal n10660 : std_logic;
signal comm_buf_7_4 : std_logic;
signal comm_buf_11_4 : std_logic;
signal comm_buf_9_4 : std_logic;
signal \n16452_cascade_\ : std_logic;
signal n16455 : std_logic;
signal comm_buf_5_4 : std_logic;
signal comm_buf_4_4 : std_logic;
signal n15400 : std_logic;
signal \n15399_cascade_\ : std_logic;
signal n16476 : std_logic;
signal \n15633_cascade_\ : std_logic;
signal \n16458_cascade_\ : std_logic;
signal \n16461_cascade_\ : std_logic;
signal \n76_cascade_\ : std_logic;
signal \n4_adj_1195_cascade_\ : std_logic;
signal n15632 : std_logic;
signal n15589 : std_logic;
signal \n87_adj_1165_cascade_\ : std_logic;
signal \n69_adj_1161_cascade_\ : std_logic;
signal n130 : std_logic;
signal n8050 : std_logic;
signal n8089 : std_logic;
signal n96_adj_1159 : std_logic;
signal \n130_adj_1156_cascade_\ : std_logic;
signal n15587 : std_logic;
signal \n8051_cascade_\ : std_logic;
signal cmd_rdadctmp_19_adj_1130 : std_logic;
signal cmd_rdadctmp_8 : std_logic;
signal buf_adcdata1_0 : std_logic;
signal cmd_rdadctmp_23 : std_logic;
signal buf_adcdata1_15 : std_logic;
signal cmd_rdadctmp_20_adj_1129 : std_logic;
signal \ADC_VAC2.bit_cnt_4\ : std_logic;
signal \ADC_VAC2.bit_cnt_3\ : std_logic;
signal \ADC_VAC2.bit_cnt_5\ : std_logic;
signal \ADC_VAC2.bit_cnt_2\ : std_logic;
signal \ADC_VAC2.n15596\ : std_logic;
signal \ADC_VAC3.n15334_cascade_\ : std_logic;
signal \ADC_VAC3.n15358_cascade_\ : std_logic;
signal \ADC_VAC3.n15602_cascade_\ : std_logic;
signal \ADC_VAC3.n15260\ : std_logic;
signal \ADC_VAC3.n15259\ : std_logic;
signal \ADC_VAC3.n17\ : std_logic;
signal \ADC_VAC3.bit_cnt_0\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \ADC_VAC3.bit_cnt_1\ : std_logic;
signal \ADC_VAC3.n13995\ : std_logic;
signal \ADC_VAC3.bit_cnt_2\ : std_logic;
signal \ADC_VAC3.n13996\ : std_logic;
signal \ADC_VAC3.bit_cnt_3\ : std_logic;
signal \ADC_VAC3.n13997\ : std_logic;
signal \ADC_VAC3.bit_cnt_4\ : std_logic;
signal \ADC_VAC3.n13998\ : std_logic;
signal \ADC_VAC3.bit_cnt_5\ : std_logic;
signal \ADC_VAC3.n13999\ : std_logic;
signal \ADC_VAC3.bit_cnt_6\ : std_logic;
signal \ADC_VAC3.n14000\ : std_logic;
signal \ADC_VAC3.n14001\ : std_logic;
signal \ADC_VAC3.bit_cnt_7\ : std_logic;
signal cmd_rdadctmp_31 : std_logic;
signal buf_adcdata1_23 : std_logic;
signal \M_DRDY3\ : std_logic;
signal adc_state_1_adj_1079 : std_logic;
signal \ADC_VAC3.n9514\ : std_logic;
signal \DTRIG_N_957_adj_1114\ : std_logic;
signal \ADC_VAC3.n9514_cascade_\ : std_logic;
signal \ADC_VAC3.n10744\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \ADC_VAC4.n14002\ : std_logic;
signal \ADC_VAC4.n14003\ : std_logic;
signal \ADC_VAC4.n14004\ : std_logic;
signal \ADC_VAC4.n14005\ : std_logic;
signal \ADC_VAC4.n14006\ : std_logic;
signal \ADC_VAC4.n14007\ : std_logic;
signal \ADC_VAC4.n14008\ : std_logic;
signal \comm_spi.n16908\ : std_logic;
signal \comm_spi.n10459\ : std_logic;
signal \comm_spi.n10460\ : std_logic;
signal \comm_spi.data_tx_7__N_828\ : std_logic;
signal buf_adcdata4_21 : std_logic;
signal cmd_rdadctmp_29_adj_1120 : std_logic;
signal cmd_rdadctmp_30_adj_1119 : std_logic;
signal cmd_rdadctmp_31_adj_1118 : std_logic;
signal buf_data3_7 : std_logic;
signal comm_buf_8_7 : std_logic;
signal buf_data3_6 : std_logic;
signal comm_buf_8_6 : std_logic;
signal buf_data3_5 : std_logic;
signal comm_buf_8_5 : std_logic;
signal buf_data3_4 : std_logic;
signal comm_buf_8_4 : std_logic;
signal buf_data3_3 : std_logic;
signal comm_buf_8_3 : std_logic;
signal buf_data3_2 : std_logic;
signal comm_buf_8_2 : std_logic;
signal buf_data3_1 : std_logic;
signal comm_buf_8_1 : std_logic;
signal buf_data3_0 : std_logic;
signal comm_buf_8_0 : std_logic;
signal buf_data3_23 : std_logic;
signal comm_buf_6_7 : std_logic;
signal buf_data3_22 : std_logic;
signal comm_buf_6_6 : std_logic;
signal buf_data3_21 : std_logic;
signal comm_buf_6_5 : std_logic;
signal buf_data3_20 : std_logic;
signal comm_buf_6_4 : std_logic;
signal buf_data3_19 : std_logic;
signal comm_buf_6_3 : std_logic;
signal buf_data3_18 : std_logic;
signal comm_buf_6_2 : std_logic;
signal \n8907_cascade_\ : std_logic;
signal n8943 : std_logic;
signal \n8943_cascade_\ : std_logic;
signal n10625 : std_logic;
signal n9123 : std_logic;
signal \n9123_cascade_\ : std_logic;
signal n10653 : std_logic;
signal buf_data3_16 : std_logic;
signal comm_buf_6_0 : std_logic;
signal buf_data3_17 : std_logic;
signal comm_buf_6_1 : std_logic;
signal n8907 : std_logic;
signal n10618 : std_logic;
signal buf_data4_10 : std_logic;
signal comm_buf_10_2 : std_logic;
signal buf_data4_11 : std_logic;
signal comm_buf_10_3 : std_logic;
signal buf_data4_12 : std_logic;
signal comm_buf_10_4 : std_logic;
signal buf_data4_15 : std_logic;
signal comm_buf_10_7 : std_logic;
signal buf_data4_8 : std_logic;
signal comm_buf_10_0 : std_logic;
signal \n16434_cascade_\ : std_logic;
signal \n16437_cascade_\ : std_logic;
signal n109 : std_logic;
signal \n8054_cascade_\ : std_logic;
signal n59 : std_logic;
signal cmd_rdadctmp_25_adj_1087 : std_logic;
signal cmd_rdadctmp_7_adj_1105 : std_logic;
signal \n16500_cascade_\ : std_logic;
signal \n16503_cascade_\ : std_logic;
signal n4_adj_1280 : std_logic;
signal \n8047_cascade_\ : std_logic;
signal n10576 : std_logic;
signal cmd_rdadctmp_9 : std_logic;
signal buf_control_3 : std_logic;
signal n69_adj_1029 : std_logic;
signal buf_adcdata4_14 : std_logic;
signal buf_adcdata3_20 : std_logic;
signal n61 : std_logic;
signal buf_control_4 : std_logic;
signal n69 : std_logic;
signal buf_control_0 : std_logic;
signal buf_data2_8 : std_logic;
signal buf_adcdata4_8 : std_logic;
signal n4064 : std_logic;
signal cmd_rdadctmp_5_adj_1107 : std_logic;
signal cmd_rdadctmp_6_adj_1106 : std_logic;
signal cmd_rdadctmp_28_adj_1084 : std_logic;
signal buf_adcdata1_9 : std_logic;
signal cmd_rdadctmp_17 : std_logic;
signal cmd_rdadctmp_19 : std_logic;
signal buf_adcdata1_11 : std_logic;
signal buf_adcdata3_8 : std_logic;
signal \ADC_VAC4.bit_cnt_4\ : std_logic;
signal \ADC_VAC4.bit_cnt_3\ : std_logic;
signal \ADC_VAC4.bit_cnt_1\ : std_logic;
signal \ADC_VAC4.bit_cnt_2\ : std_logic;
signal \ADC_VAC4.bit_cnt_6\ : std_logic;
signal \ADC_VAC4.bit_cnt_0\ : std_logic;
signal \ADC_VAC4.n15330_cascade_\ : std_logic;
signal \ADC_VAC4.bit_cnt_7\ : std_logic;
signal \ADC_VAC4.bit_cnt_5\ : std_logic;
signal \ADC_VAC4.n15354\ : std_logic;
signal \ADC_VAC4.n15619_cascade_\ : std_logic;
signal \ADC_VAC4.n9631\ : std_logic;
signal \ADC_VAC4.n9631_cascade_\ : std_logic;
signal \ADC_VAC4.n10783\ : std_logic;
signal buf_adcdata4_20 : std_logic;
signal \comm_spi.n16905_cascade_\ : std_logic;
signal \comm_spi.data_tx_7__N_809\ : std_logic;
signal comm_tx_buf_2 : std_logic;
signal \comm_spi.data_tx_7__N_810\ : std_logic;
signal \comm_spi.n16905\ : std_logic;
signal \comm_spi.n10463\ : std_logic;
signal \comm_spi.n10464\ : std_logic;
signal buf_data4_21 : std_logic;
signal comm_buf_9_5 : std_logic;
signal buf_data4_22 : std_logic;
signal comm_buf_9_6 : std_logic;
signal buf_data4_23 : std_logic;
signal comm_buf_9_7 : std_logic;
signal buf_data4_18 : std_logic;
signal comm_buf_9_2 : std_logic;
signal buf_data4_17 : std_logic;
signal comm_buf_9_1 : std_logic;
signal \n15161_cascade_\ : std_logic;
signal n8997 : std_logic;
signal \n8997_cascade_\ : std_logic;
signal n10632 : std_logic;
signal buf_data4_16 : std_logic;
signal comm_buf_9_0 : std_logic;
signal n9027 : std_logic;
signal n10639 : std_logic;
signal comm_buf_11_1 : std_logic;
signal n16422 : std_logic;
signal buf_data4_9 : std_logic;
signal comm_buf_10_1 : std_logic;
signal n8763 : std_logic;
signal n13470 : std_logic;
signal n13497 : std_logic;
signal \n13497_cascade_\ : std_logic;
signal \n9045_cascade_\ : std_logic;
signal comm_buf_11_6 : std_logic;
signal n16488 : std_logic;
signal buf_data4_14 : std_logic;
signal comm_buf_10_6 : std_logic;
signal \n13457_cascade_\ : std_logic;
signal \n15565_cascade_\ : std_logic;
signal \n13_adj_1257_cascade_\ : std_logic;
signal n8823 : std_logic;
signal n41 : std_logic;
signal n13457 : std_logic;
signal n13458 : std_logic;
signal buf_data4_13 : std_logic;
signal comm_buf_10_5 : std_logic;
signal n9045 : std_logic;
signal n10646 : std_logic;
signal \n11_adj_1279_cascade_\ : std_logic;
signal n8654 : std_logic;
signal n5 : std_logic;
signal n15221 : std_logic;
signal \n17_cascade_\ : std_logic;
signal \n8702_cascade_\ : std_logic;
signal bit_cnt_3 : std_logic;
signal bit_cnt_2 : std_logic;
signal bit_cnt_0 : std_logic;
signal \n16524_cascade_\ : std_logic;
signal \n16527_cascade_\ : std_logic;
signal \n4_adj_1264_cascade_\ : std_logic;
signal n8055 : std_logic;
signal buf_adcdata4_15 : std_logic;
signal n15144 : std_logic;
signal buf_adcdata4_17 : std_logic;
signal n71 : std_logic;
signal cmd_rdadctmp_26_adj_1123 : std_logic;
signal cmd_rdadctmp_27_adj_1085 : std_logic;
signal buf_adcdata3_23 : std_logic;
signal cmd_rdadctmp_27_adj_1122 : std_logic;
signal cmd_rdadctmp_28_adj_1121 : std_logic;
signal cmd_rdadctmp_23_adj_1126 : std_logic;
signal cmd_rdadctmp_24_adj_1125 : std_logic;
signal cmd_rdadctmp_25_adj_1124 : std_logic;
signal \M_POW\ : std_logic;
signal buf_adcdata3_19 : std_logic;
signal n87 : std_logic;
signal n8272 : std_logic;
signal cmd_rdadctmp_26_adj_1086 : std_logic;
signal buf_adcdata3_18 : std_logic;
signal n15811 : std_logic;
signal cmd_rdadctmp_21_adj_1128 : std_logic;
signal cmd_rdadctmp_22_adj_1127 : std_logic;
signal buf_adcdata3_16 : std_logic;
signal n90 : std_logic;
signal \n15156_cascade_\ : std_logic;
signal n9694 : std_logic;
signal \ADC_VAC4.n15257_cascade_\ : std_logic;
signal \ADC_VAC4.n15258\ : std_logic;
signal \ADC_VAC4.n15278\ : std_logic;
signal \M_DRDY4\ : std_logic;
signal \n14_cascade_\ : std_logic;
signal n15156 : std_logic;
signal \M_CS4\ : std_logic;
signal buf_data2_11 : std_logic;
signal buf_adcdata4_11 : std_logic;
signal n4061 : std_logic;
signal \ADC_VAC4.n17\ : std_logic;
signal adc_state_0_adj_1117 : std_logic;
signal \DTRIG_N_957_adj_1150\ : std_logic;
signal adc_state_1_adj_1116 : std_logic;
signal \ADC_VAC4.n12\ : std_logic;
signal \ADC_VAC4.n14930\ : std_logic;
signal \comm_spi.n10467\ : std_logic;
signal \comm_spi.n10468\ : std_logic;
signal \comm_spi.data_tx_7__N_822\ : std_logic;
signal \DDS_CS1\ : std_logic;
signal comm_tx_buf_7 : std_logic;
signal comm_tx_buf_6 : std_logic;
signal \comm_spi.n16884\ : std_logic;
signal buf_data1_23 : std_logic;
signal \n18_cascade_\ : std_logic;
signal \n15466_cascade_\ : std_logic;
signal n104 : std_logic;
signal n56 : std_logic;
signal buf_adcdata3_1 : std_logic;
signal buf_data1_1 : std_logic;
signal n4151 : std_logic;
signal \n15567_cascade_\ : std_logic;
signal n7_adj_1255 : std_logic;
signal n6 : std_logic;
signal \n5_adj_1235_cascade_\ : std_logic;
signal \n15535_cascade_\ : std_logic;
signal \n15_cascade_\ : std_logic;
signal n9021 : std_logic;
signal n4814 : std_logic;
signal \n4814_cascade_\ : std_logic;
signal n5_adj_1235 : std_logic;
signal \n13475_cascade_\ : std_logic;
signal \n15802_cascade_\ : std_logic;
signal n10_adj_1249 : std_logic;
signal \n15657_cascade_\ : std_logic;
signal n13_adj_1042 : std_logic;
signal \comm_spi.n10479\ : std_logic;
signal \comm_spi.data_tx_7__N_806\ : std_logic;
signal n15576 : std_logic;
signal n15691 : std_logic;
signal n15475 : std_logic;
signal n15835 : std_logic;
signal n15542 : std_logic;
signal n15679 : std_logic;
signal n15543 : std_logic;
signal buf_adcdata3_17 : std_logic;
signal \M_DCSEL\ : std_logic;
signal \n90_adj_1023_cascade_\ : std_logic;
signal n69_adj_1113 : std_logic;
signal n96 : std_logic;
signal buf_device_acadc_4 : std_logic;
signal \M_OSR0\ : std_logic;
signal n15555 : std_logic;
signal \n3_cascade_\ : std_logic;
signal \n10_adj_1242_cascade_\ : std_logic;
signal n8_adj_1212 : std_logic;
signal eis_end : std_logic;
signal \INVeis_end_328C_net\ : std_logic;
signal \n15171_cascade_\ : std_logic;
signal \raw_buf1_N_775\ : std_logic;
signal n14087 : std_logic;
signal \n15356_cascade_\ : std_logic;
signal \n15695_cascade_\ : std_logic;
signal n15696 : std_logic;
signal \n15700_cascade_\ : std_logic;
signal n3 : std_logic;
signal \INVeis_state_i0C_net\ : std_logic;
signal n8459 : std_logic;
signal \data_index_9_N_258_4\ : std_logic;
signal \eis_end_N_773\ : std_logic;
signal \eis_end_N_773_cascade_\ : std_logic;
signal n15510 : std_logic;
signal n8_adj_1227 : std_logic;
signal cmd_rdadctmp_24_adj_1088 : std_logic;
signal \data_index_9_N_258_1\ : std_logic;
signal buf_data2_13 : std_logic;
signal buf_adcdata4_13 : std_logic;
signal n4059 : std_logic;
signal n8_adj_1233 : std_logic;
signal \n8_adj_1233_cascade_\ : std_logic;
signal \M_FLT0\ : std_logic;
signal n66_adj_1166 : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \INVacadc_skipcnt_i0_i0C_net\ : std_logic;
signal n13966 : std_logic;
signal \n13966_THRU_CRY_0_THRU_CO\ : std_logic;
signal \n13966_THRU_CRY_1_THRU_CO\ : std_logic;
signal \n13966_THRU_CRY_2_THRU_CO\ : std_logic;
signal \n13966_THRU_CRY_3_THRU_CO\ : std_logic;
signal \n13966_THRU_CRY_4_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n13966_THRU_CRY_5_THRU_CO\ : std_logic;
signal \n13966_THRU_CRY_6_THRU_CO\ : std_logic;
signal acadc_skipcnt_1 : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal n13967 : std_logic;
signal n13968 : std_logic;
signal acadc_skipcnt_4 : std_logic;
signal n13969 : std_logic;
signal n13970 : std_logic;
signal n13971 : std_logic;
signal n13972 : std_logic;
signal n13973 : std_logic;
signal n13974 : std_logic;
signal \INVacadc_skipcnt_i0_i1C_net\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal n13975 : std_logic;
signal n13976 : std_logic;
signal n13977 : std_logic;
signal n13978 : std_logic;
signal n13979 : std_logic;
signal n13980 : std_logic;
signal \INVacadc_skipcnt_i0_i9C_net\ : std_logic;
signal buf_data2_22 : std_logic;
signal buf_adcdata4_22 : std_logic;
signal n4102 : std_logic;
signal \comm_spi.n16902\ : std_logic;
signal \comm_spi.n10476\ : std_logic;
signal \comm_spi.n10480\ : std_logic;
signal \comm_spi.data_tx_7__N_816\ : std_logic;
signal \comm_spi.n10472\ : std_logic;
signal \comm_spi.n10471\ : std_logic;
signal \comm_spi.n10475\ : std_logic;
signal \comm_spi.data_tx_7__N_807\ : std_logic;
signal \comm_spi.n16896\ : std_logic;
signal n15474 : std_logic;
signal n15478 : std_logic;
signal n15680 : std_logic;
signal \INVcomm_spi.data_valid_85C_net\ : std_logic;
signal \comm_spi.n10449\ : std_logic;
signal \comm_spi.n10448\ : std_logic;
signal \INVcomm_spi.imiso_83_7340_7341_setC_net\ : std_logic;
signal n15387 : std_logic;
signal n15390 : std_logic;
signal \CLOCK_DDS.tmp_buf_10\ : std_logic;
signal \CLOCK_DDS.tmp_buf_11\ : std_logic;
signal \CLOCK_DDS.tmp_buf_12\ : std_logic;
signal \CLOCK_DDS.tmp_buf_13\ : std_logic;
signal \CLOCK_DDS.tmp_buf_14\ : std_logic;
signal buf_dds_9 : std_logic;
signal \CLOCK_DDS.tmp_buf_9\ : std_logic;
signal \CLOCK_DDS.tmp_buf_8\ : std_logic;
signal \n4260_cascade_\ : std_logic;
signal n15402 : std_logic;
signal \ICE_CHKCABLE\ : std_logic;
signal \n90_adj_1154_cascade_\ : std_logic;
signal n72 : std_logic;
signal \M_OSR1\ : std_logic;
signal n15479 : std_logic;
signal cmd_rdadctmp_31_adj_1081 : std_logic;
signal \n8_adj_1221_cascade_\ : std_logic;
signal n4205 : std_logic;
signal buf_device_acadc_7 : std_logic;
signal buf_dds_14 : std_logic;
signal n4219 : std_logic;
signal req_data_cnt_15 : std_logic;
signal req_data_cnt_9 : std_logic;
signal n22 : std_logic;
signal \n24_adj_1216_cascade_\ : std_logic;
signal n30_adj_1278 : std_logic;
signal \n6791_cascade_\ : std_logic;
signal \n8_adj_1178_cascade_\ : std_logic;
signal n7_adj_1177 : std_logic;
signal \n7_adj_1177_cascade_\ : std_logic;
signal n8_adj_1178 : std_logic;
signal \data_index_9_N_258_0\ : std_logic;
signal acadc_skipcnt_0 : std_logic;
signal acadc_skipcnt_6 : std_logic;
signal n18_adj_1276 : std_logic;
signal \n17_adj_1277_cascade_\ : std_logic;
signal n31 : std_logic;
signal \n31_cascade_\ : std_logic;
signal n15187 : std_logic;
signal n8_adj_1231 : std_logic;
signal \data_index_9_N_258_2\ : std_logic;
signal \M_FLT1\ : std_logic;
signal acadc_skipcnt_14 : std_logic;
signal acadc_skipcnt_11 : std_logic;
signal \acadc_skipCount_11\ : std_logic;
signal \n23_adj_1199_cascade_\ : std_logic;
signal n30 : std_logic;
signal acadc_skipcnt_10 : std_logic;
signal \acadc_skipCount_12\ : std_logic;
signal acadc_skipcnt_12 : std_logic;
signal n21 : std_logic;
signal data_index_0 : std_logic;
signal \data_index_9_N_647_0\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal data_index_1 : std_logic;
signal n7_adj_1232 : std_logic;
signal n14031 : std_logic;
signal data_index_2 : std_logic;
signal n7_adj_1230 : std_logic;
signal n14032 : std_logic;
signal n14033 : std_logic;
signal data_index_4 : std_logic;
signal n7_adj_1226 : std_logic;
signal n14034 : std_logic;
signal n14035 : std_logic;
signal n14036 : std_logic;
signal data_index_7 : std_logic;
signal n14037 : std_logic;
signal n14038 : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal data_index_3 : std_logic;
signal \M_DRDY2\ : std_logic;
signal n10532 : std_logic;
signal n15344 : std_logic;
signal n15171 : std_logic;
signal \n15328_cascade_\ : std_logic;
signal acadc_trig : std_logic;
signal \INVacadc_trig_329C_net\ : std_logic;
signal data_index_6 : std_logic;
signal n8_adj_1221 : std_logic;
signal n7_adj_1220 : std_logic;
signal \data_index_9_N_258_7\ : std_logic;
signal n7_adj_1222 : std_logic;
signal n8_adj_1223 : std_logic;
signal \data_index_9_N_258_6\ : std_logic;
signal \ICE_SPI_MISO\ : std_logic;
signal \comm_spi.n10446\ : std_logic;
signal \INVcomm_spi.MISO_48_7334_7335_resetC_net\ : std_logic;
signal \comm_spi.data_tx_7__N_813\ : std_logic;
signal comm_tx_buf_3 : std_logic;
signal \comm_spi.data_tx_7__N_825\ : std_logic;
signal buf_data1_22 : std_logic;
signal n66 : std_logic;
signal \comm_spi.n10452\ : std_logic;
signal \comm_spi.n10451\ : std_logic;
signal \comm_spi.n10444\ : std_logic;
signal \comm_spi.n10445\ : std_logic;
signal \INVcomm_spi.MISO_48_7334_7335_setC_net\ : std_logic;
signal \comm_spi.data_tx_7__N_805\ : std_logic;
signal n10640 : std_logic;
signal n15176 : std_logic;
signal n15396 : std_logic;
signal n15670 : std_logic;
signal n13475 : std_logic;
signal n15_adj_1203 : std_logic;
signal tmp_buf_15 : std_logic;
signal \CLOCK_DDS.tmp_buf_0\ : std_logic;
signal \CLOCK_DDS.tmp_buf_1\ : std_logic;
signal \CLOCK_DDS.tmp_buf_2\ : std_logic;
signal \CLOCK_DDS.tmp_buf_3\ : std_logic;
signal \CLOCK_DDS.tmp_buf_4\ : std_logic;
signal \CLOCK_DDS.tmp_buf_5\ : std_logic;
signal \CLOCK_DDS.tmp_buf_6\ : std_logic;
signal \CLOCK_DDS.tmp_buf_7\ : std_logic;
signal \CLOCK_DDS.n9759\ : std_logic;
signal n10823 : std_logic;
signal \CLOCK_DDS.n9_adj_1021\ : std_logic;
signal bit_cnt_1 : std_logic;
signal n15556 : std_logic;
signal n60_adj_1157 : std_logic;
signal n4252 : std_logic;
signal n4202 : std_logic;
signal n4247 : std_logic;
signal buf_dds_15 : std_logic;
signal req_data_cnt_13 : std_logic;
signal req_data_cnt_8 : std_logic;
signal n15812 : std_logic;
signal buf_device_acadc_6 : std_logic;
signal buf_data1_16 : std_logic;
signal n99 : std_logic;
signal req_data_cnt_7 : std_logic;
signal n4214 : std_logic;
signal buf_dds_7 : std_logic;
signal n7567 : std_logic;
signal n21_adj_1204 : std_logic;
signal comm_buf_1_4 : std_logic;
signal buf_dds_4 : std_logic;
signal buf_control_5 : std_logic;
signal buf_data1_10 : std_logic;
signal \n4195_cascade_\ : std_logic;
signal n4232 : std_logic;
signal acadc_skipcnt_9 : std_logic;
signal acadc_skipcnt_15 : std_logic;
signal n24_adj_1174 : std_logic;
signal req_data_cnt_14 : std_logic;
signal n23_adj_1194 : std_logic;
signal \acadc_skipCount_4\ : std_logic;
signal n9224 : std_logic;
signal buf_device_acadc_5 : std_logic;
signal \acadc_skipCount_9\ : std_logic;
signal n15834 : std_logic;
signal n19_adj_1234 : std_logic;
signal \n20_adj_1253_cascade_\ : std_logic;
signal n29 : std_logic;
signal n84 : std_logic;
signal n15546 : std_logic;
signal data_index_5 : std_logic;
signal buf_dds_12 : std_logic;
signal acadc_skipcnt_2 : std_logic;
signal \acadc_skipCount_7\ : std_logic;
signal acadc_skipcnt_7 : std_logic;
signal \acadc_skipCount_2\ : std_logic;
signal n22_adj_1170 : std_logic;
signal n8_adj_1229 : std_logic;
signal n7_adj_1228 : std_logic;
signal \data_index_9_N_258_3\ : std_logic;
signal n8456 : std_logic;
signal acadc_skipcnt_3 : std_logic;
signal acadc_skipcnt_5 : std_logic;
signal acadc_skipcnt_8 : std_logic;
signal \acadc_skipCount_8\ : std_logic;
signal \n20_cascade_\ : std_logic;
signal n26 : std_logic;
signal acadc_skipcnt_13 : std_logic;
signal \acadc_skipCount_13\ : std_logic;
signal n14_adj_1160 : std_logic;
signal cmd_rdadctmp_16 : std_logic;
signal buf_adcdata1_8 : std_logic;
signal eis_state_0 : std_logic;
signal \eis_end_N_770\ : std_logic;
signal \ICE_GPMO_0\ : std_logic;
signal data_index_8 : std_logic;
signal buf_data1_3 : std_logic;
signal buf_adcdata3_3 : std_logic;
signal n4149 : std_logic;
signal comm_tx_buf_5 : std_logic;
signal \comm_spi.data_tx_7__N_819\ : std_logic;
signal n8561 : std_logic;
signal \n15460_cascade_\ : std_logic;
signal \n19_cascade_\ : std_logic;
signal n15463 : std_logic;
signal n23 : std_logic;
signal \n19_adj_1151_cascade_\ : std_logic;
signal comm_length_2 : std_logic;
signal comm_index_2 : std_logic;
signal comm_length_3 : std_logic;
signal comm_index_3 : std_logic;
signal \n6_adj_1281_cascade_\ : std_logic;
signal comm_index_1 : std_logic;
signal n2 : std_logic;
signal \n15119_cascade_\ : std_logic;
signal comm_length_1 : std_logic;
signal \n13_cascade_\ : std_logic;
signal n6_adj_1273 : std_logic;
signal n5_adj_1282 : std_logic;
signal comm_length_0 : std_logic;
signal n10566 : std_logic;
signal n13 : std_logic;
signal n12649 : std_logic;
signal \n8525_cascade_\ : std_logic;
signal n4075 : std_logic;
signal n8133 : std_logic;
signal trig_dds : std_logic;
signal buf_dds_0 : std_logic;
signal buf_dds_8 : std_logic;
signal buf_data1_15 : std_logic;
signal \n4190_cascade_\ : std_logic;
signal n4227 : std_logic;
signal n4262 : std_logic;
signal comm_buf_0_5 : std_logic;
signal \n14_adj_1202_cascade_\ : std_logic;
signal buf_dds_13 : std_logic;
signal n15690 : std_logic;
signal req_data_cnt_12 : std_logic;
signal n13_adj_1026 : std_logic;
signal buf_data1_17 : std_logic;
signal \n78_cascade_\ : std_logic;
signal n99_adj_1024 : std_logic;
signal n4257 : std_logic;
signal comm_buf_1_6 : std_logic;
signal buf_data1_21 : std_logic;
signal n66_adj_1158 : std_logic;
signal buf_dds_5 : std_logic;
signal \acadc_skipCount_10\ : std_logic;
signal \n7485_cascade_\ : std_logic;
signal tacadc_rst : std_logic;
signal req_data_cnt_10 : std_logic;
signal n90_adj_1167 : std_logic;
signal n72_adj_1162 : std_logic;
signal comm_buf_0_0 : std_logic;
signal req_data_cnt_4 : std_logic;
signal n18_adj_1217 : std_logic;
signal buf_dds_6 : std_logic;
signal comm_buf_0_1 : std_logic;
signal n7485 : std_logic;
signal eis_stop : std_logic;
signal cmd_rdadctmp_23_adj_1053 : std_logic;
signal buf_adcdata2_15 : std_logic;
signal comm_buf_0_2 : std_logic;
signal buf_dds_10 : std_logic;
signal \acadc_skipCount_0\ : std_logic;
signal n17_adj_1214 : std_logic;
signal req_data_cnt_0 : std_logic;
signal \acadc_skipCount_6\ : std_logic;
signal buf_data1_14 : std_logic;
signal \n4191_cascade_\ : std_logic;
signal n4215 : std_logic;
signal \n4228_cascade_\ : std_logic;
signal n4203 : std_logic;
signal \n4248_cascade_\ : std_logic;
signal n4258 : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal n13951 : std_logic;
signal data_cntvec_2 : std_logic;
signal n13952 : std_logic;
signal n13953 : std_logic;
signal n13954 : std_logic;
signal n13955 : std_logic;
signal data_cntvec_6 : std_logic;
signal n13956 : std_logic;
signal data_cntvec_7 : std_logic;
signal n13957 : std_logic;
signal n13958 : std_logic;
signal \INVdata_cntvec_i0_i0C_net\ : std_logic;
signal data_cntvec_8 : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal data_cntvec_9 : std_logic;
signal n13959 : std_logic;
signal data_cntvec_10 : std_logic;
signal n13960 : std_logic;
signal data_cntvec_11 : std_logic;
signal n13961 : std_logic;
signal data_cntvec_12 : std_logic;
signal n13962 : std_logic;
signal data_cntvec_13 : std_logic;
signal n13963 : std_logic;
signal data_cntvec_14 : std_logic;
signal n13964 : std_logic;
signal n13965 : std_logic;
signal data_cntvec_15 : std_logic;
signal \INVdata_cntvec_i0_i8C_net\ : std_logic;
signal data_count_0 : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal data_count_1 : std_logic;
signal n13942 : std_logic;
signal data_count_2 : std_logic;
signal n13943 : std_logic;
signal data_count_3 : std_logic;
signal n13944 : std_logic;
signal data_count_4 : std_logic;
signal n13945 : std_logic;
signal data_count_5 : std_logic;
signal n13946 : std_logic;
signal data_count_6 : std_logic;
signal n13947 : std_logic;
signal data_count_7 : std_logic;
signal n13948 : std_logic;
signal n13949 : std_logic;
signal \INVdata_count_i0_i0C_net\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal data_count_8 : std_logic;
signal \INVdata_count_i0_i8C_net\ : std_logic;
signal dds_state_2 : std_logic;
signal \ADC_VAC2.n15280\ : std_logic;
signal adc_state_1_adj_1043 : std_logic;
signal \ADC_VAC2.n12\ : std_logic;
signal \ADC_VAC2.n14926\ : std_logic;
signal \ADC_VAC2.n9413\ : std_logic;
signal \DTRIG_N_957_adj_1077\ : std_logic;
signal \ADC_VAC2.n10706\ : std_logic;
signal \comm_spi.bit_cnt_2\ : std_logic;
signal \comm_spi.bit_cnt_1\ : std_logic;
signal \comm_spi.bit_cnt_0\ : std_logic;
signal \INVcomm_spi.bit_cnt_1603__i3C_net\ : std_logic;
signal \n15668_cascade_\ : std_logic;
signal n1523 : std_logic;
signal \n1523_cascade_\ : std_logic;
signal \n2_adj_1200_cascade_\ : std_logic;
signal n16464 : std_logic;
signal \n16467_cascade_\ : std_logic;
signal n8_adj_1201 : std_logic;
signal n15527 : std_logic;
signal n14_adj_1189 : std_logic;
signal n13_adj_1032 : std_logic;
signal \n13_adj_1032_cascade_\ : std_logic;
signal n8519 : std_logic;
signal n22_adj_1115 : std_logic;
signal n15651 : std_logic;
signal n15526 : std_logic;
signal buf_data1_20 : std_logic;
signal \n8058_cascade_\ : std_logic;
signal comm_buf_0_4 : std_logic;
signal n15584 : std_logic;
signal \n83_cascade_\ : std_logic;
signal n15581 : std_logic;
signal cmd_rdadctmp_29_adj_1083 : std_logic;
signal buf_adcdata3_21 : std_logic;
signal cmd_rdadctmp_23_adj_1089 : std_logic;
signal buf_adcdata3_15 : std_logic;
signal buf_data1_18 : std_logic;
signal n75_adj_1164 : std_logic;
signal comm_buf_1_0 : std_logic;
signal data_cntvec_0 : std_logic;
signal buf_data1_8 : std_logic;
signal \n4197_cascade_\ : std_logic;
signal n4221 : std_logic;
signal \n4234_cascade_\ : std_logic;
signal n4209 : std_logic;
signal \n4254_cascade_\ : std_logic;
signal n4264 : std_logic;
signal \n32_cascade_\ : std_logic;
signal n15557 : std_logic;
signal data_idxvec_0 : std_logic;
signal \data_idxvec_15_N_673_0\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal n14040 : std_logic;
signal data_idxvec_2 : std_logic;
signal n14041 : std_logic;
signal n14042 : std_logic;
signal n14_adj_1196 : std_logic;
signal n14043 : std_logic;
signal n14_adj_1213 : std_logic;
signal n14044 : std_logic;
signal data_idxvec_6 : std_logic;
signal n14045 : std_logic;
signal n14_adj_1168 : std_logic;
signal data_idxvec_7 : std_logic;
signal n14046 : std_logic;
signal n14047 : std_logic;
signal n14_adj_1211 : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal n14_adj_1210 : std_logic;
signal data_idxvec_9 : std_logic;
signal n14048 : std_logic;
signal n14_adj_1209 : std_logic;
signal data_idxvec_10 : std_logic;
signal n14049 : std_logic;
signal n14050 : std_logic;
signal n14_adj_1207 : std_logic;
signal data_idxvec_12 : std_logic;
signal n14051 : std_logic;
signal n14_adj_1202 : std_logic;
signal data_idxvec_13 : std_logic;
signal n14052 : std_logic;
signal n14_adj_1206 : std_logic;
signal data_idxvec_14 : std_logic;
signal n14053 : std_logic;
signal n14_adj_1205 : std_logic;
signal n14054 : std_logic;
signal n9187 : std_logic;
signal buf_adcdata3_13 : std_logic;
signal n14_adj_1198 : std_logic;
signal cmd_rdadctmp_22 : std_logic;
signal buf_adcdata1_14 : std_logic;
signal req_data_cnt_11 : std_logic;
signal n14_adj_1169 : std_logic;
signal req_data_cnt_6 : std_logic;
signal n4204 : std_logic;
signal \n4249_cascade_\ : std_logic;
signal \n4259_cascade_\ : std_logic;
signal comm_buf_1_5 : std_logic;
signal data_idxvec_4 : std_logic;
signal data_cntvec_4 : std_logic;
signal buf_data1_12 : std_logic;
signal \n4193_cascade_\ : std_logic;
signal req_data_cnt_5 : std_logic;
signal \acadc_skipCount_5\ : std_logic;
signal n4216 : std_logic;
signal data_idxvec_5 : std_logic;
signal data_cntvec_5 : std_logic;
signal buf_data1_13 : std_logic;
signal \n4192_cascade_\ : std_logic;
signal n4229 : std_logic;
signal cmd_rdadctmp_18_adj_1058 : std_logic;
signal buf_adcdata2_10 : std_logic;
signal data_idxvec_1 : std_logic;
signal data_cntvec_1 : std_logic;
signal cmd_rdadctmp_16_adj_1096 : std_logic;
signal req_data_cnt_3 : std_logic;
signal \acadc_skipCount_3\ : std_logic;
signal eis_state_1 : std_logic;
signal n9790 : std_logic;
signal n10483 : std_logic;
signal \comm_spi.n16887\ : std_logic;
signal \comm_spi.n10438\ : std_logic;
signal \comm_spi.iclk_N_802\ : std_logic;
signal \comm_spi.n16890\ : std_logic;
signal \comm_spi.n10455\ : std_logic;
signal \comm_spi.n16890_cascade_\ : std_logic;
signal \comm_spi.bit_cnt_3\ : std_logic;
signal \comm_spi.n12175\ : std_logic;
signal comm_buf_1_7 : std_logic;
signal comm_buf_0_7 : std_logic;
signal comm_index_0 : std_logic;
signal n15381 : std_logic;
signal \n12846_cascade_\ : std_logic;
signal n4_adj_1179 : std_logic;
signal n15204 : std_logic;
signal \n4_adj_1184_cascade_\ : std_logic;
signal n15290 : std_logic;
signal \n15241_cascade_\ : std_logic;
signal n15108 : std_logic;
signal n15128 : std_logic;
signal n8530 : std_logic;
signal n15198 : std_logic;
signal n15266 : std_logic;
signal \n15410_cascade_\ : std_logic;
signal n15130 : std_logic;
signal n15408 : std_logic;
signal n10394 : std_logic;
signal n16190 : std_logic;
signal n15635 : std_logic;
signal n12_adj_1027 : std_logic;
signal n12622 : std_logic;
signal n14_adj_1152 : std_logic;
signal n93 : std_logic;
signal n27 : std_logic;
signal n4 : std_logic;
signal \n15309_cascade_\ : std_logic;
signal \comm_state_3_N_402_3\ : std_logic;
signal n15637 : std_logic;
signal n13_adj_1040 : std_logic;
signal n22_adj_1078 : std_logic;
signal comm_rx_buf_7 : std_logic;
signal comm_cmd_7 : std_logic;
signal comm_rx_buf_0 : std_logic;
signal comm_rx_buf_2 : std_logic;
signal comm_buf_1_2 : std_logic;
signal comm_rx_buf_4 : std_logic;
signal \n10363_cascade_\ : std_logic;
signal comm_rx_buf_5 : std_logic;
signal n8062 : std_logic;
signal \n8085_cascade_\ : std_logic;
signal n24 : std_logic;
signal comm_rx_buf_6 : std_logic;
signal buf_data1_19 : std_logic;
signal data_idxvec_11 : std_logic;
signal n75 : std_logic;
signal \n12_cascade_\ : std_logic;
signal n6301 : std_logic;
signal n8253 : std_logic;
signal n14_adj_1197 : std_logic;
signal req_data_cnt_2 : std_logic;
signal comm_cmd_5 : std_logic;
signal comm_cmd_4 : std_logic;
signal comm_cmd_6 : std_logic;
signal n8043 : std_logic;
signal n7511 : std_logic;
signal comm_buf_1_1 : std_logic;
signal eis_start : std_logic;
signal data_idxvec_8 : std_logic;
signal n78_adj_1022 : std_logic;
signal buf_dds_3 : std_logic;
signal n8 : std_logic;
signal n15188 : std_logic;
signal n12702 : std_logic;
signal \n15188_cascade_\ : std_logic;
signal n8085 : std_logic;
signal \n6_adj_1171_cascade_\ : std_logic;
signal n15190 : std_logic;
signal buf_adcdata3_12 : std_logic;
signal cmd_rdadctmp_21_adj_1091 : std_logic;
signal n4_adj_1041 : std_logic;
signal comm_buf_0_6 : std_logic;
signal n8250 : std_logic;
signal \acadc_skipCount_14\ : std_logic;
signal data_idxvec_15 : std_logic;
signal \acadc_skipCount_15\ : std_logic;
signal n15468 : std_logic;
signal n4217 : std_logic;
signal n4230 : std_logic;
signal n4250 : std_logic;
signal cmd_rdadctmp_22_adj_1090 : std_logic;
signal buf_adcdata3_14 : std_logic;
signal n1 : std_logic;
signal n8525 : std_logic;
signal buf_dds_11 : std_logic;
signal n12 : std_logic;
signal n13_adj_1025 : std_logic;
signal \acadc_skipCount_1\ : std_logic;
signal req_data_cnt_1 : std_logic;
signal \n4220_cascade_\ : std_logic;
signal \n4253_cascade_\ : std_logic;
signal n4263 : std_logic;
signal buf_dds_1 : std_logic;
signal buf_adcdata3_9 : std_logic;
signal n4208 : std_logic;
signal buf_data1_9 : std_logic;
signal n4196 : std_logic;
signal n4233 : std_logic;
signal data_idxvec_3 : std_logic;
signal data_cntvec_3 : std_logic;
signal buf_data1_11 : std_logic;
signal \n4194_cascade_\ : std_logic;
signal n4218 : std_logic;
signal \n4231_cascade_\ : std_logic;
signal n4206 : std_logic;
signal \n4251_cascade_\ : std_logic;
signal buf_data2_9 : std_logic;
signal buf_adcdata4_9 : std_logic;
signal n4063 : std_logic;
signal buf_adcdata2_11 : std_logic;
signal n8_adj_1219 : std_logic;
signal n7_adj_1218 : std_logic;
signal \data_index_9_N_258_8\ : std_logic;
signal \comm_spi.n10456\ : std_logic;
signal \comm_spi.iclk\ : std_logic;
signal \comm_spi.n16893\ : std_logic;
signal \comm_spi.n10441\ : std_logic;
signal \comm_spi.n16893_cascade_\ : std_logic;
signal \comm_spi.imosi_cascade_\ : std_logic;
signal \comm_spi.DOUT_7__N_785\ : std_logic;
signal \comm_spi.imosi_N_791\ : std_logic;
signal cmd_rdadctmp_9_adj_1067 : std_logic;
signal buf_adcdata2_1 : std_logic;
signal \comm_spi.imosi\ : std_logic;
signal \comm_spi.DOUT_7__N_786\ : std_logic;
signal n15131 : std_logic;
signal n15241 : std_logic;
signal n15191 : std_logic;
signal n10148 : std_logic;
signal n7 : std_logic;
signal \comm_state_3_N_418_1\ : std_logic;
signal \n15711_cascade_\ : std_logic;
signal n8_adj_1193 : std_logic;
signal \n26_adj_1192_cascade_\ : std_logic;
signal n18_adj_1191 : std_logic;
signal n15245 : std_logic;
signal \ICE_SPI_CE0\ : std_logic;
signal \n15245_cascade_\ : std_logic;
signal comm_data_vld : std_logic;
signal n8544 : std_logic;
signal n9_adj_1028 : std_logic;
signal n9011 : std_logic;
signal \n9011_cascade_\ : std_logic;
signal n9215 : std_logic;
signal buf_data2_19 : std_logic;
signal buf_adcdata4_19 : std_logic;
signal \comm_buf_3_7_N_501_3\ : std_logic;
signal buf_control_6 : std_logic;
signal n60 : std_logic;
signal cmd_rdadctmp_8_adj_1104 : std_logic;
signal buf_adcdata3_0 : std_logic;
signal buf_adcdata3_11 : std_logic;
signal cmd_rdadctmp_30_adj_1082 : std_logic;
signal buf_adcdata3_22 : std_logic;
signal n7_adj_1190 : std_logic;
signal buf_dds_2 : std_logic;
signal n4207 : std_logic;
signal n8094 : std_logic;
signal n729 : std_logic;
signal buf_adcdata2_19 : std_logic;
signal comm_buf_0_3 : std_logic;
signal n14_adj_1208 : std_logic;
signal cmd_rdadctmp_10 : std_logic;
signal buf_adcdata1_2 : std_logic;
signal n15147 : std_logic;
signal buf_adcdata3_10 : std_logic;
signal comm_rx_buf_1 : std_logic;
signal n8618 : std_logic;
signal n10363 : std_logic;
signal cmd_rdadctmp_25_adj_1051 : std_logic;
signal buf_adcdata2_18 : std_logic;
signal n14_adj_1215 : std_logic;
signal cmd_rdadctmp_26_adj_1050 : std_logic;
signal cmd_rdadctmp_27_adj_1049 : std_logic;
signal n4_adj_1250 : std_logic;
signal buf_adcdata2_12 : std_logic;
signal comm_cmd_2 : std_logic;
signal comm_cmd_1 : std_logic;
signal n9 : std_logic;
signal comm_rx_buf_3 : std_logic;
signal n4261 : std_logic;
signal comm_buf_1_3 : std_logic;
signal n8702 : std_logic;
signal n10583 : std_logic;
signal cmd_rdadctmp_21 : std_logic;
signal buf_adcdata1_13 : std_logic;
signal cmd_rdadctmp_17_adj_1095 : std_logic;
signal cmd_rdadctmp_18_adj_1094 : std_logic;
signal buf_adcdata2_13 : std_logic;
signal cmd_rdadctmp_20 : std_logic;
signal buf_adcdata1_12 : std_logic;
signal cmd_rdadctmp_17_adj_1059 : std_logic;
signal buf_adcdata2_9 : std_logic;
signal cmd_rdadctmp_19_adj_1057 : std_logic;
signal cmd_rdadctmp_20_adj_1056 : std_logic;
signal n8302 : std_logic;
signal cmd_rdadctmp_21_adj_1055 : std_logic;
signal buf_data2_23 : std_logic;
signal buf_adcdata4_23 : std_logic;
signal n4101 : std_logic;
signal \comm_spi.n10442\ : std_logic;
signal \ICE_SPI_MOSI\ : std_logic;
signal \comm_spi.imosi_N_792\ : std_logic;
signal cmd_rdadctmp_28_adj_1048 : std_logic;
signal buf_adcdata2_20 : std_logic;
signal cmd_rdadctmp_31_adj_1045 : std_logic;
signal buf_adcdata2_23 : std_logic;
signal buf_data2_16 : std_logic;
signal comm_cmd_0 : std_logic;
signal buf_adcdata4_16 : std_logic;
signal comm_cmd_3 : std_logic;
signal n4108 : std_logic;
signal cmd_rdadctmp_10_adj_1066 : std_logic;
signal buf_adcdata2_2 : std_logic;
signal \comm_spi.data_tx_7__N_808\ : std_logic;
signal comm_tx_buf_4 : std_logic;
signal comm_clear : std_logic;
signal \comm_spi.n16899\ : std_logic;
signal cmd_rdadctmp_29_adj_1047 : std_logic;
signal buf_adcdata2_21 : std_logic;
signal \ICE_GPMI_0\ : std_logic;
signal n8576 : std_logic;
signal n8117 : std_logic;
signal n6_adj_1175 : std_logic;
signal comm_state_0 : std_logic;
signal comm_state_1 : std_logic;
signal comm_state_2 : std_logic;
signal n8129 : std_logic;
signal cmd_rdadctmp_19_adj_1093 : std_logic;
signal adc_state_0_adj_1080 : std_logic;
signal n8332 : std_logic;
signal cmd_rdadctmp_20_adj_1092 : std_logic;
signal n15640 : std_logic;
signal n10_adj_1172 : std_logic;
signal dds_state_1 : std_logic;
signal dds_state_0 : std_logic;
signal \CLOCK_DDS.n9\ : std_logic;
signal cmd_rdadctmp_24 : std_logic;
signal buf_adcdata1_16 : std_logic;
signal cmd_rdadctmp_30_adj_1046 : std_logic;
signal buf_adcdata2_22 : std_logic;
signal n15150 : std_logic;
signal cmd_rdadctmp_22_adj_1054 : std_logic;
signal adc_state_0_adj_1044 : std_logic;
signal buf_adcdata2_14 : std_logic;
signal n15153 : std_logic;
signal cmd_rdadctmp_18 : std_logic;
signal adc_state_0 : std_logic;
signal buf_adcdata1_10 : std_logic;
signal n8_adj_1225 : std_logic;
signal comm_state_3 : std_logic;
signal n6791 : std_logic;
signal n7_adj_1224 : std_logic;
signal \data_index_9_N_258_5\ : std_logic;
signal \ICE_SPI_SCLK\ : std_logic;
signal \comm_spi.n10437\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \clk_32MHz\ : std_logic;
signal \comm_spi.iclk_N_801\ : std_logic;

signal \M_CS1_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \M_MOSI1_wire\ : std_logic;
signal \M_DRDY1_wire\ : std_logic;
signal \M_CLK2_wire\ : std_logic;
signal \M_SCLK1_wire\ : std_logic;
signal \M_FLT0_wire\ : std_logic;
signal \M_CS3_wire\ : std_logic;
signal \ICE_CHKCABLE_wire\ : std_logic;
signal \M_OSR1_wire\ : std_logic;
signal \ICE_GPMO_1_wire\ : std_logic;
signal \EIS_SYNCCLK_wire\ : std_logic;
signal \M_SCLK3_wire\ : std_logic;
signal \M_OSR0_wire\ : std_logic;
signal \M_MISO4_wire\ : std_logic;
signal \M_DRDY4_wire\ : std_logic;
signal \ICE_SPI_MOSI_wire\ : std_logic;
signal \ICE_GPMO_0_wire\ : std_logic;
signal \DDS_MOSI1_wire\ : std_logic;
signal \M_SCLK4_wire\ : std_logic;
signal \M_MISO3_wire\ : std_logic;
signal \M_CS4_wire\ : std_logic;
signal \ICE_SPI_SCLK_wire\ : std_logic;
signal \M_MOSI4_wire\ : std_logic;
signal \M_MISO2_wire\ : std_logic;
signal \M_DRDY2_wire\ : std_logic;
signal \M_CLK1_wire\ : std_logic;
signal \ICE_SPI_MISO_wire\ : std_logic;
signal \ICE_GPMO_2_wire\ : std_logic;
signal \ICE_GPMI_0_wire\ : std_logic;
signal \TEST_LED_wire\ : std_logic;
signal \M_POW_wire\ : std_logic;
signal \M_MOSI3_wire\ : std_logic;
signal \M_MISO1_wire\ : std_logic;
signal \M_DRDY3_wire\ : std_logic;
signal \M_DCSEL_wire\ : std_logic;
signal \M_START_wire\ : std_logic;
signal \M_MOSI2_wire\ : std_logic;
signal \M_CLK3_wire\ : std_logic;
signal \DDS_CS1_wire\ : std_logic;
signal \M_FLT1_wire\ : std_logic;
signal \DISP_COMM_wire\ : std_logic;
signal \DDS_MCLK1_wire\ : std_logic;
signal \ICE_SPI_CE0_wire\ : std_logic;
signal \M_SCLK2_wire\ : std_logic;
signal \M_CS2_wire\ : std_logic;
signal \M_CLK4_wire\ : std_logic;
signal \DDS_SCK1_wire\ : std_logic;
signal \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    M_CS1 <= \M_CS1_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    M_MOSI1 <= \M_MOSI1_wire\;
    \M_DRDY1_wire\ <= M_DRDY1;
    M_CLK2 <= \M_CLK2_wire\;
    M_SCLK1 <= \M_SCLK1_wire\;
    M_FLT0 <= \M_FLT0_wire\;
    M_CS3 <= \M_CS3_wire\;
    \ICE_CHKCABLE_wire\ <= ICE_CHKCABLE;
    M_OSR1 <= \M_OSR1_wire\;
    \ICE_GPMO_1_wire\ <= ICE_GPMO_1;
    \EIS_SYNCCLK_wire\ <= EIS_SYNCCLK;
    M_SCLK3 <= \M_SCLK3_wire\;
    M_OSR0 <= \M_OSR0_wire\;
    \M_MISO4_wire\ <= M_MISO4;
    \M_DRDY4_wire\ <= M_DRDY4;
    \ICE_SPI_MOSI_wire\ <= ICE_SPI_MOSI;
    \ICE_GPMO_0_wire\ <= ICE_GPMO_0;
    DDS_MOSI1 <= \DDS_MOSI1_wire\;
    M_SCLK4 <= \M_SCLK4_wire\;
    \M_MISO3_wire\ <= M_MISO3;
    M_CS4 <= \M_CS4_wire\;
    \ICE_SPI_SCLK_wire\ <= ICE_SPI_SCLK;
    M_MOSI4 <= \M_MOSI4_wire\;
    \M_MISO2_wire\ <= M_MISO2;
    \M_DRDY2_wire\ <= M_DRDY2;
    M_CLK1 <= \M_CLK1_wire\;
    ICE_SPI_MISO <= \ICE_SPI_MISO_wire\;
    \ICE_GPMO_2_wire\ <= ICE_GPMO_2;
    ICE_GPMI_0 <= \ICE_GPMI_0_wire\;
    TEST_LED <= \TEST_LED_wire\;
    M_POW <= \M_POW_wire\;
    M_MOSI3 <= \M_MOSI3_wire\;
    \M_MISO1_wire\ <= M_MISO1;
    \M_DRDY3_wire\ <= M_DRDY3;
    M_DCSEL <= \M_DCSEL_wire\;
    M_START <= \M_START_wire\;
    M_MOSI2 <= \M_MOSI2_wire\;
    M_CLK3 <= \M_CLK3_wire\;
    DDS_CS1 <= \DDS_CS1_wire\;
    M_FLT1 <= \M_FLT1_wire\;
    DISP_COMM <= \DISP_COMM_wire\;
    DDS_MCLK1 <= \DDS_MCLK1_wire\;
    \ICE_SPI_CE0_wire\ <= ICE_SPI_CE0;
    M_SCLK2 <= \M_SCLK2_wire\;
    M_CS2 <= \M_CS2_wire\;
    M_CLK4 <= \M_CLK4_wire\;
    DDS_SCK1 <= \DDS_SCK1_wire\;
    \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    buf_data1_19 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(14);
    buf_data4_19 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(12);
    buf_data3_19 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(10);
    buf_data2_19 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(8);
    buf_data1_18 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(6);
    buf_data4_18 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(4);
    buf_data3_18 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(2);
    buf_data2_18 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RADDR_wire\ <= '0'&'0'&\N__42539\&\N__30500\&\N__30356\&\N__51470\&\N__28157\&\N__32453\&\N__29660\&\N__28442\&\N__29840\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_WADDR_wire\ <= '0'&'0'&\N__35843\&\N__35951\&\N__36059\&\N__36167\&\N__36278\&\N__35039\&\N__35144\&\N__35249\&\N__35354\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_WDATA_wire\ <= '0'&\N__20237\&'0'&\N__43031\&'0'&\N__26225\&'0'&\N__43580\&'0'&\N__20042\&'0'&\N__19295\&'0'&\N__26465\&'0'&\N__43937\;
    buf_data1_17 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(14);
    buf_data4_17 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(12);
    buf_data3_17 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(10);
    buf_data2_17 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(8);
    buf_data1_16 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(6);
    buf_data4_16 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(4);
    buf_data3_16 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(2);
    buf_data2_16 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RADDR_wire\ <= '0'&'0'&\N__42533\&\N__30494\&\N__30350\&\N__51464\&\N__28151\&\N__32447\&\N__29654\&\N__28436\&\N__29834\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_WADDR_wire\ <= '0'&'0'&\N__35837\&\N__35945\&\N__36053\&\N__36161\&\N__36272\&\N__35033\&\N__35138\&\N__35243\&\N__35348\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_WDATA_wire\ <= '0'&\N__20069\&'0'&\N__25798\&'0'&\N__27959\&'0'&\N__20354\&'0'&\N__48227\&'0'&\N__47371\&'0'&\N__26363\&'0'&\N__21308\;
    buf_data1_7 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(14);
    buf_data4_7 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(12);
    buf_data3_7 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(10);
    buf_data2_7 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(8);
    buf_data1_6 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(6);
    buf_data4_6 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(4);
    buf_data3_6 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(2);
    buf_data2_6 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RADDR_wire\ <= '0'&'0'&\N__42523\&\N__30481\&\N__30340\&\N__51460\&\N__28141\&\N__32440\&\N__29641\&\N__28426\&\N__29821\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_WADDR_wire\ <= '0'&'0'&\N__35821\&\N__35929\&\N__36040\&\N__36148\&\N__36262\&\N__35020\&\N__35122\&\N__35227\&\N__35332\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_WDATA_wire\ <= '0'&\N__17774\&'0'&\N__17474\&'0'&\N__18719\&'0'&\N__17618\&'0'&\N__21707\&'0'&\N__17680\&'0'&\N__19529\&'0'&\N__17639\;
    buf_data1_15 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(14);
    buf_data4_15 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(12);
    buf_data3_15 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(10);
    buf_data2_15 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(8);
    buf_data1_14 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(6);
    buf_data4_14 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(4);
    buf_data3_14 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(2);
    buf_data2_14 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RADDR_wire\ <= '0'&'0'&\N__42527\&\N__30488\&\N__30344\&\N__51457\&\N__28145\&\N__32441\&\N__29648\&\N__28430\&\N__29828\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_WADDR_wire\ <= '0'&'0'&\N__35831\&\N__35939\&\N__36047\&\N__36155\&\N__36266\&\N__35027\&\N__35132\&\N__35237\&\N__35342\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_WDATA_wire\ <= '0'&\N__22688\&'0'&\N__26002\&'0'&\N__36770\&'0'&\N__34445\&'0'&\N__37445\&'0'&\N__24107\&'0'&\N__41558\&'0'&\N__53144\;
    buf_data1_5 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(14);
    buf_data4_5 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(12);
    buf_data3_5 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(10);
    buf_data2_5 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(8);
    buf_data1_4 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(6);
    buf_data4_4 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(4);
    buf_data3_4 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(2);
    buf_data2_4 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RADDR_wire\ <= '0'&'0'&\N__42511\&\N__30469\&\N__30328\&\N__51448\&\N__28129\&\N__32428\&\N__29629\&\N__28414\&\N__29809\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_WADDR_wire\ <= '0'&'0'&\N__35809\&\N__35917\&\N__36028\&\N__36136\&\N__36250\&\N__35008\&\N__35110\&\N__35215\&\N__35320\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_WDATA_wire\ <= '0'&\N__17792\&'0'&\N__17752\&'0'&\N__19564\&'0'&\N__17657\&'0'&\N__18635\&'0'&\N__18125\&'0'&\N__18760\&'0'&\N__17885\;
    buf_data1_1 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(14);
    buf_data4_1 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(12);
    buf_data3_1 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(10);
    buf_data2_1 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(8);
    buf_data1_0 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(6);
    buf_data4_0 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(4);
    buf_data3_0 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(2);
    buf_data2_0 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RADDR_wire\ <= '0'&'0'&\N__42545\&\N__30506\&\N__30362\&\N__51476\&\N__28163\&\N__32459\&\N__29666\&\N__28448\&\N__29846\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_WADDR_wire\ <= '0'&'0'&\N__35849\&\N__35957\&\N__36065\&\N__36173\&\N__36284\&\N__35045\&\N__35150\&\N__35255\&\N__35360\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_WDATA_wire\ <= '0'&\N__21260\&'0'&\N__17993\&'0'&\N__27593\&'0'&\N__42908\&'0'&\N__22451\&'0'&\N__18029\&'0'&\N__43810\&'0'&\N__17225\;
    buf_data1_13 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(14);
    buf_data4_13 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(12);
    buf_data3_13 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(10);
    buf_data2_13 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(8);
    buf_data1_12 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(6);
    buf_data4_12 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(4);
    buf_data3_12 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(2);
    buf_data2_12 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RADDR_wire\ <= '0'&'0'&\N__42520\&\N__30482\&\N__30337\&\N__51445\&\N__28138\&\N__32431\&\N__29642\&\N__28423\&\N__29822\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_WADDR_wire\ <= '0'&'0'&\N__35825\&\N__35933\&\N__36041\&\N__36149\&\N__36259\&\N__35021\&\N__35126\&\N__35231\&\N__35336\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_WDATA_wire\ <= '0'&\N__44563\&'0'&\N__28615\&'0'&\N__37520\&'0'&\N__44486\&'0'&\N__46256\&'0'&\N__20495\&'0'&\N__40783\&'0'&\N__45680\;
    buf_data1_23 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(14);
    buf_data4_23 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(12);
    buf_data3_23 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(10);
    buf_data2_23 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(8);
    buf_data1_22 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(6);
    buf_data4_22 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(4);
    buf_data3_22 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(2);
    buf_data2_22 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RADDR_wire\ <= '0'&'0'&\N__42563\&\N__30524\&\N__30380\&\N__51494\&\N__28181\&\N__32477\&\N__29684\&\N__28466\&\N__29864\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_WADDR_wire\ <= '0'&'0'&\N__35867\&\N__35975\&\N__36083\&\N__36191\&\N__36302\&\N__35063\&\N__35168\&\N__35273\&\N__35378\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_WDATA_wire\ <= '0'&\N__22736\&'0'&\N__45878\&'0'&\N__25685\&'0'&\N__48122\&'0'&\N__21365\&'0'&\N__29078\&'0'&\N__43718\&'0'&\N__48179\;
    buf_data1_3 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(14);
    buf_data4_3 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(12);
    buf_data3_3 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(10);
    buf_data2_3 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(8);
    buf_data1_2 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(6);
    buf_data4_2 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(4);
    buf_data3_2 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(2);
    buf_data2_2 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RADDR_wire\ <= '0'&'0'&\N__42551\&\N__30512\&\N__30368\&\N__51482\&\N__28169\&\N__32465\&\N__29672\&\N__28454\&\N__29852\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_WADDR_wire\ <= '0'&'0'&\N__35855\&\N__35963\&\N__36071\&\N__36179\&\N__36290\&\N__35051\&\N__35156\&\N__35261\&\N__35366\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_WDATA_wire\ <= '0'&\N__18785\&'0'&\N__20819\&'0'&\N__32624\&'0'&\N__17582\&'0'&\N__44426\&'0'&\N__17921\&'0'&\N__18482\&'0'&\N__46666\;
    buf_data1_11 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(14);
    buf_data4_11 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(12);
    buf_data3_11 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(10);
    buf_data2_11 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(8);
    buf_data1_10 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(6);
    buf_data4_10 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(4);
    buf_data3_10 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(2);
    buf_data2_10 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RADDR_wire\ <= '0'&'0'&\N__42508\&\N__30472\&\N__30325\&\N__51433\&\N__28126\&\N__32419\&\N__29632\&\N__28411\&\N__29812\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_WADDR_wire\ <= '0'&'0'&\N__35818\&\N__35926\&\N__36031\&\N__36139\&\N__36247\&\N__35011\&\N__35119\&\N__35224\&\N__35329\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_WDATA_wire\ <= '0'&\N__24539\&'0'&\N__26552\&'0'&\N__43778\&'0'&\N__42620\&'0'&\N__52505\&'0'&\N__19708\&'0'&\N__44207\&'0'&\N__38261\;
    buf_data1_21 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(14);
    buf_data4_21 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(12);
    buf_data3_21 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(10);
    buf_data2_21 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(8);
    buf_data1_20 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(6);
    buf_data4_20 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(4);
    buf_data3_20 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(2);
    buf_data2_20 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RADDR_wire\ <= '0'&'0'&\N__42557\&\N__30518\&\N__30374\&\N__51488\&\N__28175\&\N__32471\&\N__29678\&\N__28460\&\N__29858\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_WADDR_wire\ <= '0'&'0'&\N__35861\&\N__35969\&\N__36077\&\N__36185\&\N__36296\&\N__35057\&\N__35162\&\N__35267\&\N__35372\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_WDATA_wire\ <= '0'&\N__21167\&'0'&\N__23173\&'0'&\N__36845\&'0'&\N__46331\&'0'&\N__20189\&'0'&\N__24653\&'0'&\N__24073\&'0'&\N__45707\;
    buf_data1_9 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(14);
    buf_data4_9 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(12);
    buf_data3_9 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(10);
    buf_data2_9 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(8);
    buf_data1_8 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(6);
    buf_data4_8 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(4);
    buf_data3_8 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(2);
    buf_data2_8 <= \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\(0);
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RADDR_wire\ <= '0'&'0'&\N__42496\&\N__30460\&\N__30313\&\N__51421\&\N__28114\&\N__32407\&\N__29620\&\N__28399\&\N__29800\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_WADDR_wire\ <= '0'&'0'&\N__35806\&\N__35914\&\N__36019\&\N__36127\&\N__36235\&\N__34999\&\N__35107\&\N__35212\&\N__35317\;
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_WDATA_wire\ <= '0'&\N__24602\&'0'&\N__42670\&'0'&\N__42095\&'0'&\N__46202\&'0'&\N__32147\&'0'&\N__24350\&'0'&\N__24511\&'0'&\N__20420\;

    \pll_main.zim_pll_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => OPEN,
            REFERENCECLK => \N__16769\,
            RESETB => \N__28782\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => \clk_16MHz\,
            DYNAMICDELAY => \pll_main.zim_pll_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \clk_32MHz\,
            SCLK => \GNDG0\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51259\,
            RE => \N__28823\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN_net\,
            WE => \N__28346\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51287\,
            RE => \N__28837\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN_net\,
            WE => \N__28272\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51174\,
            RE => \N__28802\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN_net\,
            WE => \N__28345\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51305\,
            RE => \N__28838\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN_net\,
            WE => \N__28322\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51209\,
            RE => \N__28821\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN_net\,
            WE => \N__28344\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51226\,
            RE => \N__28822\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN_net\,
            WE => \N__28340\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51313\,
            RE => \N__28848\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN_net\,
            WE => \N__28353\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51134\,
            RE => \N__28774\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN_net\,
            WE => \N__28364\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51192\,
            RE => \N__28807\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN_net\,
            WE => \N__28359\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51317\,
            RE => \N__28849\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN_net\,
            WE => \N__28354\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51158\,
            RE => \N__28806\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN_net\,
            WE => \N__28358\
        );

    \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RDATA_wire\,
            RADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_RADDR_wire\,
            WADDR => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_WADDR_wire\,
            MASK => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_MASK_wire\,
            WDATA => \raw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__51319\,
            RE => \N__28853\,
            WCLKE => 'H',
            WCLK => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN_net\,
            WE => \N__28363\
        );

    \ipInertedIOPad_M_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54255\,
            DIN => \N__54254\,
            DOUT => \N__54253\,
            PACKAGEPIN => \M_CS1_wire\
        );

    \ipInertedIOPad_M_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54255\,
            PADOUT => \N__54254\,
            PADIN => \N__54253\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18920\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SYSCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54246\,
            DIN => \N__54245\,
            DOUT => \N__54244\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ipInertedIOPad_ICE_SYSCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54246\,
            PADOUT => \N__54245\,
            PADIN => \N__54244\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SYSCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54237\,
            DIN => \N__54236\,
            DOUT => \N__54235\,
            PACKAGEPIN => \M_MOSI1_wire\
        );

    \ipInertedIOPad_M_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54237\,
            PADOUT => \N__54236\,
            PADIN => \N__54235\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_DRDY1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54228\,
            DIN => \N__54227\,
            DOUT => \N__54226\,
            PACKAGEPIN => \M_DRDY1_wire\
        );

    \ipInertedIOPad_M_DRDY1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54228\,
            PADOUT => \N__54227\,
            PADIN => \N__54226\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_DRDY1\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CLK2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54219\,
            DIN => \N__54218\,
            DOUT => \N__54217\,
            PACKAGEPIN => \M_CLK2_wire\
        );

    \ipInertedIOPad_M_CLK2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54219\,
            PADOUT => \N__54218\,
            PADIN => \N__54217\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16753\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_SCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54210\,
            DIN => \N__54209\,
            DOUT => \N__54208\,
            PACKAGEPIN => \M_SCLK1_wire\
        );

    \ipInertedIOPad_M_SCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54210\,
            PADOUT => \N__54209\,
            PADIN => \N__54208\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18890\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54201\,
            DIN => \N__54200\,
            DOUT => \N__54199\,
            PACKAGEPIN => \M_FLT0_wire\
        );

    \ipInertedIOPad_M_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54201\,
            PADOUT => \N__54200\,
            PADIN => \N__54199\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28568\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CS3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54192\,
            DIN => \N__54191\,
            DOUT => \N__54190\,
            PACKAGEPIN => \M_CS3_wire\
        );

    \ipInertedIOPad_M_CS3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54192\,
            PADOUT => \N__54191\,
            PADIN => \N__54190\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20708\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_CHKCABLE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54183\,
            DIN => \N__54182\,
            DOUT => \N__54181\,
            PACKAGEPIN => \ICE_CHKCABLE_wire\
        );

    \ipInertedIOPad_ICE_CHKCABLE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54183\,
            PADOUT => \N__54182\,
            PADIN => \N__54181\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_CHKCABLE\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54174\,
            DIN => \N__54173\,
            DOUT => \N__54172\,
            PACKAGEPIN => \M_OSR1_wire\
        );

    \ipInertedIOPad_M_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54174\,
            PADOUT => \N__54173\,
            PADIN => \N__54172\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29441\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__54165\,
            DIN => \N__54164\,
            DOUT => \N__54163\,
            PACKAGEPIN => \ICE_GPMO_1_wire\
        );

    \ipInertedIOPad_ICE_GPMO_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54165\,
            PADOUT => \N__54164\,
            PADIN => \N__54163\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_EIS_SYNCCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__54156\,
            DIN => \N__54155\,
            DOUT => \N__54154\,
            PACKAGEPIN => \EIS_SYNCCLK_wire\
        );

    \ipInertedIOPad_EIS_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54156\,
            PADOUT => \N__54155\,
            PADIN => \N__54154\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_CLK4\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_SCLK3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54147\,
            DIN => \N__54146\,
            DOUT => \N__54145\,
            PACKAGEPIN => \M_SCLK3_wire\
        );

    \ipInertedIOPad_M_SCLK3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54147\,
            PADOUT => \N__54146\,
            PADIN => \N__54145\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20678\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54138\,
            DIN => \N__54137\,
            DOUT => \N__54136\,
            PACKAGEPIN => \M_OSR0_wire\
        );

    \ipInertedIOPad_M_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54138\,
            PADOUT => \N__54137\,
            PADIN => \N__54136\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28085\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MISO4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54129\,
            DIN => \N__54128\,
            DOUT => \N__54127\,
            PACKAGEPIN => \M_MISO4_wire\
        );

    \ipInertedIOPad_M_MISO4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54129\,
            PADOUT => \N__54128\,
            PADIN => \N__54127\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_MISO4\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_DRDY4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54120\,
            DIN => \N__54119\,
            DOUT => \N__54118\,
            PACKAGEPIN => \M_DRDY4_wire\
        );

    \ipInertedIOPad_M_DRDY4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54120\,
            PADOUT => \N__54119\,
            PADIN => \N__54118\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_DRDY4\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MOSI_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__54111\,
            DIN => \N__54110\,
            DOUT => \N__54109\,
            PACKAGEPIN => \ICE_SPI_MOSI_wire\
        );

    \ipInertedIOPad_ICE_SPI_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54111\,
            PADOUT => \N__54110\,
            PADIN => \N__54109\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_MOSI\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__54102\,
            DIN => \N__54101\,
            DOUT => \N__54100\,
            PACKAGEPIN => \ICE_GPMO_0_wire\
        );

    \ipInertedIOPad_ICE_GPMO_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54102\,
            PADOUT => \N__54101\,
            PADIN => \N__54100\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54093\,
            DIN => \N__54092\,
            DOUT => \N__54091\,
            PACKAGEPIN => \DDS_MOSI1_wire\
        );

    \ipInertedIOPad_DDS_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54093\,
            PADOUT => \N__54092\,
            PADIN => \N__54091\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21224\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_SCLK4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54084\,
            DIN => \N__54083\,
            DOUT => \N__54082\,
            PACKAGEPIN => \M_SCLK4_wire\
        );

    \ipInertedIOPad_M_SCLK4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54084\,
            PADOUT => \N__54083\,
            PADIN => \N__54082\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21650\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MISO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54075\,
            DIN => \N__54074\,
            DOUT => \N__54073\,
            PACKAGEPIN => \M_MISO3_wire\
        );

    \ipInertedIOPad_M_MISO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54075\,
            PADOUT => \N__54074\,
            PADIN => \N__54073\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_MISO3\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CS4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54066\,
            DIN => \N__54065\,
            DOUT => \N__54064\,
            PACKAGEPIN => \M_CS4_wire\
        );

    \ipInertedIOPad_M_CS4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54066\,
            PADOUT => \N__54065\,
            PADIN => \N__54064\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26594\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_SCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__54057\,
            DIN => \N__54056\,
            DOUT => \N__54055\,
            PACKAGEPIN => \ICE_SPI_SCLK_wire\
        );

    \ipInertedIOPad_ICE_SPI_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54057\,
            PADOUT => \N__54056\,
            PADIN => \N__54055\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_SCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MOSI4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54048\,
            DIN => \N__54047\,
            DOUT => \N__54046\,
            PACKAGEPIN => \M_MOSI4_wire\
        );

    \ipInertedIOPad_M_MOSI4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54048\,
            PADOUT => \N__54047\,
            PADIN => \N__54046\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MISO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54039\,
            DIN => \N__54038\,
            DOUT => \N__54037\,
            PACKAGEPIN => \M_MISO2_wire\
        );

    \ipInertedIOPad_M_MISO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54039\,
            PADOUT => \N__54038\,
            PADIN => \N__54037\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_MISO2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_DRDY2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54030\,
            DIN => \N__54029\,
            DOUT => \N__54028\,
            PACKAGEPIN => \M_DRDY2_wire\
        );

    \ipInertedIOPad_M_DRDY2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54030\,
            PADOUT => \N__54029\,
            PADIN => \N__54028\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_DRDY2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54021\,
            DIN => \N__54020\,
            DOUT => \N__54019\,
            PACKAGEPIN => \M_CLK1_wire\
        );

    \ipInertedIOPad_M_CLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54021\,
            PADOUT => \N__54020\,
            PADIN => \N__54019\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16745\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__54012\,
            DIN => \N__54011\,
            DOUT => \N__54010\,
            PACKAGEPIN => \ICE_SPI_MISO_wire\
        );

    \ipInertedIOPad_ICE_SPI_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54012\,
            PADOUT => \N__54011\,
            PADIN => \N__54010\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30290\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__54003\,
            DIN => \N__54002\,
            DOUT => \N__54001\,
            PACKAGEPIN => \ICE_GPMO_2_wire\
        );

    \ipInertedIOPad_ICE_GPMO_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__54003\,
            PADOUT => \N__54002\,
            PADIN => \N__54001\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMI_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53994\,
            DIN => \N__53993\,
            DOUT => \N__53992\,
            PACKAGEPIN => \ICE_GPMI_0_wire\
        );

    \ipInertedIOPad_ICE_GPMI_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53994\,
            PADOUT => \N__53993\,
            PADIN => \N__53992\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__46313\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TEST_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53985\,
            DIN => \N__53984\,
            DOUT => \N__53983\,
            PACKAGEPIN => \TEST_LED_wire\
        );

    \ipInertedIOPad_TEST_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53985\,
            PADOUT => \N__53984\,
            PADIN => \N__53983\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16796\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_POW_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53976\,
            DIN => \N__53975\,
            DOUT => \N__53974\,
            PACKAGEPIN => \M_POW_wire\
        );

    \ipInertedIOPad_M_POW_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53976\,
            PADOUT => \N__53975\,
            PADIN => \N__53974\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26267\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MOSI3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53967\,
            DIN => \N__53966\,
            DOUT => \N__53965\,
            PACKAGEPIN => \M_MOSI3_wire\
        );

    \ipInertedIOPad_M_MOSI3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53967\,
            PADOUT => \N__53966\,
            PADIN => \N__53965\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MISO1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53958\,
            DIN => \N__53957\,
            DOUT => \N__53956\,
            PACKAGEPIN => \M_MISO1_wire\
        );

    \ipInertedIOPad_M_MISO1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53958\,
            PADOUT => \N__53957\,
            PADIN => \N__53956\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_MISO1\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_DRDY3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53949\,
            DIN => \N__53948\,
            DOUT => \N__53947\,
            PACKAGEPIN => \M_DRDY3_wire\
        );

    \ipInertedIOPad_M_DRDY3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53949\,
            PADOUT => \N__53948\,
            PADIN => \N__53947\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \M_DRDY3\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_DCSEL_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53940\,
            DIN => \N__53939\,
            DOUT => \N__53938\,
            PACKAGEPIN => \M_DCSEL_wire\
        );

    \ipInertedIOPad_M_DCSEL_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53940\,
            PADOUT => \N__53939\,
            PADIN => \N__53938\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27932\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_START_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53931\,
            DIN => \N__53930\,
            DOUT => \N__53929\,
            PACKAGEPIN => \M_START_wire\
        );

    \ipInertedIOPad_M_START_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53931\,
            PADOUT => \N__53930\,
            PADIN => \N__53929\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19766\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_MOSI2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53922\,
            DIN => \N__53921\,
            DOUT => \N__53920\,
            PACKAGEPIN => \M_MOSI2_wire\
        );

    \ipInertedIOPad_M_MOSI2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53922\,
            PADOUT => \N__53921\,
            PADIN => \N__53920\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CLK3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53913\,
            DIN => \N__53912\,
            DOUT => \N__53911\,
            PACKAGEPIN => \M_CLK3_wire\
        );

    \ipInertedIOPad_M_CLK3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53913\,
            PADOUT => \N__53912\,
            PADIN => \N__53911\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16749\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53904\,
            DIN => \N__53903\,
            DOUT => \N__53902\,
            PACKAGEPIN => \DDS_CS1_wire\
        );

    \ipInertedIOPad_DDS_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53904\,
            PADOUT => \N__53903\,
            PADIN => \N__53902\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26900\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53895\,
            DIN => \N__53894\,
            DOUT => \N__53893\,
            PACKAGEPIN => \M_FLT1_wire\
        );

    \ipInertedIOPad_M_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53895\,
            PADOUT => \N__53894\,
            PADIN => \N__53893\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29585\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DISP_COMM_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53886\,
            DIN => \N__53885\,
            DOUT => \N__53884\,
            PACKAGEPIN => \DISP_COMM_wire\
        );

    \ipInertedIOPad_DISP_COMM_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53886\,
            PADOUT => \N__53885\,
            PADIN => \N__53884\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16673\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53877\,
            DIN => \N__53876\,
            DOUT => \N__53875\,
            PACKAGEPIN => \DDS_MCLK1_wire\
        );

    \ipInertedIOPad_DDS_MCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53877\,
            PADOUT => \N__53876\,
            PADIN => \N__53875\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16889\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_CE0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__53868\,
            DIN => \N__53867\,
            DOUT => \N__53866\,
            PACKAGEPIN => \ICE_SPI_CE0_wire\
        );

    \ipInertedIOPad_ICE_SPI_CE0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53868\,
            PADOUT => \N__53867\,
            PADIN => \N__53866\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_CE0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_SCLK2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53859\,
            DIN => \N__53858\,
            DOUT => \N__53857\,
            PACKAGEPIN => \M_SCLK2_wire\
        );

    \ipInertedIOPad_M_SCLK2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53859\,
            PADOUT => \N__53858\,
            PADIN => \N__53857\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19361\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CS2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53850\,
            DIN => \N__53849\,
            DOUT => \N__53848\,
            PACKAGEPIN => \M_CS2_wire\
        );

    \ipInertedIOPad_M_CS2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53850\,
            PADOUT => \N__53849\,
            PADIN => \N__53848\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17387\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_M_CLK4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53841\,
            DIN => \N__53840\,
            DOUT => \N__53839\,
            PACKAGEPIN => \M_CLK4_wire\
        );

    \ipInertedIOPad_M_CLK4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53841\,
            PADOUT => \N__53840\,
            PADIN => \N__53839\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16754\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__53832\,
            DIN => \N__53831\,
            DOUT => \N__53830\,
            PACKAGEPIN => \DDS_SCK1_wire\
        );

    \ipInertedIOPad_DDS_SCK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__53832\,
            PADOUT => \N__53831\,
            PADIN => \N__53830\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21059\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__13727\ : InMux
    port map (
            O => \N__53813\,
            I => \N__53806\
        );

    \I__13726\ : InMux
    port map (
            O => \N__53812\,
            I => \N__53803\
        );

    \I__13725\ : InMux
    port map (
            O => \N__53811\,
            I => \N__53800\
        );

    \I__13724\ : InMux
    port map (
            O => \N__53810\,
            I => \N__53795\
        );

    \I__13723\ : InMux
    port map (
            O => \N__53809\,
            I => \N__53792\
        );

    \I__13722\ : LocalMux
    port map (
            O => \N__53806\,
            I => \N__53785\
        );

    \I__13721\ : LocalMux
    port map (
            O => \N__53803\,
            I => \N__53785\
        );

    \I__13720\ : LocalMux
    port map (
            O => \N__53800\,
            I => \N__53785\
        );

    \I__13719\ : InMux
    port map (
            O => \N__53799\,
            I => \N__53782\
        );

    \I__13718\ : InMux
    port map (
            O => \N__53798\,
            I => \N__53779\
        );

    \I__13717\ : LocalMux
    port map (
            O => \N__53795\,
            I => \N__53776\
        );

    \I__13716\ : LocalMux
    port map (
            O => \N__53792\,
            I => \N__53771\
        );

    \I__13715\ : Span4Mux_v
    port map (
            O => \N__53785\,
            I => \N__53766\
        );

    \I__13714\ : LocalMux
    port map (
            O => \N__53782\,
            I => \N__53766\
        );

    \I__13713\ : LocalMux
    port map (
            O => \N__53779\,
            I => \N__53761\
        );

    \I__13712\ : Span4Mux_h
    port map (
            O => \N__53776\,
            I => \N__53761\
        );

    \I__13711\ : InMux
    port map (
            O => \N__53775\,
            I => \N__53758\
        );

    \I__13710\ : InMux
    port map (
            O => \N__53774\,
            I => \N__53755\
        );

    \I__13709\ : Span4Mux_h
    port map (
            O => \N__53771\,
            I => \N__53740\
        );

    \I__13708\ : Span4Mux_v
    port map (
            O => \N__53766\,
            I => \N__53740\
        );

    \I__13707\ : Span4Mux_v
    port map (
            O => \N__53761\,
            I => \N__53740\
        );

    \I__13706\ : LocalMux
    port map (
            O => \N__53758\,
            I => \N__53740\
        );

    \I__13705\ : LocalMux
    port map (
            O => \N__53755\,
            I => \N__53740\
        );

    \I__13704\ : InMux
    port map (
            O => \N__53754\,
            I => \N__53735\
        );

    \I__13703\ : InMux
    port map (
            O => \N__53753\,
            I => \N__53735\
        );

    \I__13702\ : InMux
    port map (
            O => \N__53752\,
            I => \N__53730\
        );

    \I__13701\ : InMux
    port map (
            O => \N__53751\,
            I => \N__53727\
        );

    \I__13700\ : Span4Mux_v
    port map (
            O => \N__53740\,
            I => \N__53722\
        );

    \I__13699\ : LocalMux
    port map (
            O => \N__53735\,
            I => \N__53722\
        );

    \I__13698\ : InMux
    port map (
            O => \N__53734\,
            I => \N__53717\
        );

    \I__13697\ : InMux
    port map (
            O => \N__53733\,
            I => \N__53717\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__53730\,
            I => \N__53713\
        );

    \I__13695\ : LocalMux
    port map (
            O => \N__53727\,
            I => \N__53710\
        );

    \I__13694\ : Span4Mux_v
    port map (
            O => \N__53722\,
            I => \N__53705\
        );

    \I__13693\ : LocalMux
    port map (
            O => \N__53717\,
            I => \N__53705\
        );

    \I__13692\ : InMux
    port map (
            O => \N__53716\,
            I => \N__53699\
        );

    \I__13691\ : Span4Mux_h
    port map (
            O => \N__53713\,
            I => \N__53692\
        );

    \I__13690\ : Span4Mux_h
    port map (
            O => \N__53710\,
            I => \N__53689\
        );

    \I__13689\ : Span4Mux_v
    port map (
            O => \N__53705\,
            I => \N__53686\
        );

    \I__13688\ : InMux
    port map (
            O => \N__53704\,
            I => \N__53678\
        );

    \I__13687\ : InMux
    port map (
            O => \N__53703\,
            I => \N__53678\
        );

    \I__13686\ : InMux
    port map (
            O => \N__53702\,
            I => \N__53678\
        );

    \I__13685\ : LocalMux
    port map (
            O => \N__53699\,
            I => \N__53675\
        );

    \I__13684\ : InMux
    port map (
            O => \N__53698\,
            I => \N__53672\
        );

    \I__13683\ : InMux
    port map (
            O => \N__53697\,
            I => \N__53669\
        );

    \I__13682\ : InMux
    port map (
            O => \N__53696\,
            I => \N__53664\
        );

    \I__13681\ : InMux
    port map (
            O => \N__53695\,
            I => \N__53664\
        );

    \I__13680\ : Span4Mux_h
    port map (
            O => \N__53692\,
            I => \N__53661\
        );

    \I__13679\ : Span4Mux_v
    port map (
            O => \N__53689\,
            I => \N__53656\
        );

    \I__13678\ : Span4Mux_h
    port map (
            O => \N__53686\,
            I => \N__53656\
        );

    \I__13677\ : InMux
    port map (
            O => \N__53685\,
            I => \N__53653\
        );

    \I__13676\ : LocalMux
    port map (
            O => \N__53678\,
            I => \N__53650\
        );

    \I__13675\ : Span4Mux_h
    port map (
            O => \N__53675\,
            I => \N__53647\
        );

    \I__13674\ : LocalMux
    port map (
            O => \N__53672\,
            I => \N__53642\
        );

    \I__13673\ : LocalMux
    port map (
            O => \N__53669\,
            I => \N__53642\
        );

    \I__13672\ : LocalMux
    port map (
            O => \N__53664\,
            I => \N__53639\
        );

    \I__13671\ : Span4Mux_h
    port map (
            O => \N__53661\,
            I => \N__53636\
        );

    \I__13670\ : Sp12to4
    port map (
            O => \N__53656\,
            I => \N__53633\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__53653\,
            I => \N__53626\
        );

    \I__13668\ : Span4Mux_h
    port map (
            O => \N__53650\,
            I => \N__53626\
        );

    \I__13667\ : Span4Mux_h
    port map (
            O => \N__53647\,
            I => \N__53626\
        );

    \I__13666\ : Span4Mux_h
    port map (
            O => \N__53642\,
            I => \N__53619\
        );

    \I__13665\ : Span4Mux_v
    port map (
            O => \N__53639\,
            I => \N__53619\
        );

    \I__13664\ : Span4Mux_v
    port map (
            O => \N__53636\,
            I => \N__53619\
        );

    \I__13663\ : Span12Mux_h
    port map (
            O => \N__53633\,
            I => \N__53616\
        );

    \I__13662\ : Odrv4
    port map (
            O => \N__53626\,
            I => n15150
        );

    \I__13661\ : Odrv4
    port map (
            O => \N__53619\,
            I => n15150
        );

    \I__13660\ : Odrv12
    port map (
            O => \N__53616\,
            I => n15150
        );

    \I__13659\ : CascadeMux
    port map (
            O => \N__53609\,
            I => \N__53606\
        );

    \I__13658\ : InMux
    port map (
            O => \N__53606\,
            I => \N__53602\
        );

    \I__13657\ : InMux
    port map (
            O => \N__53605\,
            I => \N__53599\
        );

    \I__13656\ : LocalMux
    port map (
            O => \N__53602\,
            I => \N__53596\
        );

    \I__13655\ : LocalMux
    port map (
            O => \N__53599\,
            I => \N__53593\
        );

    \I__13654\ : Span4Mux_h
    port map (
            O => \N__53596\,
            I => \N__53589\
        );

    \I__13653\ : Span4Mux_h
    port map (
            O => \N__53593\,
            I => \N__53586\
        );

    \I__13652\ : InMux
    port map (
            O => \N__53592\,
            I => \N__53583\
        );

    \I__13651\ : Odrv4
    port map (
            O => \N__53589\,
            I => cmd_rdadctmp_22_adj_1054
        );

    \I__13650\ : Odrv4
    port map (
            O => \N__53586\,
            I => cmd_rdadctmp_22_adj_1054
        );

    \I__13649\ : LocalMux
    port map (
            O => \N__53583\,
            I => cmd_rdadctmp_22_adj_1054
        );

    \I__13648\ : CascadeMux
    port map (
            O => \N__53576\,
            I => \N__53566\
        );

    \I__13647\ : InMux
    port map (
            O => \N__53575\,
            I => \N__53561\
        );

    \I__13646\ : InMux
    port map (
            O => \N__53574\,
            I => \N__53561\
        );

    \I__13645\ : InMux
    port map (
            O => \N__53573\,
            I => \N__53552\
        );

    \I__13644\ : InMux
    port map (
            O => \N__53572\,
            I => \N__53552\
        );

    \I__13643\ : InMux
    port map (
            O => \N__53571\,
            I => \N__53552\
        );

    \I__13642\ : InMux
    port map (
            O => \N__53570\,
            I => \N__53552\
        );

    \I__13641\ : InMux
    port map (
            O => \N__53569\,
            I => \N__53549\
        );

    \I__13640\ : InMux
    port map (
            O => \N__53566\,
            I => \N__53546\
        );

    \I__13639\ : LocalMux
    port map (
            O => \N__53561\,
            I => \N__53543\
        );

    \I__13638\ : LocalMux
    port map (
            O => \N__53552\,
            I => \N__53540\
        );

    \I__13637\ : LocalMux
    port map (
            O => \N__53549\,
            I => \N__53528\
        );

    \I__13636\ : LocalMux
    port map (
            O => \N__53546\,
            I => \N__53510\
        );

    \I__13635\ : Span4Mux_v
    port map (
            O => \N__53543\,
            I => \N__53510\
        );

    \I__13634\ : Span4Mux_h
    port map (
            O => \N__53540\,
            I => \N__53507\
        );

    \I__13633\ : InMux
    port map (
            O => \N__53539\,
            I => \N__53494\
        );

    \I__13632\ : InMux
    port map (
            O => \N__53538\,
            I => \N__53494\
        );

    \I__13631\ : InMux
    port map (
            O => \N__53537\,
            I => \N__53494\
        );

    \I__13630\ : InMux
    port map (
            O => \N__53536\,
            I => \N__53494\
        );

    \I__13629\ : InMux
    port map (
            O => \N__53535\,
            I => \N__53494\
        );

    \I__13628\ : InMux
    port map (
            O => \N__53534\,
            I => \N__53494\
        );

    \I__13627\ : InMux
    port map (
            O => \N__53533\,
            I => \N__53489\
        );

    \I__13626\ : InMux
    port map (
            O => \N__53532\,
            I => \N__53484\
        );

    \I__13625\ : InMux
    port map (
            O => \N__53531\,
            I => \N__53484\
        );

    \I__13624\ : Span4Mux_h
    port map (
            O => \N__53528\,
            I => \N__53478\
        );

    \I__13623\ : InMux
    port map (
            O => \N__53527\,
            I => \N__53475\
        );

    \I__13622\ : InMux
    port map (
            O => \N__53526\,
            I => \N__53471\
        );

    \I__13621\ : InMux
    port map (
            O => \N__53525\,
            I => \N__53468\
        );

    \I__13620\ : InMux
    port map (
            O => \N__53524\,
            I => \N__53457\
        );

    \I__13619\ : InMux
    port map (
            O => \N__53523\,
            I => \N__53457\
        );

    \I__13618\ : InMux
    port map (
            O => \N__53522\,
            I => \N__53457\
        );

    \I__13617\ : InMux
    port map (
            O => \N__53521\,
            I => \N__53457\
        );

    \I__13616\ : InMux
    port map (
            O => \N__53520\,
            I => \N__53457\
        );

    \I__13615\ : InMux
    port map (
            O => \N__53519\,
            I => \N__53446\
        );

    \I__13614\ : InMux
    port map (
            O => \N__53518\,
            I => \N__53446\
        );

    \I__13613\ : InMux
    port map (
            O => \N__53517\,
            I => \N__53446\
        );

    \I__13612\ : InMux
    port map (
            O => \N__53516\,
            I => \N__53446\
        );

    \I__13611\ : InMux
    port map (
            O => \N__53515\,
            I => \N__53446\
        );

    \I__13610\ : Span4Mux_v
    port map (
            O => \N__53510\,
            I => \N__53439\
        );

    \I__13609\ : Span4Mux_v
    port map (
            O => \N__53507\,
            I => \N__53439\
        );

    \I__13608\ : LocalMux
    port map (
            O => \N__53494\,
            I => \N__53439\
        );

    \I__13607\ : InMux
    port map (
            O => \N__53493\,
            I => \N__53430\
        );

    \I__13606\ : InMux
    port map (
            O => \N__53492\,
            I => \N__53427\
        );

    \I__13605\ : LocalMux
    port map (
            O => \N__53489\,
            I => \N__53422\
        );

    \I__13604\ : LocalMux
    port map (
            O => \N__53484\,
            I => \N__53422\
        );

    \I__13603\ : InMux
    port map (
            O => \N__53483\,
            I => \N__53417\
        );

    \I__13602\ : InMux
    port map (
            O => \N__53482\,
            I => \N__53417\
        );

    \I__13601\ : InMux
    port map (
            O => \N__53481\,
            I => \N__53414\
        );

    \I__13600\ : Span4Mux_v
    port map (
            O => \N__53478\,
            I => \N__53409\
        );

    \I__13599\ : LocalMux
    port map (
            O => \N__53475\,
            I => \N__53409\
        );

    \I__13598\ : InMux
    port map (
            O => \N__53474\,
            I => \N__53399\
        );

    \I__13597\ : LocalMux
    port map (
            O => \N__53471\,
            I => \N__53394\
        );

    \I__13596\ : LocalMux
    port map (
            O => \N__53468\,
            I => \N__53394\
        );

    \I__13595\ : LocalMux
    port map (
            O => \N__53457\,
            I => \N__53385\
        );

    \I__13594\ : LocalMux
    port map (
            O => \N__53446\,
            I => \N__53385\
        );

    \I__13593\ : Span4Mux_h
    port map (
            O => \N__53439\,
            I => \N__53382\
        );

    \I__13592\ : InMux
    port map (
            O => \N__53438\,
            I => \N__53379\
        );

    \I__13591\ : InMux
    port map (
            O => \N__53437\,
            I => \N__53370\
        );

    \I__13590\ : InMux
    port map (
            O => \N__53436\,
            I => \N__53370\
        );

    \I__13589\ : InMux
    port map (
            O => \N__53435\,
            I => \N__53370\
        );

    \I__13588\ : InMux
    port map (
            O => \N__53434\,
            I => \N__53370\
        );

    \I__13587\ : InMux
    port map (
            O => \N__53433\,
            I => \N__53367\
        );

    \I__13586\ : LocalMux
    port map (
            O => \N__53430\,
            I => \N__53362\
        );

    \I__13585\ : LocalMux
    port map (
            O => \N__53427\,
            I => \N__53362\
        );

    \I__13584\ : Span4Mux_h
    port map (
            O => \N__53422\,
            I => \N__53357\
        );

    \I__13583\ : LocalMux
    port map (
            O => \N__53417\,
            I => \N__53357\
        );

    \I__13582\ : LocalMux
    port map (
            O => \N__53414\,
            I => \N__53349\
        );

    \I__13581\ : Span4Mux_h
    port map (
            O => \N__53409\,
            I => \N__53349\
        );

    \I__13580\ : InMux
    port map (
            O => \N__53408\,
            I => \N__53336\
        );

    \I__13579\ : InMux
    port map (
            O => \N__53407\,
            I => \N__53336\
        );

    \I__13578\ : InMux
    port map (
            O => \N__53406\,
            I => \N__53336\
        );

    \I__13577\ : InMux
    port map (
            O => \N__53405\,
            I => \N__53336\
        );

    \I__13576\ : InMux
    port map (
            O => \N__53404\,
            I => \N__53336\
        );

    \I__13575\ : InMux
    port map (
            O => \N__53403\,
            I => \N__53336\
        );

    \I__13574\ : InMux
    port map (
            O => \N__53402\,
            I => \N__53332\
        );

    \I__13573\ : LocalMux
    port map (
            O => \N__53399\,
            I => \N__53329\
        );

    \I__13572\ : Span4Mux_h
    port map (
            O => \N__53394\,
            I => \N__53326\
        );

    \I__13571\ : InMux
    port map (
            O => \N__53393\,
            I => \N__53316\
        );

    \I__13570\ : InMux
    port map (
            O => \N__53392\,
            I => \N__53316\
        );

    \I__13569\ : InMux
    port map (
            O => \N__53391\,
            I => \N__53316\
        );

    \I__13568\ : InMux
    port map (
            O => \N__53390\,
            I => \N__53316\
        );

    \I__13567\ : Span4Mux_v
    port map (
            O => \N__53385\,
            I => \N__53313\
        );

    \I__13566\ : Span4Mux_h
    port map (
            O => \N__53382\,
            I => \N__53310\
        );

    \I__13565\ : LocalMux
    port map (
            O => \N__53379\,
            I => \N__53307\
        );

    \I__13564\ : LocalMux
    port map (
            O => \N__53370\,
            I => \N__53304\
        );

    \I__13563\ : LocalMux
    port map (
            O => \N__53367\,
            I => \N__53301\
        );

    \I__13562\ : Span4Mux_v
    port map (
            O => \N__53362\,
            I => \N__53298\
        );

    \I__13561\ : Span4Mux_h
    port map (
            O => \N__53357\,
            I => \N__53295\
        );

    \I__13560\ : InMux
    port map (
            O => \N__53356\,
            I => \N__53290\
        );

    \I__13559\ : InMux
    port map (
            O => \N__53355\,
            I => \N__53285\
        );

    \I__13558\ : InMux
    port map (
            O => \N__53354\,
            I => \N__53285\
        );

    \I__13557\ : Span4Mux_h
    port map (
            O => \N__53349\,
            I => \N__53282\
        );

    \I__13556\ : LocalMux
    port map (
            O => \N__53336\,
            I => \N__53279\
        );

    \I__13555\ : InMux
    port map (
            O => \N__53335\,
            I => \N__53272\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__53332\,
            I => \N__53269\
        );

    \I__13553\ : Span4Mux_v
    port map (
            O => \N__53329\,
            I => \N__53264\
        );

    \I__13552\ : Span4Mux_h
    port map (
            O => \N__53326\,
            I => \N__53264\
        );

    \I__13551\ : InMux
    port map (
            O => \N__53325\,
            I => \N__53261\
        );

    \I__13550\ : LocalMux
    port map (
            O => \N__53316\,
            I => \N__53258\
        );

    \I__13549\ : Span4Mux_h
    port map (
            O => \N__53313\,
            I => \N__53253\
        );

    \I__13548\ : Span4Mux_h
    port map (
            O => \N__53310\,
            I => \N__53253\
        );

    \I__13547\ : Span4Mux_h
    port map (
            O => \N__53307\,
            I => \N__53248\
        );

    \I__13546\ : Span4Mux_h
    port map (
            O => \N__53304\,
            I => \N__53248\
        );

    \I__13545\ : Span4Mux_h
    port map (
            O => \N__53301\,
            I => \N__53243\
        );

    \I__13544\ : Span4Mux_h
    port map (
            O => \N__53298\,
            I => \N__53243\
        );

    \I__13543\ : Span4Mux_v
    port map (
            O => \N__53295\,
            I => \N__53240\
        );

    \I__13542\ : InMux
    port map (
            O => \N__53294\,
            I => \N__53237\
        );

    \I__13541\ : InMux
    port map (
            O => \N__53293\,
            I => \N__53234\
        );

    \I__13540\ : LocalMux
    port map (
            O => \N__53290\,
            I => \N__53229\
        );

    \I__13539\ : LocalMux
    port map (
            O => \N__53285\,
            I => \N__53229\
        );

    \I__13538\ : Span4Mux_h
    port map (
            O => \N__53282\,
            I => \N__53224\
        );

    \I__13537\ : Span4Mux_h
    port map (
            O => \N__53279\,
            I => \N__53224\
        );

    \I__13536\ : InMux
    port map (
            O => \N__53278\,
            I => \N__53216\
        );

    \I__13535\ : InMux
    port map (
            O => \N__53277\,
            I => \N__53213\
        );

    \I__13534\ : InMux
    port map (
            O => \N__53276\,
            I => \N__53210\
        );

    \I__13533\ : InMux
    port map (
            O => \N__53275\,
            I => \N__53207\
        );

    \I__13532\ : LocalMux
    port map (
            O => \N__53272\,
            I => \N__53204\
        );

    \I__13531\ : Span4Mux_h
    port map (
            O => \N__53269\,
            I => \N__53199\
        );

    \I__13530\ : Span4Mux_h
    port map (
            O => \N__53264\,
            I => \N__53199\
        );

    \I__13529\ : LocalMux
    port map (
            O => \N__53261\,
            I => \N__53192\
        );

    \I__13528\ : Span12Mux_h
    port map (
            O => \N__53258\,
            I => \N__53192\
        );

    \I__13527\ : Sp12to4
    port map (
            O => \N__53253\,
            I => \N__53192\
        );

    \I__13526\ : Span4Mux_h
    port map (
            O => \N__53248\,
            I => \N__53185\
        );

    \I__13525\ : Span4Mux_h
    port map (
            O => \N__53243\,
            I => \N__53185\
        );

    \I__13524\ : Span4Mux_h
    port map (
            O => \N__53240\,
            I => \N__53185\
        );

    \I__13523\ : LocalMux
    port map (
            O => \N__53237\,
            I => \N__53176\
        );

    \I__13522\ : LocalMux
    port map (
            O => \N__53234\,
            I => \N__53176\
        );

    \I__13521\ : Span4Mux_h
    port map (
            O => \N__53229\,
            I => \N__53176\
        );

    \I__13520\ : Span4Mux_h
    port map (
            O => \N__53224\,
            I => \N__53176\
        );

    \I__13519\ : InMux
    port map (
            O => \N__53223\,
            I => \N__53165\
        );

    \I__13518\ : InMux
    port map (
            O => \N__53222\,
            I => \N__53165\
        );

    \I__13517\ : InMux
    port map (
            O => \N__53221\,
            I => \N__53165\
        );

    \I__13516\ : InMux
    port map (
            O => \N__53220\,
            I => \N__53165\
        );

    \I__13515\ : InMux
    port map (
            O => \N__53219\,
            I => \N__53165\
        );

    \I__13514\ : LocalMux
    port map (
            O => \N__53216\,
            I => adc_state_0_adj_1044
        );

    \I__13513\ : LocalMux
    port map (
            O => \N__53213\,
            I => adc_state_0_adj_1044
        );

    \I__13512\ : LocalMux
    port map (
            O => \N__53210\,
            I => adc_state_0_adj_1044
        );

    \I__13511\ : LocalMux
    port map (
            O => \N__53207\,
            I => adc_state_0_adj_1044
        );

    \I__13510\ : Odrv12
    port map (
            O => \N__53204\,
            I => adc_state_0_adj_1044
        );

    \I__13509\ : Odrv4
    port map (
            O => \N__53199\,
            I => adc_state_0_adj_1044
        );

    \I__13508\ : Odrv12
    port map (
            O => \N__53192\,
            I => adc_state_0_adj_1044
        );

    \I__13507\ : Odrv4
    port map (
            O => \N__53185\,
            I => adc_state_0_adj_1044
        );

    \I__13506\ : Odrv4
    port map (
            O => \N__53176\,
            I => adc_state_0_adj_1044
        );

    \I__13505\ : LocalMux
    port map (
            O => \N__53165\,
            I => adc_state_0_adj_1044
        );

    \I__13504\ : InMux
    port map (
            O => \N__53144\,
            I => \N__53140\
        );

    \I__13503\ : InMux
    port map (
            O => \N__53143\,
            I => \N__53137\
        );

    \I__13502\ : LocalMux
    port map (
            O => \N__53140\,
            I => \N__53134\
        );

    \I__13501\ : LocalMux
    port map (
            O => \N__53137\,
            I => buf_adcdata2_14
        );

    \I__13500\ : Odrv4
    port map (
            O => \N__53134\,
            I => buf_adcdata2_14
        );

    \I__13499\ : InMux
    port map (
            O => \N__53129\,
            I => \N__53118\
        );

    \I__13498\ : InMux
    port map (
            O => \N__53128\,
            I => \N__53118\
        );

    \I__13497\ : InMux
    port map (
            O => \N__53127\,
            I => \N__53107\
        );

    \I__13496\ : InMux
    port map (
            O => \N__53126\,
            I => \N__53107\
        );

    \I__13495\ : InMux
    port map (
            O => \N__53125\,
            I => \N__53107\
        );

    \I__13494\ : InMux
    port map (
            O => \N__53124\,
            I => \N__53102\
        );

    \I__13493\ : InMux
    port map (
            O => \N__53123\,
            I => \N__53102\
        );

    \I__13492\ : LocalMux
    port map (
            O => \N__53118\,
            I => \N__53098\
        );

    \I__13491\ : InMux
    port map (
            O => \N__53117\,
            I => \N__53095\
        );

    \I__13490\ : InMux
    port map (
            O => \N__53116\,
            I => \N__53092\
        );

    \I__13489\ : InMux
    port map (
            O => \N__53115\,
            I => \N__53089\
        );

    \I__13488\ : InMux
    port map (
            O => \N__53114\,
            I => \N__53086\
        );

    \I__13487\ : LocalMux
    port map (
            O => \N__53107\,
            I => \N__53079\
        );

    \I__13486\ : LocalMux
    port map (
            O => \N__53102\,
            I => \N__53079\
        );

    \I__13485\ : InMux
    port map (
            O => \N__53101\,
            I => \N__53072\
        );

    \I__13484\ : Span4Mux_v
    port map (
            O => \N__53098\,
            I => \N__53065\
        );

    \I__13483\ : LocalMux
    port map (
            O => \N__53095\,
            I => \N__53065\
        );

    \I__13482\ : LocalMux
    port map (
            O => \N__53092\,
            I => \N__53065\
        );

    \I__13481\ : LocalMux
    port map (
            O => \N__53089\,
            I => \N__53060\
        );

    \I__13480\ : LocalMux
    port map (
            O => \N__53086\,
            I => \N__53057\
        );

    \I__13479\ : InMux
    port map (
            O => \N__53085\,
            I => \N__53052\
        );

    \I__13478\ : InMux
    port map (
            O => \N__53084\,
            I => \N__53052\
        );

    \I__13477\ : Span4Mux_v
    port map (
            O => \N__53079\,
            I => \N__53046\
        );

    \I__13476\ : InMux
    port map (
            O => \N__53078\,
            I => \N__53037\
        );

    \I__13475\ : InMux
    port map (
            O => \N__53077\,
            I => \N__53037\
        );

    \I__13474\ : InMux
    port map (
            O => \N__53076\,
            I => \N__53037\
        );

    \I__13473\ : InMux
    port map (
            O => \N__53075\,
            I => \N__53037\
        );

    \I__13472\ : LocalMux
    port map (
            O => \N__53072\,
            I => \N__53034\
        );

    \I__13471\ : Span4Mux_v
    port map (
            O => \N__53065\,
            I => \N__53031\
        );

    \I__13470\ : InMux
    port map (
            O => \N__53064\,
            I => \N__53028\
        );

    \I__13469\ : InMux
    port map (
            O => \N__53063\,
            I => \N__53025\
        );

    \I__13468\ : Span4Mux_v
    port map (
            O => \N__53060\,
            I => \N__53022\
        );

    \I__13467\ : Span4Mux_h
    port map (
            O => \N__53057\,
            I => \N__53019\
        );

    \I__13466\ : LocalMux
    port map (
            O => \N__53052\,
            I => \N__53016\
        );

    \I__13465\ : InMux
    port map (
            O => \N__53051\,
            I => \N__53012\
        );

    \I__13464\ : InMux
    port map (
            O => \N__53050\,
            I => \N__53009\
        );

    \I__13463\ : InMux
    port map (
            O => \N__53049\,
            I => \N__53006\
        );

    \I__13462\ : Span4Mux_h
    port map (
            O => \N__53046\,
            I => \N__53001\
        );

    \I__13461\ : LocalMux
    port map (
            O => \N__53037\,
            I => \N__53001\
        );

    \I__13460\ : Span4Mux_v
    port map (
            O => \N__53034\,
            I => \N__52998\
        );

    \I__13459\ : Span4Mux_h
    port map (
            O => \N__53031\,
            I => \N__52995\
        );

    \I__13458\ : LocalMux
    port map (
            O => \N__53028\,
            I => \N__52990\
        );

    \I__13457\ : LocalMux
    port map (
            O => \N__53025\,
            I => \N__52990\
        );

    \I__13456\ : Span4Mux_h
    port map (
            O => \N__53022\,
            I => \N__52987\
        );

    \I__13455\ : Span4Mux_h
    port map (
            O => \N__53019\,
            I => \N__52984\
        );

    \I__13454\ : Span4Mux_h
    port map (
            O => \N__53016\,
            I => \N__52981\
        );

    \I__13453\ : InMux
    port map (
            O => \N__53015\,
            I => \N__52978\
        );

    \I__13452\ : LocalMux
    port map (
            O => \N__53012\,
            I => \N__52969\
        );

    \I__13451\ : LocalMux
    port map (
            O => \N__53009\,
            I => \N__52969\
        );

    \I__13450\ : LocalMux
    port map (
            O => \N__53006\,
            I => \N__52969\
        );

    \I__13449\ : Span4Mux_h
    port map (
            O => \N__53001\,
            I => \N__52969\
        );

    \I__13448\ : Sp12to4
    port map (
            O => \N__52998\,
            I => \N__52966\
        );

    \I__13447\ : Sp12to4
    port map (
            O => \N__52995\,
            I => \N__52963\
        );

    \I__13446\ : Span4Mux_v
    port map (
            O => \N__52990\,
            I => \N__52956\
        );

    \I__13445\ : Span4Mux_h
    port map (
            O => \N__52987\,
            I => \N__52956\
        );

    \I__13444\ : Span4Mux_h
    port map (
            O => \N__52984\,
            I => \N__52956\
        );

    \I__13443\ : Span4Mux_h
    port map (
            O => \N__52981\,
            I => \N__52953\
        );

    \I__13442\ : LocalMux
    port map (
            O => \N__52978\,
            I => \N__52944\
        );

    \I__13441\ : Sp12to4
    port map (
            O => \N__52969\,
            I => \N__52944\
        );

    \I__13440\ : Span12Mux_h
    port map (
            O => \N__52966\,
            I => \N__52944\
        );

    \I__13439\ : Span12Mux_h
    port map (
            O => \N__52963\,
            I => \N__52944\
        );

    \I__13438\ : Span4Mux_h
    port map (
            O => \N__52956\,
            I => \N__52941\
        );

    \I__13437\ : Odrv4
    port map (
            O => \N__52953\,
            I => n15153
        );

    \I__13436\ : Odrv12
    port map (
            O => \N__52944\,
            I => n15153
        );

    \I__13435\ : Odrv4
    port map (
            O => \N__52941\,
            I => n15153
        );

    \I__13434\ : CascadeMux
    port map (
            O => \N__52934\,
            I => \N__52931\
        );

    \I__13433\ : InMux
    port map (
            O => \N__52931\,
            I => \N__52928\
        );

    \I__13432\ : LocalMux
    port map (
            O => \N__52928\,
            I => \N__52925\
        );

    \I__13431\ : Span4Mux_h
    port map (
            O => \N__52925\,
            I => \N__52922\
        );

    \I__13430\ : Span4Mux_h
    port map (
            O => \N__52922\,
            I => \N__52918\
        );

    \I__13429\ : CascadeMux
    port map (
            O => \N__52921\,
            I => \N__52914\
        );

    \I__13428\ : Span4Mux_h
    port map (
            O => \N__52918\,
            I => \N__52911\
        );

    \I__13427\ : InMux
    port map (
            O => \N__52917\,
            I => \N__52908\
        );

    \I__13426\ : InMux
    port map (
            O => \N__52914\,
            I => \N__52905\
        );

    \I__13425\ : Odrv4
    port map (
            O => \N__52911\,
            I => cmd_rdadctmp_18
        );

    \I__13424\ : LocalMux
    port map (
            O => \N__52908\,
            I => cmd_rdadctmp_18
        );

    \I__13423\ : LocalMux
    port map (
            O => \N__52905\,
            I => cmd_rdadctmp_18
        );

    \I__13422\ : CascadeMux
    port map (
            O => \N__52898\,
            I => \N__52885\
        );

    \I__13421\ : InMux
    port map (
            O => \N__52897\,
            I => \N__52871\
        );

    \I__13420\ : InMux
    port map (
            O => \N__52896\,
            I => \N__52868\
        );

    \I__13419\ : InMux
    port map (
            O => \N__52895\,
            I => \N__52863\
        );

    \I__13418\ : InMux
    port map (
            O => \N__52894\,
            I => \N__52863\
        );

    \I__13417\ : InMux
    port map (
            O => \N__52893\,
            I => \N__52860\
        );

    \I__13416\ : InMux
    port map (
            O => \N__52892\,
            I => \N__52857\
        );

    \I__13415\ : CascadeMux
    port map (
            O => \N__52891\,
            I => \N__52854\
        );

    \I__13414\ : CascadeMux
    port map (
            O => \N__52890\,
            I => \N__52841\
        );

    \I__13413\ : CascadeMux
    port map (
            O => \N__52889\,
            I => \N__52838\
        );

    \I__13412\ : InMux
    port map (
            O => \N__52888\,
            I => \N__52814\
        );

    \I__13411\ : InMux
    port map (
            O => \N__52885\,
            I => \N__52814\
        );

    \I__13410\ : InMux
    port map (
            O => \N__52884\,
            I => \N__52814\
        );

    \I__13409\ : InMux
    port map (
            O => \N__52883\,
            I => \N__52814\
        );

    \I__13408\ : InMux
    port map (
            O => \N__52882\,
            I => \N__52814\
        );

    \I__13407\ : InMux
    port map (
            O => \N__52881\,
            I => \N__52814\
        );

    \I__13406\ : InMux
    port map (
            O => \N__52880\,
            I => \N__52814\
        );

    \I__13405\ : InMux
    port map (
            O => \N__52879\,
            I => \N__52814\
        );

    \I__13404\ : CascadeMux
    port map (
            O => \N__52878\,
            I => \N__52810\
        );

    \I__13403\ : InMux
    port map (
            O => \N__52877\,
            I => \N__52806\
        );

    \I__13402\ : InMux
    port map (
            O => \N__52876\,
            I => \N__52799\
        );

    \I__13401\ : InMux
    port map (
            O => \N__52875\,
            I => \N__52799\
        );

    \I__13400\ : InMux
    port map (
            O => \N__52874\,
            I => \N__52799\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__52871\,
            I => \N__52790\
        );

    \I__13398\ : LocalMux
    port map (
            O => \N__52868\,
            I => \N__52785\
        );

    \I__13397\ : LocalMux
    port map (
            O => \N__52863\,
            I => \N__52785\
        );

    \I__13396\ : LocalMux
    port map (
            O => \N__52860\,
            I => \N__52782\
        );

    \I__13395\ : LocalMux
    port map (
            O => \N__52857\,
            I => \N__52779\
        );

    \I__13394\ : InMux
    port map (
            O => \N__52854\,
            I => \N__52775\
        );

    \I__13393\ : InMux
    port map (
            O => \N__52853\,
            I => \N__52763\
        );

    \I__13392\ : InMux
    port map (
            O => \N__52852\,
            I => \N__52763\
        );

    \I__13391\ : InMux
    port map (
            O => \N__52851\,
            I => \N__52763\
        );

    \I__13390\ : InMux
    port map (
            O => \N__52850\,
            I => \N__52763\
        );

    \I__13389\ : InMux
    port map (
            O => \N__52849\,
            I => \N__52763\
        );

    \I__13388\ : InMux
    port map (
            O => \N__52848\,
            I => \N__52760\
        );

    \I__13387\ : InMux
    port map (
            O => \N__52847\,
            I => \N__52757\
        );

    \I__13386\ : InMux
    port map (
            O => \N__52846\,
            I => \N__52754\
        );

    \I__13385\ : InMux
    port map (
            O => \N__52845\,
            I => \N__52751\
        );

    \I__13384\ : InMux
    port map (
            O => \N__52844\,
            I => \N__52748\
        );

    \I__13383\ : InMux
    port map (
            O => \N__52841\,
            I => \N__52745\
        );

    \I__13382\ : InMux
    port map (
            O => \N__52838\,
            I => \N__52742\
        );

    \I__13381\ : InMux
    port map (
            O => \N__52837\,
            I => \N__52739\
        );

    \I__13380\ : InMux
    port map (
            O => \N__52836\,
            I => \N__52736\
        );

    \I__13379\ : InMux
    port map (
            O => \N__52835\,
            I => \N__52725\
        );

    \I__13378\ : InMux
    port map (
            O => \N__52834\,
            I => \N__52725\
        );

    \I__13377\ : InMux
    port map (
            O => \N__52833\,
            I => \N__52725\
        );

    \I__13376\ : InMux
    port map (
            O => \N__52832\,
            I => \N__52725\
        );

    \I__13375\ : InMux
    port map (
            O => \N__52831\,
            I => \N__52725\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__52814\,
            I => \N__52722\
        );

    \I__13373\ : InMux
    port map (
            O => \N__52813\,
            I => \N__52719\
        );

    \I__13372\ : InMux
    port map (
            O => \N__52810\,
            I => \N__52714\
        );

    \I__13371\ : InMux
    port map (
            O => \N__52809\,
            I => \N__52714\
        );

    \I__13370\ : LocalMux
    port map (
            O => \N__52806\,
            I => \N__52711\
        );

    \I__13369\ : LocalMux
    port map (
            O => \N__52799\,
            I => \N__52708\
        );

    \I__13368\ : InMux
    port map (
            O => \N__52798\,
            I => \N__52699\
        );

    \I__13367\ : InMux
    port map (
            O => \N__52797\,
            I => \N__52699\
        );

    \I__13366\ : InMux
    port map (
            O => \N__52796\,
            I => \N__52699\
        );

    \I__13365\ : InMux
    port map (
            O => \N__52795\,
            I => \N__52699\
        );

    \I__13364\ : InMux
    port map (
            O => \N__52794\,
            I => \N__52696\
        );

    \I__13363\ : InMux
    port map (
            O => \N__52793\,
            I => \N__52693\
        );

    \I__13362\ : Span4Mux_v
    port map (
            O => \N__52790\,
            I => \N__52690\
        );

    \I__13361\ : Span4Mux_v
    port map (
            O => \N__52785\,
            I => \N__52683\
        );

    \I__13360\ : Span4Mux_v
    port map (
            O => \N__52782\,
            I => \N__52683\
        );

    \I__13359\ : Span4Mux_v
    port map (
            O => \N__52779\,
            I => \N__52683\
        );

    \I__13358\ : CascadeMux
    port map (
            O => \N__52778\,
            I => \N__52680\
        );

    \I__13357\ : LocalMux
    port map (
            O => \N__52775\,
            I => \N__52667\
        );

    \I__13356\ : InMux
    port map (
            O => \N__52774\,
            I => \N__52664\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__52763\,
            I => \N__52659\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__52760\,
            I => \N__52659\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__52757\,
            I => \N__52656\
        );

    \I__13352\ : LocalMux
    port map (
            O => \N__52754\,
            I => \N__52653\
        );

    \I__13351\ : LocalMux
    port map (
            O => \N__52751\,
            I => \N__52650\
        );

    \I__13350\ : LocalMux
    port map (
            O => \N__52748\,
            I => \N__52645\
        );

    \I__13349\ : LocalMux
    port map (
            O => \N__52745\,
            I => \N__52645\
        );

    \I__13348\ : LocalMux
    port map (
            O => \N__52742\,
            I => \N__52636\
        );

    \I__13347\ : LocalMux
    port map (
            O => \N__52739\,
            I => \N__52636\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__52736\,
            I => \N__52636\
        );

    \I__13345\ : LocalMux
    port map (
            O => \N__52725\,
            I => \N__52636\
        );

    \I__13344\ : Span4Mux_h
    port map (
            O => \N__52722\,
            I => \N__52631\
        );

    \I__13343\ : LocalMux
    port map (
            O => \N__52719\,
            I => \N__52631\
        );

    \I__13342\ : LocalMux
    port map (
            O => \N__52714\,
            I => \N__52628\
        );

    \I__13341\ : Span4Mux_v
    port map (
            O => \N__52711\,
            I => \N__52621\
        );

    \I__13340\ : Span4Mux_v
    port map (
            O => \N__52708\,
            I => \N__52621\
        );

    \I__13339\ : LocalMux
    port map (
            O => \N__52699\,
            I => \N__52621\
        );

    \I__13338\ : LocalMux
    port map (
            O => \N__52696\,
            I => \N__52607\
        );

    \I__13337\ : LocalMux
    port map (
            O => \N__52693\,
            I => \N__52607\
        );

    \I__13336\ : Sp12to4
    port map (
            O => \N__52690\,
            I => \N__52607\
        );

    \I__13335\ : Sp12to4
    port map (
            O => \N__52683\,
            I => \N__52607\
        );

    \I__13334\ : InMux
    port map (
            O => \N__52680\,
            I => \N__52598\
        );

    \I__13333\ : InMux
    port map (
            O => \N__52679\,
            I => \N__52598\
        );

    \I__13332\ : InMux
    port map (
            O => \N__52678\,
            I => \N__52595\
        );

    \I__13331\ : InMux
    port map (
            O => \N__52677\,
            I => \N__52578\
        );

    \I__13330\ : InMux
    port map (
            O => \N__52676\,
            I => \N__52578\
        );

    \I__13329\ : InMux
    port map (
            O => \N__52675\,
            I => \N__52578\
        );

    \I__13328\ : InMux
    port map (
            O => \N__52674\,
            I => \N__52578\
        );

    \I__13327\ : InMux
    port map (
            O => \N__52673\,
            I => \N__52578\
        );

    \I__13326\ : InMux
    port map (
            O => \N__52672\,
            I => \N__52578\
        );

    \I__13325\ : InMux
    port map (
            O => \N__52671\,
            I => \N__52578\
        );

    \I__13324\ : InMux
    port map (
            O => \N__52670\,
            I => \N__52578\
        );

    \I__13323\ : Span4Mux_h
    port map (
            O => \N__52667\,
            I => \N__52571\
        );

    \I__13322\ : LocalMux
    port map (
            O => \N__52664\,
            I => \N__52571\
        );

    \I__13321\ : Span4Mux_v
    port map (
            O => \N__52659\,
            I => \N__52571\
        );

    \I__13320\ : Span4Mux_v
    port map (
            O => \N__52656\,
            I => \N__52564\
        );

    \I__13319\ : Span4Mux_v
    port map (
            O => \N__52653\,
            I => \N__52564\
        );

    \I__13318\ : Span4Mux_v
    port map (
            O => \N__52650\,
            I => \N__52564\
        );

    \I__13317\ : Span4Mux_h
    port map (
            O => \N__52645\,
            I => \N__52559\
        );

    \I__13316\ : Span4Mux_h
    port map (
            O => \N__52636\,
            I => \N__52559\
        );

    \I__13315\ : Span4Mux_v
    port map (
            O => \N__52631\,
            I => \N__52552\
        );

    \I__13314\ : Span4Mux_v
    port map (
            O => \N__52628\,
            I => \N__52552\
        );

    \I__13313\ : Span4Mux_v
    port map (
            O => \N__52621\,
            I => \N__52552\
        );

    \I__13312\ : InMux
    port map (
            O => \N__52620\,
            I => \N__52545\
        );

    \I__13311\ : InMux
    port map (
            O => \N__52619\,
            I => \N__52545\
        );

    \I__13310\ : InMux
    port map (
            O => \N__52618\,
            I => \N__52545\
        );

    \I__13309\ : InMux
    port map (
            O => \N__52617\,
            I => \N__52540\
        );

    \I__13308\ : InMux
    port map (
            O => \N__52616\,
            I => \N__52540\
        );

    \I__13307\ : Span12Mux_h
    port map (
            O => \N__52607\,
            I => \N__52537\
        );

    \I__13306\ : InMux
    port map (
            O => \N__52606\,
            I => \N__52528\
        );

    \I__13305\ : InMux
    port map (
            O => \N__52605\,
            I => \N__52528\
        );

    \I__13304\ : InMux
    port map (
            O => \N__52604\,
            I => \N__52528\
        );

    \I__13303\ : InMux
    port map (
            O => \N__52603\,
            I => \N__52528\
        );

    \I__13302\ : LocalMux
    port map (
            O => \N__52598\,
            I => adc_state_0
        );

    \I__13301\ : LocalMux
    port map (
            O => \N__52595\,
            I => adc_state_0
        );

    \I__13300\ : LocalMux
    port map (
            O => \N__52578\,
            I => adc_state_0
        );

    \I__13299\ : Odrv4
    port map (
            O => \N__52571\,
            I => adc_state_0
        );

    \I__13298\ : Odrv4
    port map (
            O => \N__52564\,
            I => adc_state_0
        );

    \I__13297\ : Odrv4
    port map (
            O => \N__52559\,
            I => adc_state_0
        );

    \I__13296\ : Odrv4
    port map (
            O => \N__52552\,
            I => adc_state_0
        );

    \I__13295\ : LocalMux
    port map (
            O => \N__52545\,
            I => adc_state_0
        );

    \I__13294\ : LocalMux
    port map (
            O => \N__52540\,
            I => adc_state_0
        );

    \I__13293\ : Odrv12
    port map (
            O => \N__52537\,
            I => adc_state_0
        );

    \I__13292\ : LocalMux
    port map (
            O => \N__52528\,
            I => adc_state_0
        );

    \I__13291\ : InMux
    port map (
            O => \N__52505\,
            I => \N__52501\
        );

    \I__13290\ : InMux
    port map (
            O => \N__52504\,
            I => \N__52498\
        );

    \I__13289\ : LocalMux
    port map (
            O => \N__52501\,
            I => \N__52495\
        );

    \I__13288\ : LocalMux
    port map (
            O => \N__52498\,
            I => buf_adcdata1_10
        );

    \I__13287\ : Odrv4
    port map (
            O => \N__52495\,
            I => buf_adcdata1_10
        );

    \I__13286\ : InMux
    port map (
            O => \N__52490\,
            I => \N__52486\
        );

    \I__13285\ : CascadeMux
    port map (
            O => \N__52489\,
            I => \N__52483\
        );

    \I__13284\ : LocalMux
    port map (
            O => \N__52486\,
            I => \N__52480\
        );

    \I__13283\ : InMux
    port map (
            O => \N__52483\,
            I => \N__52477\
        );

    \I__13282\ : Span12Mux_s11_v
    port map (
            O => \N__52480\,
            I => \N__52474\
        );

    \I__13281\ : LocalMux
    port map (
            O => \N__52477\,
            I => n8_adj_1225
        );

    \I__13280\ : Odrv12
    port map (
            O => \N__52474\,
            I => n8_adj_1225
        );

    \I__13279\ : InMux
    port map (
            O => \N__52469\,
            I => \N__52463\
        );

    \I__13278\ : InMux
    port map (
            O => \N__52468\,
            I => \N__52439\
        );

    \I__13277\ : InMux
    port map (
            O => \N__52467\,
            I => \N__52436\
        );

    \I__13276\ : InMux
    port map (
            O => \N__52466\,
            I => \N__52427\
        );

    \I__13275\ : LocalMux
    port map (
            O => \N__52463\,
            I => \N__52420\
        );

    \I__13274\ : CascadeMux
    port map (
            O => \N__52462\,
            I => \N__52415\
        );

    \I__13273\ : CascadeMux
    port map (
            O => \N__52461\,
            I => \N__52411\
        );

    \I__13272\ : CascadeMux
    port map (
            O => \N__52460\,
            I => \N__52407\
        );

    \I__13271\ : CascadeMux
    port map (
            O => \N__52459\,
            I => \N__52403\
        );

    \I__13270\ : CascadeMux
    port map (
            O => \N__52458\,
            I => \N__52399\
        );

    \I__13269\ : CascadeMux
    port map (
            O => \N__52457\,
            I => \N__52395\
        );

    \I__13268\ : CascadeMux
    port map (
            O => \N__52456\,
            I => \N__52391\
        );

    \I__13267\ : InMux
    port map (
            O => \N__52455\,
            I => \N__52387\
        );

    \I__13266\ : CascadeMux
    port map (
            O => \N__52454\,
            I => \N__52381\
        );

    \I__13265\ : InMux
    port map (
            O => \N__52453\,
            I => \N__52377\
        );

    \I__13264\ : InMux
    port map (
            O => \N__52452\,
            I => \N__52369\
        );

    \I__13263\ : InMux
    port map (
            O => \N__52451\,
            I => \N__52369\
        );

    \I__13262\ : InMux
    port map (
            O => \N__52450\,
            I => \N__52369\
        );

    \I__13261\ : InMux
    port map (
            O => \N__52449\,
            I => \N__52364\
        );

    \I__13260\ : InMux
    port map (
            O => \N__52448\,
            I => \N__52364\
        );

    \I__13259\ : CascadeMux
    port map (
            O => \N__52447\,
            I => \N__52361\
        );

    \I__13258\ : CascadeMux
    port map (
            O => \N__52446\,
            I => \N__52357\
        );

    \I__13257\ : InMux
    port map (
            O => \N__52445\,
            I => \N__52351\
        );

    \I__13256\ : InMux
    port map (
            O => \N__52444\,
            I => \N__52351\
        );

    \I__13255\ : InMux
    port map (
            O => \N__52443\,
            I => \N__52346\
        );

    \I__13254\ : InMux
    port map (
            O => \N__52442\,
            I => \N__52342\
        );

    \I__13253\ : LocalMux
    port map (
            O => \N__52439\,
            I => \N__52337\
        );

    \I__13252\ : LocalMux
    port map (
            O => \N__52436\,
            I => \N__52337\
        );

    \I__13251\ : InMux
    port map (
            O => \N__52435\,
            I => \N__52332\
        );

    \I__13250\ : InMux
    port map (
            O => \N__52434\,
            I => \N__52332\
        );

    \I__13249\ : InMux
    port map (
            O => \N__52433\,
            I => \N__52327\
        );

    \I__13248\ : InMux
    port map (
            O => \N__52432\,
            I => \N__52327\
        );

    \I__13247\ : InMux
    port map (
            O => \N__52431\,
            I => \N__52322\
        );

    \I__13246\ : InMux
    port map (
            O => \N__52430\,
            I => \N__52322\
        );

    \I__13245\ : LocalMux
    port map (
            O => \N__52427\,
            I => \N__52319\
        );

    \I__13244\ : InMux
    port map (
            O => \N__52426\,
            I => \N__52314\
        );

    \I__13243\ : InMux
    port map (
            O => \N__52425\,
            I => \N__52314\
        );

    \I__13242\ : SRMux
    port map (
            O => \N__52424\,
            I => \N__52306\
        );

    \I__13241\ : CascadeMux
    port map (
            O => \N__52423\,
            I => \N__52303\
        );

    \I__13240\ : Span4Mux_h
    port map (
            O => \N__52420\,
            I => \N__52297\
        );

    \I__13239\ : InMux
    port map (
            O => \N__52419\,
            I => \N__52280\
        );

    \I__13238\ : InMux
    port map (
            O => \N__52418\,
            I => \N__52280\
        );

    \I__13237\ : InMux
    port map (
            O => \N__52415\,
            I => \N__52280\
        );

    \I__13236\ : InMux
    port map (
            O => \N__52414\,
            I => \N__52280\
        );

    \I__13235\ : InMux
    port map (
            O => \N__52411\,
            I => \N__52280\
        );

    \I__13234\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52280\
        );

    \I__13233\ : InMux
    port map (
            O => \N__52407\,
            I => \N__52280\
        );

    \I__13232\ : InMux
    port map (
            O => \N__52406\,
            I => \N__52280\
        );

    \I__13231\ : InMux
    port map (
            O => \N__52403\,
            I => \N__52265\
        );

    \I__13230\ : InMux
    port map (
            O => \N__52402\,
            I => \N__52265\
        );

    \I__13229\ : InMux
    port map (
            O => \N__52399\,
            I => \N__52265\
        );

    \I__13228\ : InMux
    port map (
            O => \N__52398\,
            I => \N__52265\
        );

    \I__13227\ : InMux
    port map (
            O => \N__52395\,
            I => \N__52265\
        );

    \I__13226\ : InMux
    port map (
            O => \N__52394\,
            I => \N__52265\
        );

    \I__13225\ : InMux
    port map (
            O => \N__52391\,
            I => \N__52265\
        );

    \I__13224\ : CascadeMux
    port map (
            O => \N__52390\,
            I => \N__52262\
        );

    \I__13223\ : LocalMux
    port map (
            O => \N__52387\,
            I => \N__52259\
        );

    \I__13222\ : InMux
    port map (
            O => \N__52386\,
            I => \N__52254\
        );

    \I__13221\ : InMux
    port map (
            O => \N__52385\,
            I => \N__52254\
        );

    \I__13220\ : InMux
    port map (
            O => \N__52384\,
            I => \N__52247\
        );

    \I__13219\ : InMux
    port map (
            O => \N__52381\,
            I => \N__52247\
        );

    \I__13218\ : InMux
    port map (
            O => \N__52380\,
            I => \N__52247\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__52377\,
            I => \N__52244\
        );

    \I__13216\ : InMux
    port map (
            O => \N__52376\,
            I => \N__52241\
        );

    \I__13215\ : LocalMux
    port map (
            O => \N__52369\,
            I => \N__52233\
        );

    \I__13214\ : LocalMux
    port map (
            O => \N__52364\,
            I => \N__52233\
        );

    \I__13213\ : InMux
    port map (
            O => \N__52361\,
            I => \N__52230\
        );

    \I__13212\ : InMux
    port map (
            O => \N__52360\,
            I => \N__52225\
        );

    \I__13211\ : InMux
    port map (
            O => \N__52357\,
            I => \N__52225\
        );

    \I__13210\ : CascadeMux
    port map (
            O => \N__52356\,
            I => \N__52222\
        );

    \I__13209\ : LocalMux
    port map (
            O => \N__52351\,
            I => \N__52214\
        );

    \I__13208\ : InMux
    port map (
            O => \N__52350\,
            I => \N__52211\
        );

    \I__13207\ : InMux
    port map (
            O => \N__52349\,
            I => \N__52208\
        );

    \I__13206\ : LocalMux
    port map (
            O => \N__52346\,
            I => \N__52205\
        );

    \I__13205\ : InMux
    port map (
            O => \N__52345\,
            I => \N__52202\
        );

    \I__13204\ : LocalMux
    port map (
            O => \N__52342\,
            I => \N__52187\
        );

    \I__13203\ : Span4Mux_v
    port map (
            O => \N__52337\,
            I => \N__52187\
        );

    \I__13202\ : LocalMux
    port map (
            O => \N__52332\,
            I => \N__52187\
        );

    \I__13201\ : LocalMux
    port map (
            O => \N__52327\,
            I => \N__52187\
        );

    \I__13200\ : LocalMux
    port map (
            O => \N__52322\,
            I => \N__52187\
        );

    \I__13199\ : Span4Mux_h
    port map (
            O => \N__52319\,
            I => \N__52187\
        );

    \I__13198\ : LocalMux
    port map (
            O => \N__52314\,
            I => \N__52187\
        );

    \I__13197\ : InMux
    port map (
            O => \N__52313\,
            I => \N__52172\
        );

    \I__13196\ : InMux
    port map (
            O => \N__52312\,
            I => \N__52172\
        );

    \I__13195\ : InMux
    port map (
            O => \N__52311\,
            I => \N__52172\
        );

    \I__13194\ : InMux
    port map (
            O => \N__52310\,
            I => \N__52172\
        );

    \I__13193\ : InMux
    port map (
            O => \N__52309\,
            I => \N__52172\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__52306\,
            I => \N__52169\
        );

    \I__13191\ : InMux
    port map (
            O => \N__52303\,
            I => \N__52166\
        );

    \I__13190\ : InMux
    port map (
            O => \N__52302\,
            I => \N__52162\
        );

    \I__13189\ : InMux
    port map (
            O => \N__52301\,
            I => \N__52159\
        );

    \I__13188\ : InMux
    port map (
            O => \N__52300\,
            I => \N__52156\
        );

    \I__13187\ : Span4Mux_v
    port map (
            O => \N__52297\,
            I => \N__52149\
        );

    \I__13186\ : LocalMux
    port map (
            O => \N__52280\,
            I => \N__52149\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__52265\,
            I => \N__52149\
        );

    \I__13184\ : InMux
    port map (
            O => \N__52262\,
            I => \N__52146\
        );

    \I__13183\ : Span4Mux_v
    port map (
            O => \N__52259\,
            I => \N__52143\
        );

    \I__13182\ : LocalMux
    port map (
            O => \N__52254\,
            I => \N__52140\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__52247\,
            I => \N__52133\
        );

    \I__13180\ : Span4Mux_h
    port map (
            O => \N__52244\,
            I => \N__52133\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__52241\,
            I => \N__52133\
        );

    \I__13178\ : InMux
    port map (
            O => \N__52240\,
            I => \N__52126\
        );

    \I__13177\ : InMux
    port map (
            O => \N__52239\,
            I => \N__52126\
        );

    \I__13176\ : InMux
    port map (
            O => \N__52238\,
            I => \N__52126\
        );

    \I__13175\ : Span4Mux_h
    port map (
            O => \N__52233\,
            I => \N__52119\
        );

    \I__13174\ : LocalMux
    port map (
            O => \N__52230\,
            I => \N__52119\
        );

    \I__13173\ : LocalMux
    port map (
            O => \N__52225\,
            I => \N__52119\
        );

    \I__13172\ : InMux
    port map (
            O => \N__52222\,
            I => \N__52110\
        );

    \I__13171\ : InMux
    port map (
            O => \N__52221\,
            I => \N__52110\
        );

    \I__13170\ : InMux
    port map (
            O => \N__52220\,
            I => \N__52110\
        );

    \I__13169\ : InMux
    port map (
            O => \N__52219\,
            I => \N__52110\
        );

    \I__13168\ : InMux
    port map (
            O => \N__52218\,
            I => \N__52105\
        );

    \I__13167\ : InMux
    port map (
            O => \N__52217\,
            I => \N__52105\
        );

    \I__13166\ : Span4Mux_h
    port map (
            O => \N__52214\,
            I => \N__52102\
        );

    \I__13165\ : LocalMux
    port map (
            O => \N__52211\,
            I => \N__52091\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__52208\,
            I => \N__52091\
        );

    \I__13163\ : Span4Mux_h
    port map (
            O => \N__52205\,
            I => \N__52091\
        );

    \I__13162\ : LocalMux
    port map (
            O => \N__52202\,
            I => \N__52091\
        );

    \I__13161\ : Span4Mux_v
    port map (
            O => \N__52187\,
            I => \N__52091\
        );

    \I__13160\ : InMux
    port map (
            O => \N__52186\,
            I => \N__52086\
        );

    \I__13159\ : InMux
    port map (
            O => \N__52185\,
            I => \N__52086\
        );

    \I__13158\ : InMux
    port map (
            O => \N__52184\,
            I => \N__52083\
        );

    \I__13157\ : InMux
    port map (
            O => \N__52183\,
            I => \N__52078\
        );

    \I__13156\ : LocalMux
    port map (
            O => \N__52172\,
            I => \N__52075\
        );

    \I__13155\ : Span4Mux_v
    port map (
            O => \N__52169\,
            I => \N__52070\
        );

    \I__13154\ : LocalMux
    port map (
            O => \N__52166\,
            I => \N__52067\
        );

    \I__13153\ : CascadeMux
    port map (
            O => \N__52165\,
            I => \N__52063\
        );

    \I__13152\ : LocalMux
    port map (
            O => \N__52162\,
            I => \N__52058\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__52159\,
            I => \N__52051\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__52156\,
            I => \N__52051\
        );

    \I__13149\ : Span4Mux_v
    port map (
            O => \N__52149\,
            I => \N__52051\
        );

    \I__13148\ : LocalMux
    port map (
            O => \N__52146\,
            I => \N__52046\
        );

    \I__13147\ : Span4Mux_v
    port map (
            O => \N__52143\,
            I => \N__52046\
        );

    \I__13146\ : Span4Mux_h
    port map (
            O => \N__52140\,
            I => \N__52039\
        );

    \I__13145\ : Span4Mux_v
    port map (
            O => \N__52133\,
            I => \N__52039\
        );

    \I__13144\ : LocalMux
    port map (
            O => \N__52126\,
            I => \N__52039\
        );

    \I__13143\ : Span4Mux_h
    port map (
            O => \N__52119\,
            I => \N__52034\
        );

    \I__13142\ : LocalMux
    port map (
            O => \N__52110\,
            I => \N__52034\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__52105\,
            I => \N__52025\
        );

    \I__13140\ : Span4Mux_h
    port map (
            O => \N__52102\,
            I => \N__52025\
        );

    \I__13139\ : Span4Mux_v
    port map (
            O => \N__52091\,
            I => \N__52025\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__52086\,
            I => \N__52022\
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__52083\,
            I => \N__52019\
        );

    \I__13136\ : InMux
    port map (
            O => \N__52082\,
            I => \N__52016\
        );

    \I__13135\ : InMux
    port map (
            O => \N__52081\,
            I => \N__52013\
        );

    \I__13134\ : LocalMux
    port map (
            O => \N__52078\,
            I => \N__52010\
        );

    \I__13133\ : Span12Mux_v
    port map (
            O => \N__52075\,
            I => \N__52007\
        );

    \I__13132\ : InMux
    port map (
            O => \N__52074\,
            I => \N__52004\
        );

    \I__13131\ : InMux
    port map (
            O => \N__52073\,
            I => \N__52001\
        );

    \I__13130\ : Span4Mux_h
    port map (
            O => \N__52070\,
            I => \N__51996\
        );

    \I__13129\ : Span4Mux_v
    port map (
            O => \N__52067\,
            I => \N__51996\
        );

    \I__13128\ : InMux
    port map (
            O => \N__52066\,
            I => \N__51991\
        );

    \I__13127\ : InMux
    port map (
            O => \N__52063\,
            I => \N__51991\
        );

    \I__13126\ : InMux
    port map (
            O => \N__52062\,
            I => \N__51986\
        );

    \I__13125\ : InMux
    port map (
            O => \N__52061\,
            I => \N__51986\
        );

    \I__13124\ : Span4Mux_v
    port map (
            O => \N__52058\,
            I => \N__51977\
        );

    \I__13123\ : Span4Mux_v
    port map (
            O => \N__52051\,
            I => \N__51977\
        );

    \I__13122\ : Span4Mux_v
    port map (
            O => \N__52046\,
            I => \N__51977\
        );

    \I__13121\ : Span4Mux_h
    port map (
            O => \N__52039\,
            I => \N__51977\
        );

    \I__13120\ : Span4Mux_h
    port map (
            O => \N__52034\,
            I => \N__51974\
        );

    \I__13119\ : InMux
    port map (
            O => \N__52033\,
            I => \N__51969\
        );

    \I__13118\ : InMux
    port map (
            O => \N__52032\,
            I => \N__51969\
        );

    \I__13117\ : Span4Mux_h
    port map (
            O => \N__52025\,
            I => \N__51964\
        );

    \I__13116\ : Span4Mux_h
    port map (
            O => \N__52022\,
            I => \N__51964\
        );

    \I__13115\ : Span12Mux_h
    port map (
            O => \N__52019\,
            I => \N__51953\
        );

    \I__13114\ : LocalMux
    port map (
            O => \N__52016\,
            I => \N__51953\
        );

    \I__13113\ : LocalMux
    port map (
            O => \N__52013\,
            I => \N__51953\
        );

    \I__13112\ : Span12Mux_s10_v
    port map (
            O => \N__52010\,
            I => \N__51953\
        );

    \I__13111\ : Span12Mux_h
    port map (
            O => \N__52007\,
            I => \N__51953\
        );

    \I__13110\ : LocalMux
    port map (
            O => \N__52004\,
            I => comm_state_3
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__52001\,
            I => comm_state_3
        );

    \I__13108\ : Odrv4
    port map (
            O => \N__51996\,
            I => comm_state_3
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__51991\,
            I => comm_state_3
        );

    \I__13106\ : LocalMux
    port map (
            O => \N__51986\,
            I => comm_state_3
        );

    \I__13105\ : Odrv4
    port map (
            O => \N__51977\,
            I => comm_state_3
        );

    \I__13104\ : Odrv4
    port map (
            O => \N__51974\,
            I => comm_state_3
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__51969\,
            I => comm_state_3
        );

    \I__13102\ : Odrv4
    port map (
            O => \N__51964\,
            I => comm_state_3
        );

    \I__13101\ : Odrv12
    port map (
            O => \N__51953\,
            I => comm_state_3
        );

    \I__13100\ : CascadeMux
    port map (
            O => \N__51932\,
            I => \N__51924\
        );

    \I__13099\ : CascadeMux
    port map (
            O => \N__51931\,
            I => \N__51919\
        );

    \I__13098\ : CascadeMux
    port map (
            O => \N__51930\,
            I => \N__51910\
        );

    \I__13097\ : CascadeMux
    port map (
            O => \N__51929\,
            I => \N__51906\
        );

    \I__13096\ : CascadeMux
    port map (
            O => \N__51928\,
            I => \N__51903\
        );

    \I__13095\ : InMux
    port map (
            O => \N__51927\,
            I => \N__51900\
        );

    \I__13094\ : InMux
    port map (
            O => \N__51924\,
            I => \N__51890\
        );

    \I__13093\ : InMux
    port map (
            O => \N__51923\,
            I => \N__51887\
        );

    \I__13092\ : InMux
    port map (
            O => \N__51922\,
            I => \N__51884\
        );

    \I__13091\ : InMux
    port map (
            O => \N__51919\,
            I => \N__51881\
        );

    \I__13090\ : CascadeMux
    port map (
            O => \N__51918\,
            I => \N__51876\
        );

    \I__13089\ : CascadeMux
    port map (
            O => \N__51917\,
            I => \N__51873\
        );

    \I__13088\ : CascadeMux
    port map (
            O => \N__51916\,
            I => \N__51870\
        );

    \I__13087\ : InMux
    port map (
            O => \N__51915\,
            I => \N__51863\
        );

    \I__13086\ : CascadeMux
    port map (
            O => \N__51914\,
            I => \N__51860\
        );

    \I__13085\ : CascadeMux
    port map (
            O => \N__51913\,
            I => \N__51857\
        );

    \I__13084\ : InMux
    port map (
            O => \N__51910\,
            I => \N__51854\
        );

    \I__13083\ : CascadeMux
    port map (
            O => \N__51909\,
            I => \N__51848\
        );

    \I__13082\ : InMux
    port map (
            O => \N__51906\,
            I => \N__51845\
        );

    \I__13081\ : InMux
    port map (
            O => \N__51903\,
            I => \N__51838\
        );

    \I__13080\ : LocalMux
    port map (
            O => \N__51900\,
            I => \N__51835\
        );

    \I__13079\ : InMux
    port map (
            O => \N__51899\,
            I => \N__51830\
        );

    \I__13078\ : InMux
    port map (
            O => \N__51898\,
            I => \N__51830\
        );

    \I__13077\ : CascadeMux
    port map (
            O => \N__51897\,
            I => \N__51826\
        );

    \I__13076\ : InMux
    port map (
            O => \N__51896\,
            I => \N__51822\
        );

    \I__13075\ : InMux
    port map (
            O => \N__51895\,
            I => \N__51817\
        );

    \I__13074\ : InMux
    port map (
            O => \N__51894\,
            I => \N__51817\
        );

    \I__13073\ : InMux
    port map (
            O => \N__51893\,
            I => \N__51814\
        );

    \I__13072\ : LocalMux
    port map (
            O => \N__51890\,
            I => \N__51811\
        );

    \I__13071\ : LocalMux
    port map (
            O => \N__51887\,
            I => \N__51808\
        );

    \I__13070\ : LocalMux
    port map (
            O => \N__51884\,
            I => \N__51805\
        );

    \I__13069\ : LocalMux
    port map (
            O => \N__51881\,
            I => \N__51802\
        );

    \I__13068\ : InMux
    port map (
            O => \N__51880\,
            I => \N__51797\
        );

    \I__13067\ : InMux
    port map (
            O => \N__51879\,
            I => \N__51797\
        );

    \I__13066\ : InMux
    port map (
            O => \N__51876\,
            I => \N__51794\
        );

    \I__13065\ : InMux
    port map (
            O => \N__51873\,
            I => \N__51787\
        );

    \I__13064\ : InMux
    port map (
            O => \N__51870\,
            I => \N__51787\
        );

    \I__13063\ : InMux
    port map (
            O => \N__51869\,
            I => \N__51787\
        );

    \I__13062\ : InMux
    port map (
            O => \N__51868\,
            I => \N__51784\
        );

    \I__13061\ : InMux
    port map (
            O => \N__51867\,
            I => \N__51779\
        );

    \I__13060\ : InMux
    port map (
            O => \N__51866\,
            I => \N__51779\
        );

    \I__13059\ : LocalMux
    port map (
            O => \N__51863\,
            I => \N__51776\
        );

    \I__13058\ : InMux
    port map (
            O => \N__51860\,
            I => \N__51771\
        );

    \I__13057\ : InMux
    port map (
            O => \N__51857\,
            I => \N__51771\
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__51854\,
            I => \N__51763\
        );

    \I__13055\ : InMux
    port map (
            O => \N__51853\,
            I => \N__51758\
        );

    \I__13054\ : InMux
    port map (
            O => \N__51852\,
            I => \N__51758\
        );

    \I__13053\ : InMux
    port map (
            O => \N__51851\,
            I => \N__51753\
        );

    \I__13052\ : InMux
    port map (
            O => \N__51848\,
            I => \N__51753\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__51845\,
            I => \N__51750\
        );

    \I__13050\ : CascadeMux
    port map (
            O => \N__51844\,
            I => \N__51746\
        );

    \I__13049\ : CascadeMux
    port map (
            O => \N__51843\,
            I => \N__51743\
        );

    \I__13048\ : CascadeMux
    port map (
            O => \N__51842\,
            I => \N__51740\
        );

    \I__13047\ : InMux
    port map (
            O => \N__51841\,
            I => \N__51734\
        );

    \I__13046\ : LocalMux
    port map (
            O => \N__51838\,
            I => \N__51731\
        );

    \I__13045\ : Span4Mux_h
    port map (
            O => \N__51835\,
            I => \N__51726\
        );

    \I__13044\ : LocalMux
    port map (
            O => \N__51830\,
            I => \N__51726\
        );

    \I__13043\ : CascadeMux
    port map (
            O => \N__51829\,
            I => \N__51722\
        );

    \I__13042\ : InMux
    port map (
            O => \N__51826\,
            I => \N__51719\
        );

    \I__13041\ : CascadeMux
    port map (
            O => \N__51825\,
            I => \N__51716\
        );

    \I__13040\ : LocalMux
    port map (
            O => \N__51822\,
            I => \N__51711\
        );

    \I__13039\ : LocalMux
    port map (
            O => \N__51817\,
            I => \N__51711\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__51814\,
            I => \N__51708\
        );

    \I__13037\ : Span4Mux_v
    port map (
            O => \N__51811\,
            I => \N__51705\
        );

    \I__13036\ : Span4Mux_v
    port map (
            O => \N__51808\,
            I => \N__51700\
        );

    \I__13035\ : Span4Mux_v
    port map (
            O => \N__51805\,
            I => \N__51700\
        );

    \I__13034\ : Span4Mux_v
    port map (
            O => \N__51802\,
            I => \N__51683\
        );

    \I__13033\ : LocalMux
    port map (
            O => \N__51797\,
            I => \N__51683\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__51794\,
            I => \N__51683\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__51787\,
            I => \N__51683\
        );

    \I__13030\ : LocalMux
    port map (
            O => \N__51784\,
            I => \N__51683\
        );

    \I__13029\ : LocalMux
    port map (
            O => \N__51779\,
            I => \N__51683\
        );

    \I__13028\ : Span4Mux_v
    port map (
            O => \N__51776\,
            I => \N__51683\
        );

    \I__13027\ : LocalMux
    port map (
            O => \N__51771\,
            I => \N__51683\
        );

    \I__13026\ : CascadeMux
    port map (
            O => \N__51770\,
            I => \N__51680\
        );

    \I__13025\ : CascadeMux
    port map (
            O => \N__51769\,
            I => \N__51676\
        );

    \I__13024\ : CascadeMux
    port map (
            O => \N__51768\,
            I => \N__51672\
        );

    \I__13023\ : CascadeMux
    port map (
            O => \N__51767\,
            I => \N__51669\
        );

    \I__13022\ : CascadeMux
    port map (
            O => \N__51766\,
            I => \N__51665\
        );

    \I__13021\ : Span4Mux_h
    port map (
            O => \N__51763\,
            I => \N__51658\
        );

    \I__13020\ : LocalMux
    port map (
            O => \N__51758\,
            I => \N__51658\
        );

    \I__13019\ : LocalMux
    port map (
            O => \N__51753\,
            I => \N__51655\
        );

    \I__13018\ : Span4Mux_v
    port map (
            O => \N__51750\,
            I => \N__51652\
        );

    \I__13017\ : InMux
    port map (
            O => \N__51749\,
            I => \N__51643\
        );

    \I__13016\ : InMux
    port map (
            O => \N__51746\,
            I => \N__51643\
        );

    \I__13015\ : InMux
    port map (
            O => \N__51743\,
            I => \N__51643\
        );

    \I__13014\ : InMux
    port map (
            O => \N__51740\,
            I => \N__51643\
        );

    \I__13013\ : CascadeMux
    port map (
            O => \N__51739\,
            I => \N__51640\
        );

    \I__13012\ : CascadeMux
    port map (
            O => \N__51738\,
            I => \N__51637\
        );

    \I__13011\ : CascadeMux
    port map (
            O => \N__51737\,
            I => \N__51633\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__51734\,
            I => \N__51630\
        );

    \I__13009\ : Span4Mux_h
    port map (
            O => \N__51731\,
            I => \N__51625\
        );

    \I__13008\ : Span4Mux_h
    port map (
            O => \N__51726\,
            I => \N__51625\
        );

    \I__13007\ : InMux
    port map (
            O => \N__51725\,
            I => \N__51620\
        );

    \I__13006\ : InMux
    port map (
            O => \N__51722\,
            I => \N__51620\
        );

    \I__13005\ : LocalMux
    port map (
            O => \N__51719\,
            I => \N__51617\
        );

    \I__13004\ : InMux
    port map (
            O => \N__51716\,
            I => \N__51614\
        );

    \I__13003\ : Span4Mux_v
    port map (
            O => \N__51711\,
            I => \N__51607\
        );

    \I__13002\ : Span4Mux_v
    port map (
            O => \N__51708\,
            I => \N__51607\
        );

    \I__13001\ : Span4Mux_v
    port map (
            O => \N__51705\,
            I => \N__51607\
        );

    \I__13000\ : Span4Mux_v
    port map (
            O => \N__51700\,
            I => \N__51602\
        );

    \I__12999\ : Span4Mux_v
    port map (
            O => \N__51683\,
            I => \N__51602\
        );

    \I__12998\ : InMux
    port map (
            O => \N__51680\,
            I => \N__51599\
        );

    \I__12997\ : InMux
    port map (
            O => \N__51679\,
            I => \N__51594\
        );

    \I__12996\ : InMux
    port map (
            O => \N__51676\,
            I => \N__51594\
        );

    \I__12995\ : InMux
    port map (
            O => \N__51675\,
            I => \N__51583\
        );

    \I__12994\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51583\
        );

    \I__12993\ : InMux
    port map (
            O => \N__51669\,
            I => \N__51583\
        );

    \I__12992\ : InMux
    port map (
            O => \N__51668\,
            I => \N__51583\
        );

    \I__12991\ : InMux
    port map (
            O => \N__51665\,
            I => \N__51583\
        );

    \I__12990\ : InMux
    port map (
            O => \N__51664\,
            I => \N__51578\
        );

    \I__12989\ : InMux
    port map (
            O => \N__51663\,
            I => \N__51578\
        );

    \I__12988\ : Span4Mux_h
    port map (
            O => \N__51658\,
            I => \N__51569\
        );

    \I__12987\ : Span4Mux_v
    port map (
            O => \N__51655\,
            I => \N__51569\
        );

    \I__12986\ : Span4Mux_h
    port map (
            O => \N__51652\,
            I => \N__51569\
        );

    \I__12985\ : LocalMux
    port map (
            O => \N__51643\,
            I => \N__51569\
        );

    \I__12984\ : InMux
    port map (
            O => \N__51640\,
            I => \N__51566\
        );

    \I__12983\ : InMux
    port map (
            O => \N__51637\,
            I => \N__51561\
        );

    \I__12982\ : InMux
    port map (
            O => \N__51636\,
            I => \N__51561\
        );

    \I__12981\ : InMux
    port map (
            O => \N__51633\,
            I => \N__51558\
        );

    \I__12980\ : Span12Mux_v
    port map (
            O => \N__51630\,
            I => \N__51555\
        );

    \I__12979\ : Span4Mux_v
    port map (
            O => \N__51625\,
            I => \N__51550\
        );

    \I__12978\ : LocalMux
    port map (
            O => \N__51620\,
            I => \N__51550\
        );

    \I__12977\ : Span12Mux_v
    port map (
            O => \N__51617\,
            I => \N__51541\
        );

    \I__12976\ : LocalMux
    port map (
            O => \N__51614\,
            I => \N__51541\
        );

    \I__12975\ : Sp12to4
    port map (
            O => \N__51607\,
            I => \N__51541\
        );

    \I__12974\ : Sp12to4
    port map (
            O => \N__51602\,
            I => \N__51541\
        );

    \I__12973\ : LocalMux
    port map (
            O => \N__51599\,
            I => \N__51530\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__51594\,
            I => \N__51530\
        );

    \I__12971\ : LocalMux
    port map (
            O => \N__51583\,
            I => \N__51530\
        );

    \I__12970\ : LocalMux
    port map (
            O => \N__51578\,
            I => \N__51530\
        );

    \I__12969\ : Span4Mux_v
    port map (
            O => \N__51569\,
            I => \N__51530\
        );

    \I__12968\ : LocalMux
    port map (
            O => \N__51566\,
            I => n6791
        );

    \I__12967\ : LocalMux
    port map (
            O => \N__51561\,
            I => n6791
        );

    \I__12966\ : LocalMux
    port map (
            O => \N__51558\,
            I => n6791
        );

    \I__12965\ : Odrv12
    port map (
            O => \N__51555\,
            I => n6791
        );

    \I__12964\ : Odrv4
    port map (
            O => \N__51550\,
            I => n6791
        );

    \I__12963\ : Odrv12
    port map (
            O => \N__51541\,
            I => n6791
        );

    \I__12962\ : Odrv4
    port map (
            O => \N__51530\,
            I => n6791
        );

    \I__12961\ : InMux
    port map (
            O => \N__51515\,
            I => \N__51512\
        );

    \I__12960\ : LocalMux
    port map (
            O => \N__51512\,
            I => \N__51509\
        );

    \I__12959\ : Span4Mux_h
    port map (
            O => \N__51509\,
            I => \N__51505\
        );

    \I__12958\ : InMux
    port map (
            O => \N__51508\,
            I => \N__51502\
        );

    \I__12957\ : Span4Mux_h
    port map (
            O => \N__51505\,
            I => \N__51499\
        );

    \I__12956\ : LocalMux
    port map (
            O => \N__51502\,
            I => n7_adj_1224
        );

    \I__12955\ : Odrv4
    port map (
            O => \N__51499\,
            I => n7_adj_1224
        );

    \I__12954\ : CascadeMux
    port map (
            O => \N__51494\,
            I => \N__51491\
        );

    \I__12953\ : CascadeBuf
    port map (
            O => \N__51491\,
            I => \N__51488\
        );

    \I__12952\ : CascadeMux
    port map (
            O => \N__51488\,
            I => \N__51485\
        );

    \I__12951\ : CascadeBuf
    port map (
            O => \N__51485\,
            I => \N__51482\
        );

    \I__12950\ : CascadeMux
    port map (
            O => \N__51482\,
            I => \N__51479\
        );

    \I__12949\ : CascadeBuf
    port map (
            O => \N__51479\,
            I => \N__51476\
        );

    \I__12948\ : CascadeMux
    port map (
            O => \N__51476\,
            I => \N__51473\
        );

    \I__12947\ : CascadeBuf
    port map (
            O => \N__51473\,
            I => \N__51470\
        );

    \I__12946\ : CascadeMux
    port map (
            O => \N__51470\,
            I => \N__51467\
        );

    \I__12945\ : CascadeBuf
    port map (
            O => \N__51467\,
            I => \N__51464\
        );

    \I__12944\ : CascadeMux
    port map (
            O => \N__51464\,
            I => \N__51461\
        );

    \I__12943\ : CascadeBuf
    port map (
            O => \N__51461\,
            I => \N__51457\
        );

    \I__12942\ : CascadeMux
    port map (
            O => \N__51460\,
            I => \N__51454\
        );

    \I__12941\ : CascadeMux
    port map (
            O => \N__51457\,
            I => \N__51451\
        );

    \I__12940\ : CascadeBuf
    port map (
            O => \N__51454\,
            I => \N__51448\
        );

    \I__12939\ : CascadeBuf
    port map (
            O => \N__51451\,
            I => \N__51445\
        );

    \I__12938\ : CascadeMux
    port map (
            O => \N__51448\,
            I => \N__51442\
        );

    \I__12937\ : CascadeMux
    port map (
            O => \N__51445\,
            I => \N__51439\
        );

    \I__12936\ : InMux
    port map (
            O => \N__51442\,
            I => \N__51436\
        );

    \I__12935\ : CascadeBuf
    port map (
            O => \N__51439\,
            I => \N__51433\
        );

    \I__12934\ : LocalMux
    port map (
            O => \N__51436\,
            I => \N__51430\
        );

    \I__12933\ : CascadeMux
    port map (
            O => \N__51433\,
            I => \N__51427\
        );

    \I__12932\ : Span12Mux_s11_h
    port map (
            O => \N__51430\,
            I => \N__51424\
        );

    \I__12931\ : CascadeBuf
    port map (
            O => \N__51427\,
            I => \N__51421\
        );

    \I__12930\ : Span12Mux_h
    port map (
            O => \N__51424\,
            I => \N__51418\
        );

    \I__12929\ : CascadeMux
    port map (
            O => \N__51421\,
            I => \N__51415\
        );

    \I__12928\ : Span12Mux_v
    port map (
            O => \N__51418\,
            I => \N__51412\
        );

    \I__12927\ : InMux
    port map (
            O => \N__51415\,
            I => \N__51409\
        );

    \I__12926\ : Odrv12
    port map (
            O => \N__51412\,
            I => \data_index_9_N_258_5\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__51409\,
            I => \data_index_9_N_258_5\
        );

    \I__12924\ : InMux
    port map (
            O => \N__51404\,
            I => \N__51401\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__51401\,
            I => \N__51398\
        );

    \I__12922\ : Span4Mux_v
    port map (
            O => \N__51398\,
            I => \N__51394\
        );

    \I__12921\ : InMux
    port map (
            O => \N__51397\,
            I => \N__51391\
        );

    \I__12920\ : Span4Mux_h
    port map (
            O => \N__51394\,
            I => \N__51385\
        );

    \I__12919\ : LocalMux
    port map (
            O => \N__51391\,
            I => \N__51385\
        );

    \I__12918\ : InMux
    port map (
            O => \N__51390\,
            I => \N__51382\
        );

    \I__12917\ : Span4Mux_v
    port map (
            O => \N__51385\,
            I => \N__51379\
        );

    \I__12916\ : LocalMux
    port map (
            O => \N__51382\,
            I => \N__51376\
        );

    \I__12915\ : Span4Mux_h
    port map (
            O => \N__51379\,
            I => \N__51371\
        );

    \I__12914\ : Span4Mux_h
    port map (
            O => \N__51376\,
            I => \N__51368\
        );

    \I__12913\ : InMux
    port map (
            O => \N__51375\,
            I => \N__51365\
        );

    \I__12912\ : InMux
    port map (
            O => \N__51374\,
            I => \N__51362\
        );

    \I__12911\ : Sp12to4
    port map (
            O => \N__51371\,
            I => \N__51359\
        );

    \I__12910\ : Span4Mux_h
    port map (
            O => \N__51368\,
            I => \N__51354\
        );

    \I__12909\ : LocalMux
    port map (
            O => \N__51365\,
            I => \N__51354\
        );

    \I__12908\ : LocalMux
    port map (
            O => \N__51362\,
            I => \N__51351\
        );

    \I__12907\ : Span12Mux_s4_h
    port map (
            O => \N__51359\,
            I => \N__51346\
        );

    \I__12906\ : Sp12to4
    port map (
            O => \N__51354\,
            I => \N__51346\
        );

    \I__12905\ : Span12Mux_v
    port map (
            O => \N__51351\,
            I => \N__51343\
        );

    \I__12904\ : Span12Mux_v
    port map (
            O => \N__51346\,
            I => \N__51340\
        );

    \I__12903\ : Odrv12
    port map (
            O => \N__51343\,
            I => \ICE_SPI_SCLK\
        );

    \I__12902\ : Odrv12
    port map (
            O => \N__51340\,
            I => \ICE_SPI_SCLK\
        );

    \I__12901\ : InMux
    port map (
            O => \N__51335\,
            I => \N__51332\
        );

    \I__12900\ : LocalMux
    port map (
            O => \N__51332\,
            I => \N__51329\
        );

    \I__12899\ : Span4Mux_v
    port map (
            O => \N__51329\,
            I => \N__51326\
        );

    \I__12898\ : Span4Mux_h
    port map (
            O => \N__51326\,
            I => \N__51323\
        );

    \I__12897\ : Odrv4
    port map (
            O => \N__51323\,
            I => \comm_spi.n10437\
        );

    \I__12896\ : ClkMux
    port map (
            O => \N__51320\,
            I => \N__50675\
        );

    \I__12895\ : ClkMux
    port map (
            O => \N__51319\,
            I => \N__50675\
        );

    \I__12894\ : ClkMux
    port map (
            O => \N__51318\,
            I => \N__50675\
        );

    \I__12893\ : ClkMux
    port map (
            O => \N__51317\,
            I => \N__50675\
        );

    \I__12892\ : ClkMux
    port map (
            O => \N__51316\,
            I => \N__50675\
        );

    \I__12891\ : ClkMux
    port map (
            O => \N__51315\,
            I => \N__50675\
        );

    \I__12890\ : ClkMux
    port map (
            O => \N__51314\,
            I => \N__50675\
        );

    \I__12889\ : ClkMux
    port map (
            O => \N__51313\,
            I => \N__50675\
        );

    \I__12888\ : ClkMux
    port map (
            O => \N__51312\,
            I => \N__50675\
        );

    \I__12887\ : ClkMux
    port map (
            O => \N__51311\,
            I => \N__50675\
        );

    \I__12886\ : ClkMux
    port map (
            O => \N__51310\,
            I => \N__50675\
        );

    \I__12885\ : ClkMux
    port map (
            O => \N__51309\,
            I => \N__50675\
        );

    \I__12884\ : ClkMux
    port map (
            O => \N__51308\,
            I => \N__50675\
        );

    \I__12883\ : ClkMux
    port map (
            O => \N__51307\,
            I => \N__50675\
        );

    \I__12882\ : ClkMux
    port map (
            O => \N__51306\,
            I => \N__50675\
        );

    \I__12881\ : ClkMux
    port map (
            O => \N__51305\,
            I => \N__50675\
        );

    \I__12880\ : ClkMux
    port map (
            O => \N__51304\,
            I => \N__50675\
        );

    \I__12879\ : ClkMux
    port map (
            O => \N__51303\,
            I => \N__50675\
        );

    \I__12878\ : ClkMux
    port map (
            O => \N__51302\,
            I => \N__50675\
        );

    \I__12877\ : ClkMux
    port map (
            O => \N__51301\,
            I => \N__50675\
        );

    \I__12876\ : ClkMux
    port map (
            O => \N__51300\,
            I => \N__50675\
        );

    \I__12875\ : ClkMux
    port map (
            O => \N__51299\,
            I => \N__50675\
        );

    \I__12874\ : ClkMux
    port map (
            O => \N__51298\,
            I => \N__50675\
        );

    \I__12873\ : ClkMux
    port map (
            O => \N__51297\,
            I => \N__50675\
        );

    \I__12872\ : ClkMux
    port map (
            O => \N__51296\,
            I => \N__50675\
        );

    \I__12871\ : ClkMux
    port map (
            O => \N__51295\,
            I => \N__50675\
        );

    \I__12870\ : ClkMux
    port map (
            O => \N__51294\,
            I => \N__50675\
        );

    \I__12869\ : ClkMux
    port map (
            O => \N__51293\,
            I => \N__50675\
        );

    \I__12868\ : ClkMux
    port map (
            O => \N__51292\,
            I => \N__50675\
        );

    \I__12867\ : ClkMux
    port map (
            O => \N__51291\,
            I => \N__50675\
        );

    \I__12866\ : ClkMux
    port map (
            O => \N__51290\,
            I => \N__50675\
        );

    \I__12865\ : ClkMux
    port map (
            O => \N__51289\,
            I => \N__50675\
        );

    \I__12864\ : ClkMux
    port map (
            O => \N__51288\,
            I => \N__50675\
        );

    \I__12863\ : ClkMux
    port map (
            O => \N__51287\,
            I => \N__50675\
        );

    \I__12862\ : ClkMux
    port map (
            O => \N__51286\,
            I => \N__50675\
        );

    \I__12861\ : ClkMux
    port map (
            O => \N__51285\,
            I => \N__50675\
        );

    \I__12860\ : ClkMux
    port map (
            O => \N__51284\,
            I => \N__50675\
        );

    \I__12859\ : ClkMux
    port map (
            O => \N__51283\,
            I => \N__50675\
        );

    \I__12858\ : ClkMux
    port map (
            O => \N__51282\,
            I => \N__50675\
        );

    \I__12857\ : ClkMux
    port map (
            O => \N__51281\,
            I => \N__50675\
        );

    \I__12856\ : ClkMux
    port map (
            O => \N__51280\,
            I => \N__50675\
        );

    \I__12855\ : ClkMux
    port map (
            O => \N__51279\,
            I => \N__50675\
        );

    \I__12854\ : ClkMux
    port map (
            O => \N__51278\,
            I => \N__50675\
        );

    \I__12853\ : ClkMux
    port map (
            O => \N__51277\,
            I => \N__50675\
        );

    \I__12852\ : ClkMux
    port map (
            O => \N__51276\,
            I => \N__50675\
        );

    \I__12851\ : ClkMux
    port map (
            O => \N__51275\,
            I => \N__50675\
        );

    \I__12850\ : ClkMux
    port map (
            O => \N__51274\,
            I => \N__50675\
        );

    \I__12849\ : ClkMux
    port map (
            O => \N__51273\,
            I => \N__50675\
        );

    \I__12848\ : ClkMux
    port map (
            O => \N__51272\,
            I => \N__50675\
        );

    \I__12847\ : ClkMux
    port map (
            O => \N__51271\,
            I => \N__50675\
        );

    \I__12846\ : ClkMux
    port map (
            O => \N__51270\,
            I => \N__50675\
        );

    \I__12845\ : ClkMux
    port map (
            O => \N__51269\,
            I => \N__50675\
        );

    \I__12844\ : ClkMux
    port map (
            O => \N__51268\,
            I => \N__50675\
        );

    \I__12843\ : ClkMux
    port map (
            O => \N__51267\,
            I => \N__50675\
        );

    \I__12842\ : ClkMux
    port map (
            O => \N__51266\,
            I => \N__50675\
        );

    \I__12841\ : ClkMux
    port map (
            O => \N__51265\,
            I => \N__50675\
        );

    \I__12840\ : ClkMux
    port map (
            O => \N__51264\,
            I => \N__50675\
        );

    \I__12839\ : ClkMux
    port map (
            O => \N__51263\,
            I => \N__50675\
        );

    \I__12838\ : ClkMux
    port map (
            O => \N__51262\,
            I => \N__50675\
        );

    \I__12837\ : ClkMux
    port map (
            O => \N__51261\,
            I => \N__50675\
        );

    \I__12836\ : ClkMux
    port map (
            O => \N__51260\,
            I => \N__50675\
        );

    \I__12835\ : ClkMux
    port map (
            O => \N__51259\,
            I => \N__50675\
        );

    \I__12834\ : ClkMux
    port map (
            O => \N__51258\,
            I => \N__50675\
        );

    \I__12833\ : ClkMux
    port map (
            O => \N__51257\,
            I => \N__50675\
        );

    \I__12832\ : ClkMux
    port map (
            O => \N__51256\,
            I => \N__50675\
        );

    \I__12831\ : ClkMux
    port map (
            O => \N__51255\,
            I => \N__50675\
        );

    \I__12830\ : ClkMux
    port map (
            O => \N__51254\,
            I => \N__50675\
        );

    \I__12829\ : ClkMux
    port map (
            O => \N__51253\,
            I => \N__50675\
        );

    \I__12828\ : ClkMux
    port map (
            O => \N__51252\,
            I => \N__50675\
        );

    \I__12827\ : ClkMux
    port map (
            O => \N__51251\,
            I => \N__50675\
        );

    \I__12826\ : ClkMux
    port map (
            O => \N__51250\,
            I => \N__50675\
        );

    \I__12825\ : ClkMux
    port map (
            O => \N__51249\,
            I => \N__50675\
        );

    \I__12824\ : ClkMux
    port map (
            O => \N__51248\,
            I => \N__50675\
        );

    \I__12823\ : ClkMux
    port map (
            O => \N__51247\,
            I => \N__50675\
        );

    \I__12822\ : ClkMux
    port map (
            O => \N__51246\,
            I => \N__50675\
        );

    \I__12821\ : ClkMux
    port map (
            O => \N__51245\,
            I => \N__50675\
        );

    \I__12820\ : ClkMux
    port map (
            O => \N__51244\,
            I => \N__50675\
        );

    \I__12819\ : ClkMux
    port map (
            O => \N__51243\,
            I => \N__50675\
        );

    \I__12818\ : ClkMux
    port map (
            O => \N__51242\,
            I => \N__50675\
        );

    \I__12817\ : ClkMux
    port map (
            O => \N__51241\,
            I => \N__50675\
        );

    \I__12816\ : ClkMux
    port map (
            O => \N__51240\,
            I => \N__50675\
        );

    \I__12815\ : ClkMux
    port map (
            O => \N__51239\,
            I => \N__50675\
        );

    \I__12814\ : ClkMux
    port map (
            O => \N__51238\,
            I => \N__50675\
        );

    \I__12813\ : ClkMux
    port map (
            O => \N__51237\,
            I => \N__50675\
        );

    \I__12812\ : ClkMux
    port map (
            O => \N__51236\,
            I => \N__50675\
        );

    \I__12811\ : ClkMux
    port map (
            O => \N__51235\,
            I => \N__50675\
        );

    \I__12810\ : ClkMux
    port map (
            O => \N__51234\,
            I => \N__50675\
        );

    \I__12809\ : ClkMux
    port map (
            O => \N__51233\,
            I => \N__50675\
        );

    \I__12808\ : ClkMux
    port map (
            O => \N__51232\,
            I => \N__50675\
        );

    \I__12807\ : ClkMux
    port map (
            O => \N__51231\,
            I => \N__50675\
        );

    \I__12806\ : ClkMux
    port map (
            O => \N__51230\,
            I => \N__50675\
        );

    \I__12805\ : ClkMux
    port map (
            O => \N__51229\,
            I => \N__50675\
        );

    \I__12804\ : ClkMux
    port map (
            O => \N__51228\,
            I => \N__50675\
        );

    \I__12803\ : ClkMux
    port map (
            O => \N__51227\,
            I => \N__50675\
        );

    \I__12802\ : ClkMux
    port map (
            O => \N__51226\,
            I => \N__50675\
        );

    \I__12801\ : ClkMux
    port map (
            O => \N__51225\,
            I => \N__50675\
        );

    \I__12800\ : ClkMux
    port map (
            O => \N__51224\,
            I => \N__50675\
        );

    \I__12799\ : ClkMux
    port map (
            O => \N__51223\,
            I => \N__50675\
        );

    \I__12798\ : ClkMux
    port map (
            O => \N__51222\,
            I => \N__50675\
        );

    \I__12797\ : ClkMux
    port map (
            O => \N__51221\,
            I => \N__50675\
        );

    \I__12796\ : ClkMux
    port map (
            O => \N__51220\,
            I => \N__50675\
        );

    \I__12795\ : ClkMux
    port map (
            O => \N__51219\,
            I => \N__50675\
        );

    \I__12794\ : ClkMux
    port map (
            O => \N__51218\,
            I => \N__50675\
        );

    \I__12793\ : ClkMux
    port map (
            O => \N__51217\,
            I => \N__50675\
        );

    \I__12792\ : ClkMux
    port map (
            O => \N__51216\,
            I => \N__50675\
        );

    \I__12791\ : ClkMux
    port map (
            O => \N__51215\,
            I => \N__50675\
        );

    \I__12790\ : ClkMux
    port map (
            O => \N__51214\,
            I => \N__50675\
        );

    \I__12789\ : ClkMux
    port map (
            O => \N__51213\,
            I => \N__50675\
        );

    \I__12788\ : ClkMux
    port map (
            O => \N__51212\,
            I => \N__50675\
        );

    \I__12787\ : ClkMux
    port map (
            O => \N__51211\,
            I => \N__50675\
        );

    \I__12786\ : ClkMux
    port map (
            O => \N__51210\,
            I => \N__50675\
        );

    \I__12785\ : ClkMux
    port map (
            O => \N__51209\,
            I => \N__50675\
        );

    \I__12784\ : ClkMux
    port map (
            O => \N__51208\,
            I => \N__50675\
        );

    \I__12783\ : ClkMux
    port map (
            O => \N__51207\,
            I => \N__50675\
        );

    \I__12782\ : ClkMux
    port map (
            O => \N__51206\,
            I => \N__50675\
        );

    \I__12781\ : ClkMux
    port map (
            O => \N__51205\,
            I => \N__50675\
        );

    \I__12780\ : ClkMux
    port map (
            O => \N__51204\,
            I => \N__50675\
        );

    \I__12779\ : ClkMux
    port map (
            O => \N__51203\,
            I => \N__50675\
        );

    \I__12778\ : ClkMux
    port map (
            O => \N__51202\,
            I => \N__50675\
        );

    \I__12777\ : ClkMux
    port map (
            O => \N__51201\,
            I => \N__50675\
        );

    \I__12776\ : ClkMux
    port map (
            O => \N__51200\,
            I => \N__50675\
        );

    \I__12775\ : ClkMux
    port map (
            O => \N__51199\,
            I => \N__50675\
        );

    \I__12774\ : ClkMux
    port map (
            O => \N__51198\,
            I => \N__50675\
        );

    \I__12773\ : ClkMux
    port map (
            O => \N__51197\,
            I => \N__50675\
        );

    \I__12772\ : ClkMux
    port map (
            O => \N__51196\,
            I => \N__50675\
        );

    \I__12771\ : ClkMux
    port map (
            O => \N__51195\,
            I => \N__50675\
        );

    \I__12770\ : ClkMux
    port map (
            O => \N__51194\,
            I => \N__50675\
        );

    \I__12769\ : ClkMux
    port map (
            O => \N__51193\,
            I => \N__50675\
        );

    \I__12768\ : ClkMux
    port map (
            O => \N__51192\,
            I => \N__50675\
        );

    \I__12767\ : ClkMux
    port map (
            O => \N__51191\,
            I => \N__50675\
        );

    \I__12766\ : ClkMux
    port map (
            O => \N__51190\,
            I => \N__50675\
        );

    \I__12765\ : ClkMux
    port map (
            O => \N__51189\,
            I => \N__50675\
        );

    \I__12764\ : ClkMux
    port map (
            O => \N__51188\,
            I => \N__50675\
        );

    \I__12763\ : ClkMux
    port map (
            O => \N__51187\,
            I => \N__50675\
        );

    \I__12762\ : ClkMux
    port map (
            O => \N__51186\,
            I => \N__50675\
        );

    \I__12761\ : ClkMux
    port map (
            O => \N__51185\,
            I => \N__50675\
        );

    \I__12760\ : ClkMux
    port map (
            O => \N__51184\,
            I => \N__50675\
        );

    \I__12759\ : ClkMux
    port map (
            O => \N__51183\,
            I => \N__50675\
        );

    \I__12758\ : ClkMux
    port map (
            O => \N__51182\,
            I => \N__50675\
        );

    \I__12757\ : ClkMux
    port map (
            O => \N__51181\,
            I => \N__50675\
        );

    \I__12756\ : ClkMux
    port map (
            O => \N__51180\,
            I => \N__50675\
        );

    \I__12755\ : ClkMux
    port map (
            O => \N__51179\,
            I => \N__50675\
        );

    \I__12754\ : ClkMux
    port map (
            O => \N__51178\,
            I => \N__50675\
        );

    \I__12753\ : ClkMux
    port map (
            O => \N__51177\,
            I => \N__50675\
        );

    \I__12752\ : ClkMux
    port map (
            O => \N__51176\,
            I => \N__50675\
        );

    \I__12751\ : ClkMux
    port map (
            O => \N__51175\,
            I => \N__50675\
        );

    \I__12750\ : ClkMux
    port map (
            O => \N__51174\,
            I => \N__50675\
        );

    \I__12749\ : ClkMux
    port map (
            O => \N__51173\,
            I => \N__50675\
        );

    \I__12748\ : ClkMux
    port map (
            O => \N__51172\,
            I => \N__50675\
        );

    \I__12747\ : ClkMux
    port map (
            O => \N__51171\,
            I => \N__50675\
        );

    \I__12746\ : ClkMux
    port map (
            O => \N__51170\,
            I => \N__50675\
        );

    \I__12745\ : ClkMux
    port map (
            O => \N__51169\,
            I => \N__50675\
        );

    \I__12744\ : ClkMux
    port map (
            O => \N__51168\,
            I => \N__50675\
        );

    \I__12743\ : ClkMux
    port map (
            O => \N__51167\,
            I => \N__50675\
        );

    \I__12742\ : ClkMux
    port map (
            O => \N__51166\,
            I => \N__50675\
        );

    \I__12741\ : ClkMux
    port map (
            O => \N__51165\,
            I => \N__50675\
        );

    \I__12740\ : ClkMux
    port map (
            O => \N__51164\,
            I => \N__50675\
        );

    \I__12739\ : ClkMux
    port map (
            O => \N__51163\,
            I => \N__50675\
        );

    \I__12738\ : ClkMux
    port map (
            O => \N__51162\,
            I => \N__50675\
        );

    \I__12737\ : ClkMux
    port map (
            O => \N__51161\,
            I => \N__50675\
        );

    \I__12736\ : ClkMux
    port map (
            O => \N__51160\,
            I => \N__50675\
        );

    \I__12735\ : ClkMux
    port map (
            O => \N__51159\,
            I => \N__50675\
        );

    \I__12734\ : ClkMux
    port map (
            O => \N__51158\,
            I => \N__50675\
        );

    \I__12733\ : ClkMux
    port map (
            O => \N__51157\,
            I => \N__50675\
        );

    \I__12732\ : ClkMux
    port map (
            O => \N__51156\,
            I => \N__50675\
        );

    \I__12731\ : ClkMux
    port map (
            O => \N__51155\,
            I => \N__50675\
        );

    \I__12730\ : ClkMux
    port map (
            O => \N__51154\,
            I => \N__50675\
        );

    \I__12729\ : ClkMux
    port map (
            O => \N__51153\,
            I => \N__50675\
        );

    \I__12728\ : ClkMux
    port map (
            O => \N__51152\,
            I => \N__50675\
        );

    \I__12727\ : ClkMux
    port map (
            O => \N__51151\,
            I => \N__50675\
        );

    \I__12726\ : ClkMux
    port map (
            O => \N__51150\,
            I => \N__50675\
        );

    \I__12725\ : ClkMux
    port map (
            O => \N__51149\,
            I => \N__50675\
        );

    \I__12724\ : ClkMux
    port map (
            O => \N__51148\,
            I => \N__50675\
        );

    \I__12723\ : ClkMux
    port map (
            O => \N__51147\,
            I => \N__50675\
        );

    \I__12722\ : ClkMux
    port map (
            O => \N__51146\,
            I => \N__50675\
        );

    \I__12721\ : ClkMux
    port map (
            O => \N__51145\,
            I => \N__50675\
        );

    \I__12720\ : ClkMux
    port map (
            O => \N__51144\,
            I => \N__50675\
        );

    \I__12719\ : ClkMux
    port map (
            O => \N__51143\,
            I => \N__50675\
        );

    \I__12718\ : ClkMux
    port map (
            O => \N__51142\,
            I => \N__50675\
        );

    \I__12717\ : ClkMux
    port map (
            O => \N__51141\,
            I => \N__50675\
        );

    \I__12716\ : ClkMux
    port map (
            O => \N__51140\,
            I => \N__50675\
        );

    \I__12715\ : ClkMux
    port map (
            O => \N__51139\,
            I => \N__50675\
        );

    \I__12714\ : ClkMux
    port map (
            O => \N__51138\,
            I => \N__50675\
        );

    \I__12713\ : ClkMux
    port map (
            O => \N__51137\,
            I => \N__50675\
        );

    \I__12712\ : ClkMux
    port map (
            O => \N__51136\,
            I => \N__50675\
        );

    \I__12711\ : ClkMux
    port map (
            O => \N__51135\,
            I => \N__50675\
        );

    \I__12710\ : ClkMux
    port map (
            O => \N__51134\,
            I => \N__50675\
        );

    \I__12709\ : ClkMux
    port map (
            O => \N__51133\,
            I => \N__50675\
        );

    \I__12708\ : ClkMux
    port map (
            O => \N__51132\,
            I => \N__50675\
        );

    \I__12707\ : ClkMux
    port map (
            O => \N__51131\,
            I => \N__50675\
        );

    \I__12706\ : ClkMux
    port map (
            O => \N__51130\,
            I => \N__50675\
        );

    \I__12705\ : ClkMux
    port map (
            O => \N__51129\,
            I => \N__50675\
        );

    \I__12704\ : ClkMux
    port map (
            O => \N__51128\,
            I => \N__50675\
        );

    \I__12703\ : ClkMux
    port map (
            O => \N__51127\,
            I => \N__50675\
        );

    \I__12702\ : ClkMux
    port map (
            O => \N__51126\,
            I => \N__50675\
        );

    \I__12701\ : ClkMux
    port map (
            O => \N__51125\,
            I => \N__50675\
        );

    \I__12700\ : ClkMux
    port map (
            O => \N__51124\,
            I => \N__50675\
        );

    \I__12699\ : ClkMux
    port map (
            O => \N__51123\,
            I => \N__50675\
        );

    \I__12698\ : ClkMux
    port map (
            O => \N__51122\,
            I => \N__50675\
        );

    \I__12697\ : ClkMux
    port map (
            O => \N__51121\,
            I => \N__50675\
        );

    \I__12696\ : ClkMux
    port map (
            O => \N__51120\,
            I => \N__50675\
        );

    \I__12695\ : ClkMux
    port map (
            O => \N__51119\,
            I => \N__50675\
        );

    \I__12694\ : ClkMux
    port map (
            O => \N__51118\,
            I => \N__50675\
        );

    \I__12693\ : ClkMux
    port map (
            O => \N__51117\,
            I => \N__50675\
        );

    \I__12692\ : ClkMux
    port map (
            O => \N__51116\,
            I => \N__50675\
        );

    \I__12691\ : ClkMux
    port map (
            O => \N__51115\,
            I => \N__50675\
        );

    \I__12690\ : ClkMux
    port map (
            O => \N__51114\,
            I => \N__50675\
        );

    \I__12689\ : ClkMux
    port map (
            O => \N__51113\,
            I => \N__50675\
        );

    \I__12688\ : ClkMux
    port map (
            O => \N__51112\,
            I => \N__50675\
        );

    \I__12687\ : ClkMux
    port map (
            O => \N__51111\,
            I => \N__50675\
        );

    \I__12686\ : ClkMux
    port map (
            O => \N__51110\,
            I => \N__50675\
        );

    \I__12685\ : ClkMux
    port map (
            O => \N__51109\,
            I => \N__50675\
        );

    \I__12684\ : ClkMux
    port map (
            O => \N__51108\,
            I => \N__50675\
        );

    \I__12683\ : ClkMux
    port map (
            O => \N__51107\,
            I => \N__50675\
        );

    \I__12682\ : ClkMux
    port map (
            O => \N__51106\,
            I => \N__50675\
        );

    \I__12681\ : GlobalMux
    port map (
            O => \N__50675\,
            I => \clk_32MHz\
        );

    \I__12680\ : SRMux
    port map (
            O => \N__50672\,
            I => \N__50669\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__50669\,
            I => \N__50666\
        );

    \I__12678\ : Span4Mux_h
    port map (
            O => \N__50666\,
            I => \N__50663\
        );

    \I__12677\ : Odrv4
    port map (
            O => \N__50663\,
            I => \comm_spi.iclk_N_801\
        );

    \I__12676\ : CEMux
    port map (
            O => \N__50660\,
            I => \N__50657\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__50657\,
            I => \N__50653\
        );

    \I__12674\ : CEMux
    port map (
            O => \N__50656\,
            I => \N__50650\
        );

    \I__12673\ : Span4Mux_v
    port map (
            O => \N__50653\,
            I => \N__50647\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__50650\,
            I => \N__50644\
        );

    \I__12671\ : Span4Mux_h
    port map (
            O => \N__50647\,
            I => \N__50641\
        );

    \I__12670\ : Span4Mux_h
    port map (
            O => \N__50644\,
            I => \N__50638\
        );

    \I__12669\ : Odrv4
    port map (
            O => \N__50641\,
            I => n8576
        );

    \I__12668\ : Odrv4
    port map (
            O => \N__50638\,
            I => n8576
        );

    \I__12667\ : CEMux
    port map (
            O => \N__50633\,
            I => \N__50630\
        );

    \I__12666\ : LocalMux
    port map (
            O => \N__50630\,
            I => \N__50627\
        );

    \I__12665\ : Span4Mux_h
    port map (
            O => \N__50627\,
            I => \N__50624\
        );

    \I__12664\ : Odrv4
    port map (
            O => \N__50624\,
            I => n8117
        );

    \I__12663\ : InMux
    port map (
            O => \N__50621\,
            I => \N__50618\
        );

    \I__12662\ : LocalMux
    port map (
            O => \N__50618\,
            I => \N__50615\
        );

    \I__12661\ : Span4Mux_h
    port map (
            O => \N__50615\,
            I => \N__50612\
        );

    \I__12660\ : Odrv4
    port map (
            O => \N__50612\,
            I => n6_adj_1175
        );

    \I__12659\ : InMux
    port map (
            O => \N__50609\,
            I => \N__50606\
        );

    \I__12658\ : LocalMux
    port map (
            O => \N__50606\,
            I => \N__50590\
        );

    \I__12657\ : InMux
    port map (
            O => \N__50605\,
            I => \N__50583\
        );

    \I__12656\ : InMux
    port map (
            O => \N__50604\,
            I => \N__50583\
        );

    \I__12655\ : InMux
    port map (
            O => \N__50603\,
            I => \N__50583\
        );

    \I__12654\ : InMux
    port map (
            O => \N__50602\,
            I => \N__50575\
        );

    \I__12653\ : InMux
    port map (
            O => \N__50601\,
            I => \N__50575\
        );

    \I__12652\ : InMux
    port map (
            O => \N__50600\,
            I => \N__50570\
        );

    \I__12651\ : InMux
    port map (
            O => \N__50599\,
            I => \N__50570\
        );

    \I__12650\ : InMux
    port map (
            O => \N__50598\,
            I => \N__50565\
        );

    \I__12649\ : InMux
    port map (
            O => \N__50597\,
            I => \N__50565\
        );

    \I__12648\ : InMux
    port map (
            O => \N__50596\,
            I => \N__50562\
        );

    \I__12647\ : InMux
    port map (
            O => \N__50595\,
            I => \N__50555\
        );

    \I__12646\ : InMux
    port map (
            O => \N__50594\,
            I => \N__50547\
        );

    \I__12645\ : InMux
    port map (
            O => \N__50593\,
            I => \N__50544\
        );

    \I__12644\ : Span4Mux_v
    port map (
            O => \N__50590\,
            I => \N__50541\
        );

    \I__12643\ : LocalMux
    port map (
            O => \N__50583\,
            I => \N__50538\
        );

    \I__12642\ : InMux
    port map (
            O => \N__50582\,
            I => \N__50533\
        );

    \I__12641\ : InMux
    port map (
            O => \N__50581\,
            I => \N__50528\
        );

    \I__12640\ : InMux
    port map (
            O => \N__50580\,
            I => \N__50528\
        );

    \I__12639\ : LocalMux
    port map (
            O => \N__50575\,
            I => \N__50525\
        );

    \I__12638\ : LocalMux
    port map (
            O => \N__50570\,
            I => \N__50520\
        );

    \I__12637\ : LocalMux
    port map (
            O => \N__50565\,
            I => \N__50520\
        );

    \I__12636\ : LocalMux
    port map (
            O => \N__50562\,
            I => \N__50517\
        );

    \I__12635\ : InMux
    port map (
            O => \N__50561\,
            I => \N__50514\
        );

    \I__12634\ : InMux
    port map (
            O => \N__50560\,
            I => \N__50493\
        );

    \I__12633\ : InMux
    port map (
            O => \N__50559\,
            I => \N__50493\
        );

    \I__12632\ : InMux
    port map (
            O => \N__50558\,
            I => \N__50490\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__50555\,
            I => \N__50487\
        );

    \I__12630\ : InMux
    port map (
            O => \N__50554\,
            I => \N__50478\
        );

    \I__12629\ : InMux
    port map (
            O => \N__50553\,
            I => \N__50478\
        );

    \I__12628\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50478\
        );

    \I__12627\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50478\
        );

    \I__12626\ : CascadeMux
    port map (
            O => \N__50550\,
            I => \N__50473\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__50547\,
            I => \N__50468\
        );

    \I__12624\ : LocalMux
    port map (
            O => \N__50544\,
            I => \N__50468\
        );

    \I__12623\ : Span4Mux_h
    port map (
            O => \N__50541\,
            I => \N__50465\
        );

    \I__12622\ : Span12Mux_v
    port map (
            O => \N__50538\,
            I => \N__50462\
        );

    \I__12621\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50459\
        );

    \I__12620\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50456\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__50533\,
            I => \N__50447\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__50528\,
            I => \N__50447\
        );

    \I__12617\ : Span4Mux_v
    port map (
            O => \N__50525\,
            I => \N__50447\
        );

    \I__12616\ : Span4Mux_v
    port map (
            O => \N__50520\,
            I => \N__50447\
        );

    \I__12615\ : Span4Mux_h
    port map (
            O => \N__50517\,
            I => \N__50442\
        );

    \I__12614\ : LocalMux
    port map (
            O => \N__50514\,
            I => \N__50442\
        );

    \I__12613\ : InMux
    port map (
            O => \N__50513\,
            I => \N__50439\
        );

    \I__12612\ : InMux
    port map (
            O => \N__50512\,
            I => \N__50428\
        );

    \I__12611\ : InMux
    port map (
            O => \N__50511\,
            I => \N__50428\
        );

    \I__12610\ : InMux
    port map (
            O => \N__50510\,
            I => \N__50428\
        );

    \I__12609\ : InMux
    port map (
            O => \N__50509\,
            I => \N__50428\
        );

    \I__12608\ : InMux
    port map (
            O => \N__50508\,
            I => \N__50428\
        );

    \I__12607\ : InMux
    port map (
            O => \N__50507\,
            I => \N__50421\
        );

    \I__12606\ : InMux
    port map (
            O => \N__50506\,
            I => \N__50421\
        );

    \I__12605\ : InMux
    port map (
            O => \N__50505\,
            I => \N__50421\
        );

    \I__12604\ : InMux
    port map (
            O => \N__50504\,
            I => \N__50416\
        );

    \I__12603\ : InMux
    port map (
            O => \N__50503\,
            I => \N__50416\
        );

    \I__12602\ : InMux
    port map (
            O => \N__50502\,
            I => \N__50413\
        );

    \I__12601\ : InMux
    port map (
            O => \N__50501\,
            I => \N__50408\
        );

    \I__12600\ : InMux
    port map (
            O => \N__50500\,
            I => \N__50408\
        );

    \I__12599\ : InMux
    port map (
            O => \N__50499\,
            I => \N__50403\
        );

    \I__12598\ : InMux
    port map (
            O => \N__50498\,
            I => \N__50403\
        );

    \I__12597\ : LocalMux
    port map (
            O => \N__50493\,
            I => \N__50394\
        );

    \I__12596\ : LocalMux
    port map (
            O => \N__50490\,
            I => \N__50394\
        );

    \I__12595\ : Span4Mux_v
    port map (
            O => \N__50487\,
            I => \N__50394\
        );

    \I__12594\ : LocalMux
    port map (
            O => \N__50478\,
            I => \N__50394\
        );

    \I__12593\ : InMux
    port map (
            O => \N__50477\,
            I => \N__50387\
        );

    \I__12592\ : InMux
    port map (
            O => \N__50476\,
            I => \N__50387\
        );

    \I__12591\ : InMux
    port map (
            O => \N__50473\,
            I => \N__50387\
        );

    \I__12590\ : Span4Mux_v
    port map (
            O => \N__50468\,
            I => \N__50384\
        );

    \I__12589\ : Sp12to4
    port map (
            O => \N__50465\,
            I => \N__50377\
        );

    \I__12588\ : Span12Mux_h
    port map (
            O => \N__50462\,
            I => \N__50377\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__50459\,
            I => \N__50377\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__50456\,
            I => \N__50370\
        );

    \I__12585\ : Span4Mux_h
    port map (
            O => \N__50447\,
            I => \N__50370\
        );

    \I__12584\ : Span4Mux_v
    port map (
            O => \N__50442\,
            I => \N__50370\
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__50439\,
            I => comm_state_0
        );

    \I__12582\ : LocalMux
    port map (
            O => \N__50428\,
            I => comm_state_0
        );

    \I__12581\ : LocalMux
    port map (
            O => \N__50421\,
            I => comm_state_0
        );

    \I__12580\ : LocalMux
    port map (
            O => \N__50416\,
            I => comm_state_0
        );

    \I__12579\ : LocalMux
    port map (
            O => \N__50413\,
            I => comm_state_0
        );

    \I__12578\ : LocalMux
    port map (
            O => \N__50408\,
            I => comm_state_0
        );

    \I__12577\ : LocalMux
    port map (
            O => \N__50403\,
            I => comm_state_0
        );

    \I__12576\ : Odrv4
    port map (
            O => \N__50394\,
            I => comm_state_0
        );

    \I__12575\ : LocalMux
    port map (
            O => \N__50387\,
            I => comm_state_0
        );

    \I__12574\ : Odrv4
    port map (
            O => \N__50384\,
            I => comm_state_0
        );

    \I__12573\ : Odrv12
    port map (
            O => \N__50377\,
            I => comm_state_0
        );

    \I__12572\ : Odrv4
    port map (
            O => \N__50370\,
            I => comm_state_0
        );

    \I__12571\ : InMux
    port map (
            O => \N__50345\,
            I => \N__50334\
        );

    \I__12570\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50331\
        );

    \I__12569\ : InMux
    port map (
            O => \N__50343\,
            I => \N__50297\
        );

    \I__12568\ : InMux
    port map (
            O => \N__50342\,
            I => \N__50294\
        );

    \I__12567\ : InMux
    port map (
            O => \N__50341\,
            I => \N__50247\
        );

    \I__12566\ : InMux
    port map (
            O => \N__50340\,
            I => \N__50247\
        );

    \I__12565\ : InMux
    port map (
            O => \N__50339\,
            I => \N__50240\
        );

    \I__12564\ : InMux
    port map (
            O => \N__50338\,
            I => \N__50240\
        );

    \I__12563\ : InMux
    port map (
            O => \N__50337\,
            I => \N__50240\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__50334\,
            I => \N__50235\
        );

    \I__12561\ : LocalMux
    port map (
            O => \N__50331\,
            I => \N__50235\
        );

    \I__12560\ : InMux
    port map (
            O => \N__50330\,
            I => \N__50230\
        );

    \I__12559\ : InMux
    port map (
            O => \N__50329\,
            I => \N__50230\
        );

    \I__12558\ : InMux
    port map (
            O => \N__50328\,
            I => \N__50221\
        );

    \I__12557\ : InMux
    port map (
            O => \N__50327\,
            I => \N__50221\
        );

    \I__12556\ : InMux
    port map (
            O => \N__50326\,
            I => \N__50221\
        );

    \I__12555\ : InMux
    port map (
            O => \N__50325\,
            I => \N__50221\
        );

    \I__12554\ : CascadeMux
    port map (
            O => \N__50324\,
            I => \N__50216\
        );

    \I__12553\ : InMux
    port map (
            O => \N__50323\,
            I => \N__50212\
        );

    \I__12552\ : CascadeMux
    port map (
            O => \N__50322\,
            I => \N__50207\
        );

    \I__12551\ : InMux
    port map (
            O => \N__50321\,
            I => \N__50204\
        );

    \I__12550\ : InMux
    port map (
            O => \N__50320\,
            I => \N__50183\
        );

    \I__12549\ : InMux
    port map (
            O => \N__50319\,
            I => \N__50183\
        );

    \I__12548\ : InMux
    port map (
            O => \N__50318\,
            I => \N__50183\
        );

    \I__12547\ : InMux
    port map (
            O => \N__50317\,
            I => \N__50183\
        );

    \I__12546\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50183\
        );

    \I__12545\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50183\
        );

    \I__12544\ : InMux
    port map (
            O => \N__50314\,
            I => \N__50183\
        );

    \I__12543\ : InMux
    port map (
            O => \N__50313\,
            I => \N__50183\
        );

    \I__12542\ : InMux
    port map (
            O => \N__50312\,
            I => \N__50178\
        );

    \I__12541\ : InMux
    port map (
            O => \N__50311\,
            I => \N__50178\
        );

    \I__12540\ : InMux
    port map (
            O => \N__50310\,
            I => \N__50167\
        );

    \I__12539\ : InMux
    port map (
            O => \N__50309\,
            I => \N__50167\
        );

    \I__12538\ : InMux
    port map (
            O => \N__50308\,
            I => \N__50167\
        );

    \I__12537\ : InMux
    port map (
            O => \N__50307\,
            I => \N__50167\
        );

    \I__12536\ : InMux
    port map (
            O => \N__50306\,
            I => \N__50167\
        );

    \I__12535\ : InMux
    port map (
            O => \N__50305\,
            I => \N__50164\
        );

    \I__12534\ : InMux
    port map (
            O => \N__50304\,
            I => \N__50153\
        );

    \I__12533\ : InMux
    port map (
            O => \N__50303\,
            I => \N__50153\
        );

    \I__12532\ : InMux
    port map (
            O => \N__50302\,
            I => \N__50153\
        );

    \I__12531\ : InMux
    port map (
            O => \N__50301\,
            I => \N__50153\
        );

    \I__12530\ : InMux
    port map (
            O => \N__50300\,
            I => \N__50153\
        );

    \I__12529\ : LocalMux
    port map (
            O => \N__50297\,
            I => \N__50144\
        );

    \I__12528\ : LocalMux
    port map (
            O => \N__50294\,
            I => \N__50144\
        );

    \I__12527\ : CascadeMux
    port map (
            O => \N__50293\,
            I => \N__50138\
        );

    \I__12526\ : CascadeMux
    port map (
            O => \N__50292\,
            I => \N__50135\
        );

    \I__12525\ : InMux
    port map (
            O => \N__50291\,
            I => \N__50132\
        );

    \I__12524\ : CascadeMux
    port map (
            O => \N__50290\,
            I => \N__50128\
        );

    \I__12523\ : InMux
    port map (
            O => \N__50289\,
            I => \N__50124\
        );

    \I__12522\ : InMux
    port map (
            O => \N__50288\,
            I => \N__50115\
        );

    \I__12521\ : InMux
    port map (
            O => \N__50287\,
            I => \N__50115\
        );

    \I__12520\ : InMux
    port map (
            O => \N__50286\,
            I => \N__50099\
        );

    \I__12519\ : InMux
    port map (
            O => \N__50285\,
            I => \N__50099\
        );

    \I__12518\ : InMux
    port map (
            O => \N__50284\,
            I => \N__50099\
        );

    \I__12517\ : InMux
    port map (
            O => \N__50283\,
            I => \N__50094\
        );

    \I__12516\ : InMux
    port map (
            O => \N__50282\,
            I => \N__50094\
        );

    \I__12515\ : InMux
    port map (
            O => \N__50281\,
            I => \N__50085\
        );

    \I__12514\ : InMux
    port map (
            O => \N__50280\,
            I => \N__50078\
        );

    \I__12513\ : InMux
    port map (
            O => \N__50279\,
            I => \N__50078\
        );

    \I__12512\ : InMux
    port map (
            O => \N__50278\,
            I => \N__50078\
        );

    \I__12511\ : InMux
    port map (
            O => \N__50277\,
            I => \N__50069\
        );

    \I__12510\ : InMux
    port map (
            O => \N__50276\,
            I => \N__50069\
        );

    \I__12509\ : InMux
    port map (
            O => \N__50275\,
            I => \N__50069\
        );

    \I__12508\ : InMux
    port map (
            O => \N__50274\,
            I => \N__50069\
        );

    \I__12507\ : InMux
    port map (
            O => \N__50273\,
            I => \N__50060\
        );

    \I__12506\ : InMux
    port map (
            O => \N__50272\,
            I => \N__50060\
        );

    \I__12505\ : InMux
    port map (
            O => \N__50271\,
            I => \N__50060\
        );

    \I__12504\ : InMux
    port map (
            O => \N__50270\,
            I => \N__50060\
        );

    \I__12503\ : InMux
    port map (
            O => \N__50269\,
            I => \N__50057\
        );

    \I__12502\ : InMux
    port map (
            O => \N__50268\,
            I => \N__50054\
        );

    \I__12501\ : InMux
    port map (
            O => \N__50267\,
            I => \N__50051\
        );

    \I__12500\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50048\
        );

    \I__12499\ : InMux
    port map (
            O => \N__50265\,
            I => \N__50031\
        );

    \I__12498\ : InMux
    port map (
            O => \N__50264\,
            I => \N__50031\
        );

    \I__12497\ : InMux
    port map (
            O => \N__50263\,
            I => \N__50031\
        );

    \I__12496\ : InMux
    port map (
            O => \N__50262\,
            I => \N__50031\
        );

    \I__12495\ : InMux
    port map (
            O => \N__50261\,
            I => \N__50031\
        );

    \I__12494\ : InMux
    port map (
            O => \N__50260\,
            I => \N__50031\
        );

    \I__12493\ : InMux
    port map (
            O => \N__50259\,
            I => \N__50031\
        );

    \I__12492\ : InMux
    port map (
            O => \N__50258\,
            I => \N__50031\
        );

    \I__12491\ : InMux
    port map (
            O => \N__50257\,
            I => \N__50018\
        );

    \I__12490\ : InMux
    port map (
            O => \N__50256\,
            I => \N__50018\
        );

    \I__12489\ : InMux
    port map (
            O => \N__50255\,
            I => \N__50018\
        );

    \I__12488\ : InMux
    port map (
            O => \N__50254\,
            I => \N__50018\
        );

    \I__12487\ : InMux
    port map (
            O => \N__50253\,
            I => \N__50018\
        );

    \I__12486\ : InMux
    port map (
            O => \N__50252\,
            I => \N__50018\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__50247\,
            I => \N__50015\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__50240\,
            I => \N__50012\
        );

    \I__12483\ : Span4Mux_h
    port map (
            O => \N__50235\,
            I => \N__50005\
        );

    \I__12482\ : LocalMux
    port map (
            O => \N__50230\,
            I => \N__50005\
        );

    \I__12481\ : LocalMux
    port map (
            O => \N__50221\,
            I => \N__50005\
        );

    \I__12480\ : CascadeMux
    port map (
            O => \N__50220\,
            I => \N__50001\
        );

    \I__12479\ : CascadeMux
    port map (
            O => \N__50219\,
            I => \N__49997\
        );

    \I__12478\ : InMux
    port map (
            O => \N__50216\,
            I => \N__49993\
        );

    \I__12477\ : InMux
    port map (
            O => \N__50215\,
            I => \N__49990\
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__50212\,
            I => \N__49987\
        );

    \I__12475\ : InMux
    port map (
            O => \N__50211\,
            I => \N__49980\
        );

    \I__12474\ : InMux
    port map (
            O => \N__50210\,
            I => \N__49980\
        );

    \I__12473\ : InMux
    port map (
            O => \N__50207\,
            I => \N__49980\
        );

    \I__12472\ : LocalMux
    port map (
            O => \N__50204\,
            I => \N__49977\
        );

    \I__12471\ : InMux
    port map (
            O => \N__50203\,
            I => \N__49972\
        );

    \I__12470\ : InMux
    port map (
            O => \N__50202\,
            I => \N__49972\
        );

    \I__12469\ : InMux
    port map (
            O => \N__50201\,
            I => \N__49967\
        );

    \I__12468\ : InMux
    port map (
            O => \N__50200\,
            I => \N__49967\
        );

    \I__12467\ : LocalMux
    port map (
            O => \N__50183\,
            I => \N__49962\
        );

    \I__12466\ : LocalMux
    port map (
            O => \N__50178\,
            I => \N__49957\
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__50167\,
            I => \N__49957\
        );

    \I__12464\ : LocalMux
    port map (
            O => \N__50164\,
            I => \N__49952\
        );

    \I__12463\ : LocalMux
    port map (
            O => \N__50153\,
            I => \N__49952\
        );

    \I__12462\ : InMux
    port map (
            O => \N__50152\,
            I => \N__49943\
        );

    \I__12461\ : InMux
    port map (
            O => \N__50151\,
            I => \N__49943\
        );

    \I__12460\ : InMux
    port map (
            O => \N__50150\,
            I => \N__49943\
        );

    \I__12459\ : InMux
    port map (
            O => \N__50149\,
            I => \N__49943\
        );

    \I__12458\ : Span4Mux_h
    port map (
            O => \N__50144\,
            I => \N__49940\
        );

    \I__12457\ : CascadeMux
    port map (
            O => \N__50143\,
            I => \N__49935\
        );

    \I__12456\ : InMux
    port map (
            O => \N__50142\,
            I => \N__49932\
        );

    \I__12455\ : InMux
    port map (
            O => \N__50141\,
            I => \N__49929\
        );

    \I__12454\ : InMux
    port map (
            O => \N__50138\,
            I => \N__49924\
        );

    \I__12453\ : InMux
    port map (
            O => \N__50135\,
            I => \N__49924\
        );

    \I__12452\ : LocalMux
    port map (
            O => \N__50132\,
            I => \N__49921\
        );

    \I__12451\ : InMux
    port map (
            O => \N__50131\,
            I => \N__49914\
        );

    \I__12450\ : InMux
    port map (
            O => \N__50128\,
            I => \N__49914\
        );

    \I__12449\ : InMux
    port map (
            O => \N__50127\,
            I => \N__49914\
        );

    \I__12448\ : LocalMux
    port map (
            O => \N__50124\,
            I => \N__49911\
        );

    \I__12447\ : InMux
    port map (
            O => \N__50123\,
            I => \N__49902\
        );

    \I__12446\ : InMux
    port map (
            O => \N__50122\,
            I => \N__49902\
        );

    \I__12445\ : InMux
    port map (
            O => \N__50121\,
            I => \N__49902\
        );

    \I__12444\ : InMux
    port map (
            O => \N__50120\,
            I => \N__49902\
        );

    \I__12443\ : LocalMux
    port map (
            O => \N__50115\,
            I => \N__49899\
        );

    \I__12442\ : InMux
    port map (
            O => \N__50114\,
            I => \N__49882\
        );

    \I__12441\ : InMux
    port map (
            O => \N__50113\,
            I => \N__49882\
        );

    \I__12440\ : InMux
    port map (
            O => \N__50112\,
            I => \N__49882\
        );

    \I__12439\ : CascadeMux
    port map (
            O => \N__50111\,
            I => \N__49876\
        );

    \I__12438\ : InMux
    port map (
            O => \N__50110\,
            I => \N__49871\
        );

    \I__12437\ : InMux
    port map (
            O => \N__50109\,
            I => \N__49865\
        );

    \I__12436\ : InMux
    port map (
            O => \N__50108\,
            I => \N__49862\
        );

    \I__12435\ : InMux
    port map (
            O => \N__50107\,
            I => \N__49859\
        );

    \I__12434\ : InMux
    port map (
            O => \N__50106\,
            I => \N__49856\
        );

    \I__12433\ : LocalMux
    port map (
            O => \N__50099\,
            I => \N__49851\
        );

    \I__12432\ : LocalMux
    port map (
            O => \N__50094\,
            I => \N__49851\
        );

    \I__12431\ : InMux
    port map (
            O => \N__50093\,
            I => \N__49848\
        );

    \I__12430\ : InMux
    port map (
            O => \N__50092\,
            I => \N__49845\
        );

    \I__12429\ : InMux
    port map (
            O => \N__50091\,
            I => \N__49836\
        );

    \I__12428\ : InMux
    port map (
            O => \N__50090\,
            I => \N__49836\
        );

    \I__12427\ : InMux
    port map (
            O => \N__50089\,
            I => \N__49836\
        );

    \I__12426\ : InMux
    port map (
            O => \N__50088\,
            I => \N__49836\
        );

    \I__12425\ : LocalMux
    port map (
            O => \N__50085\,
            I => \N__49831\
        );

    \I__12424\ : LocalMux
    port map (
            O => \N__50078\,
            I => \N__49831\
        );

    \I__12423\ : LocalMux
    port map (
            O => \N__50069\,
            I => \N__49820\
        );

    \I__12422\ : LocalMux
    port map (
            O => \N__50060\,
            I => \N__49820\
        );

    \I__12421\ : LocalMux
    port map (
            O => \N__50057\,
            I => \N__49820\
        );

    \I__12420\ : LocalMux
    port map (
            O => \N__50054\,
            I => \N__49820\
        );

    \I__12419\ : LocalMux
    port map (
            O => \N__50051\,
            I => \N__49820\
        );

    \I__12418\ : LocalMux
    port map (
            O => \N__50048\,
            I => \N__49806\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__50031\,
            I => \N__49806\
        );

    \I__12416\ : LocalMux
    port map (
            O => \N__50018\,
            I => \N__49806\
        );

    \I__12415\ : Span4Mux_h
    port map (
            O => \N__50015\,
            I => \N__49806\
        );

    \I__12414\ : Span4Mux_h
    port map (
            O => \N__50012\,
            I => \N__49806\
        );

    \I__12413\ : Span4Mux_v
    port map (
            O => \N__50005\,
            I => \N__49806\
        );

    \I__12412\ : InMux
    port map (
            O => \N__50004\,
            I => \N__49795\
        );

    \I__12411\ : InMux
    port map (
            O => \N__50001\,
            I => \N__49795\
        );

    \I__12410\ : InMux
    port map (
            O => \N__50000\,
            I => \N__49795\
        );

    \I__12409\ : InMux
    port map (
            O => \N__49997\,
            I => \N__49795\
        );

    \I__12408\ : InMux
    port map (
            O => \N__49996\,
            I => \N__49795\
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__49993\,
            I => \N__49792\
        );

    \I__12406\ : LocalMux
    port map (
            O => \N__49990\,
            I => \N__49779\
        );

    \I__12405\ : Span4Mux_h
    port map (
            O => \N__49987\,
            I => \N__49779\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__49980\,
            I => \N__49779\
        );

    \I__12403\ : Span4Mux_h
    port map (
            O => \N__49977\,
            I => \N__49779\
        );

    \I__12402\ : LocalMux
    port map (
            O => \N__49972\,
            I => \N__49779\
        );

    \I__12401\ : LocalMux
    port map (
            O => \N__49967\,
            I => \N__49779\
        );

    \I__12400\ : InMux
    port map (
            O => \N__49966\,
            I => \N__49776\
        );

    \I__12399\ : InMux
    port map (
            O => \N__49965\,
            I => \N__49770\
        );

    \I__12398\ : Span4Mux_v
    port map (
            O => \N__49962\,
            I => \N__49763\
        );

    \I__12397\ : Span4Mux_v
    port map (
            O => \N__49957\,
            I => \N__49763\
        );

    \I__12396\ : Span4Mux_v
    port map (
            O => \N__49952\,
            I => \N__49763\
        );

    \I__12395\ : LocalMux
    port map (
            O => \N__49943\,
            I => \N__49758\
        );

    \I__12394\ : Span4Mux_h
    port map (
            O => \N__49940\,
            I => \N__49758\
        );

    \I__12393\ : InMux
    port map (
            O => \N__49939\,
            I => \N__49753\
        );

    \I__12392\ : InMux
    port map (
            O => \N__49938\,
            I => \N__49753\
        );

    \I__12391\ : InMux
    port map (
            O => \N__49935\,
            I => \N__49750\
        );

    \I__12390\ : LocalMux
    port map (
            O => \N__49932\,
            I => \N__49747\
        );

    \I__12389\ : LocalMux
    port map (
            O => \N__49929\,
            I => \N__49742\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__49924\,
            I => \N__49742\
        );

    \I__12387\ : Span4Mux_h
    port map (
            O => \N__49921\,
            I => \N__49736\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__49914\,
            I => \N__49736\
        );

    \I__12385\ : Span4Mux_v
    port map (
            O => \N__49911\,
            I => \N__49726\
        );

    \I__12384\ : LocalMux
    port map (
            O => \N__49902\,
            I => \N__49726\
        );

    \I__12383\ : Span4Mux_h
    port map (
            O => \N__49899\,
            I => \N__49726\
        );

    \I__12382\ : InMux
    port map (
            O => \N__49898\,
            I => \N__49721\
        );

    \I__12381\ : InMux
    port map (
            O => \N__49897\,
            I => \N__49721\
        );

    \I__12380\ : InMux
    port map (
            O => \N__49896\,
            I => \N__49716\
        );

    \I__12379\ : InMux
    port map (
            O => \N__49895\,
            I => \N__49716\
        );

    \I__12378\ : InMux
    port map (
            O => \N__49894\,
            I => \N__49703\
        );

    \I__12377\ : InMux
    port map (
            O => \N__49893\,
            I => \N__49703\
        );

    \I__12376\ : InMux
    port map (
            O => \N__49892\,
            I => \N__49703\
        );

    \I__12375\ : InMux
    port map (
            O => \N__49891\,
            I => \N__49703\
        );

    \I__12374\ : InMux
    port map (
            O => \N__49890\,
            I => \N__49703\
        );

    \I__12373\ : InMux
    port map (
            O => \N__49889\,
            I => \N__49703\
        );

    \I__12372\ : LocalMux
    port map (
            O => \N__49882\,
            I => \N__49700\
        );

    \I__12371\ : InMux
    port map (
            O => \N__49881\,
            I => \N__49695\
        );

    \I__12370\ : InMux
    port map (
            O => \N__49880\,
            I => \N__49695\
        );

    \I__12369\ : InMux
    port map (
            O => \N__49879\,
            I => \N__49688\
        );

    \I__12368\ : InMux
    port map (
            O => \N__49876\,
            I => \N__49688\
        );

    \I__12367\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49688\
        );

    \I__12366\ : InMux
    port map (
            O => \N__49874\,
            I => \N__49685\
        );

    \I__12365\ : LocalMux
    port map (
            O => \N__49871\,
            I => \N__49682\
        );

    \I__12364\ : InMux
    port map (
            O => \N__49870\,
            I => \N__49675\
        );

    \I__12363\ : InMux
    port map (
            O => \N__49869\,
            I => \N__49675\
        );

    \I__12362\ : InMux
    port map (
            O => \N__49868\,
            I => \N__49675\
        );

    \I__12361\ : LocalMux
    port map (
            O => \N__49865\,
            I => \N__49660\
        );

    \I__12360\ : LocalMux
    port map (
            O => \N__49862\,
            I => \N__49660\
        );

    \I__12359\ : LocalMux
    port map (
            O => \N__49859\,
            I => \N__49660\
        );

    \I__12358\ : LocalMux
    port map (
            O => \N__49856\,
            I => \N__49660\
        );

    \I__12357\ : Sp12to4
    port map (
            O => \N__49851\,
            I => \N__49660\
        );

    \I__12356\ : LocalMux
    port map (
            O => \N__49848\,
            I => \N__49660\
        );

    \I__12355\ : LocalMux
    port map (
            O => \N__49845\,
            I => \N__49660\
        );

    \I__12354\ : LocalMux
    port map (
            O => \N__49836\,
            I => \N__49653\
        );

    \I__12353\ : Span4Mux_v
    port map (
            O => \N__49831\,
            I => \N__49653\
        );

    \I__12352\ : Span4Mux_v
    port map (
            O => \N__49820\,
            I => \N__49653\
        );

    \I__12351\ : InMux
    port map (
            O => \N__49819\,
            I => \N__49650\
        );

    \I__12350\ : Span4Mux_h
    port map (
            O => \N__49806\,
            I => \N__49645\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__49795\,
            I => \N__49645\
        );

    \I__12348\ : Span4Mux_h
    port map (
            O => \N__49792\,
            I => \N__49638\
        );

    \I__12347\ : Span4Mux_v
    port map (
            O => \N__49779\,
            I => \N__49638\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__49776\,
            I => \N__49638\
        );

    \I__12345\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49631\
        );

    \I__12344\ : InMux
    port map (
            O => \N__49774\,
            I => \N__49631\
        );

    \I__12343\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49631\
        );

    \I__12342\ : LocalMux
    port map (
            O => \N__49770\,
            I => \N__49628\
        );

    \I__12341\ : Span4Mux_h
    port map (
            O => \N__49763\,
            I => \N__49615\
        );

    \I__12340\ : Span4Mux_v
    port map (
            O => \N__49758\,
            I => \N__49615\
        );

    \I__12339\ : LocalMux
    port map (
            O => \N__49753\,
            I => \N__49615\
        );

    \I__12338\ : LocalMux
    port map (
            O => \N__49750\,
            I => \N__49615\
        );

    \I__12337\ : Span4Mux_v
    port map (
            O => \N__49747\,
            I => \N__49615\
        );

    \I__12336\ : Span4Mux_h
    port map (
            O => \N__49742\,
            I => \N__49615\
        );

    \I__12335\ : InMux
    port map (
            O => \N__49741\,
            I => \N__49612\
        );

    \I__12334\ : Span4Mux_h
    port map (
            O => \N__49736\,
            I => \N__49609\
        );

    \I__12333\ : InMux
    port map (
            O => \N__49735\,
            I => \N__49602\
        );

    \I__12332\ : InMux
    port map (
            O => \N__49734\,
            I => \N__49602\
        );

    \I__12331\ : InMux
    port map (
            O => \N__49733\,
            I => \N__49602\
        );

    \I__12330\ : Span4Mux_v
    port map (
            O => \N__49726\,
            I => \N__49599\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__49721\,
            I => \N__49576\
        );

    \I__12328\ : LocalMux
    port map (
            O => \N__49716\,
            I => \N__49576\
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__49703\,
            I => \N__49576\
        );

    \I__12326\ : Span12Mux_v
    port map (
            O => \N__49700\,
            I => \N__49576\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__49695\,
            I => \N__49576\
        );

    \I__12324\ : LocalMux
    port map (
            O => \N__49688\,
            I => \N__49576\
        );

    \I__12323\ : LocalMux
    port map (
            O => \N__49685\,
            I => \N__49576\
        );

    \I__12322\ : Span12Mux_v
    port map (
            O => \N__49682\,
            I => \N__49576\
        );

    \I__12321\ : LocalMux
    port map (
            O => \N__49675\,
            I => \N__49576\
        );

    \I__12320\ : Span12Mux_v
    port map (
            O => \N__49660\,
            I => \N__49576\
        );

    \I__12319\ : Sp12to4
    port map (
            O => \N__49653\,
            I => \N__49576\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__49650\,
            I => \N__49569\
        );

    \I__12317\ : Span4Mux_h
    port map (
            O => \N__49645\,
            I => \N__49569\
        );

    \I__12316\ : Span4Mux_h
    port map (
            O => \N__49638\,
            I => \N__49569\
        );

    \I__12315\ : LocalMux
    port map (
            O => \N__49631\,
            I => comm_state_1
        );

    \I__12314\ : Odrv4
    port map (
            O => \N__49628\,
            I => comm_state_1
        );

    \I__12313\ : Odrv4
    port map (
            O => \N__49615\,
            I => comm_state_1
        );

    \I__12312\ : LocalMux
    port map (
            O => \N__49612\,
            I => comm_state_1
        );

    \I__12311\ : Odrv4
    port map (
            O => \N__49609\,
            I => comm_state_1
        );

    \I__12310\ : LocalMux
    port map (
            O => \N__49602\,
            I => comm_state_1
        );

    \I__12309\ : Odrv4
    port map (
            O => \N__49599\,
            I => comm_state_1
        );

    \I__12308\ : Odrv12
    port map (
            O => \N__49576\,
            I => comm_state_1
        );

    \I__12307\ : Odrv4
    port map (
            O => \N__49569\,
            I => comm_state_1
        );

    \I__12306\ : InMux
    port map (
            O => \N__49550\,
            I => \N__49532\
        );

    \I__12305\ : InMux
    port map (
            O => \N__49549\,
            I => \N__49528\
        );

    \I__12304\ : InMux
    port map (
            O => \N__49548\,
            I => \N__49521\
        );

    \I__12303\ : InMux
    port map (
            O => \N__49547\,
            I => \N__49521\
        );

    \I__12302\ : InMux
    port map (
            O => \N__49546\,
            I => \N__49521\
        );

    \I__12301\ : InMux
    port map (
            O => \N__49545\,
            I => \N__49514\
        );

    \I__12300\ : InMux
    port map (
            O => \N__49544\,
            I => \N__49514\
        );

    \I__12299\ : InMux
    port map (
            O => \N__49543\,
            I => \N__49514\
        );

    \I__12298\ : InMux
    port map (
            O => \N__49542\,
            I => \N__49509\
        );

    \I__12297\ : InMux
    port map (
            O => \N__49541\,
            I => \N__49509\
        );

    \I__12296\ : InMux
    port map (
            O => \N__49540\,
            I => \N__49499\
        );

    \I__12295\ : InMux
    port map (
            O => \N__49539\,
            I => \N__49499\
        );

    \I__12294\ : CascadeMux
    port map (
            O => \N__49538\,
            I => \N__49496\
        );

    \I__12293\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49493\
        );

    \I__12292\ : InMux
    port map (
            O => \N__49536\,
            I => \N__49488\
        );

    \I__12291\ : InMux
    port map (
            O => \N__49535\,
            I => \N__49488\
        );

    \I__12290\ : LocalMux
    port map (
            O => \N__49532\,
            I => \N__49485\
        );

    \I__12289\ : InMux
    port map (
            O => \N__49531\,
            I => \N__49482\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__49528\,
            I => \N__49474\
        );

    \I__12287\ : LocalMux
    port map (
            O => \N__49521\,
            I => \N__49474\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__49514\,
            I => \N__49464\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__49509\,
            I => \N__49464\
        );

    \I__12284\ : InMux
    port map (
            O => \N__49508\,
            I => \N__49453\
        );

    \I__12283\ : InMux
    port map (
            O => \N__49507\,
            I => \N__49453\
        );

    \I__12282\ : InMux
    port map (
            O => \N__49506\,
            I => \N__49453\
        );

    \I__12281\ : InMux
    port map (
            O => \N__49505\,
            I => \N__49453\
        );

    \I__12280\ : InMux
    port map (
            O => \N__49504\,
            I => \N__49453\
        );

    \I__12279\ : LocalMux
    port map (
            O => \N__49499\,
            I => \N__49450\
        );

    \I__12278\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49447\
        );

    \I__12277\ : LocalMux
    port map (
            O => \N__49493\,
            I => \N__49442\
        );

    \I__12276\ : LocalMux
    port map (
            O => \N__49488\,
            I => \N__49439\
        );

    \I__12275\ : Span4Mux_v
    port map (
            O => \N__49485\,
            I => \N__49427\
        );

    \I__12274\ : LocalMux
    port map (
            O => \N__49482\,
            I => \N__49427\
        );

    \I__12273\ : InMux
    port map (
            O => \N__49481\,
            I => \N__49422\
        );

    \I__12272\ : InMux
    port map (
            O => \N__49480\,
            I => \N__49422\
        );

    \I__12271\ : InMux
    port map (
            O => \N__49479\,
            I => \N__49419\
        );

    \I__12270\ : Span4Mux_v
    port map (
            O => \N__49474\,
            I => \N__49416\
        );

    \I__12269\ : InMux
    port map (
            O => \N__49473\,
            I => \N__49407\
        );

    \I__12268\ : InMux
    port map (
            O => \N__49472\,
            I => \N__49407\
        );

    \I__12267\ : InMux
    port map (
            O => \N__49471\,
            I => \N__49407\
        );

    \I__12266\ : InMux
    port map (
            O => \N__49470\,
            I => \N__49407\
        );

    \I__12265\ : InMux
    port map (
            O => \N__49469\,
            I => \N__49399\
        );

    \I__12264\ : Span4Mux_v
    port map (
            O => \N__49464\,
            I => \N__49394\
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__49453\,
            I => \N__49394\
        );

    \I__12262\ : Span4Mux_v
    port map (
            O => \N__49450\,
            I => \N__49389\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__49447\,
            I => \N__49389\
        );

    \I__12260\ : InMux
    port map (
            O => \N__49446\,
            I => \N__49386\
        );

    \I__12259\ : InMux
    port map (
            O => \N__49445\,
            I => \N__49383\
        );

    \I__12258\ : Span12Mux_v
    port map (
            O => \N__49442\,
            I => \N__49378\
        );

    \I__12257\ : Span12Mux_s10_h
    port map (
            O => \N__49439\,
            I => \N__49378\
        );

    \I__12256\ : InMux
    port map (
            O => \N__49438\,
            I => \N__49375\
        );

    \I__12255\ : InMux
    port map (
            O => \N__49437\,
            I => \N__49372\
        );

    \I__12254\ : InMux
    port map (
            O => \N__49436\,
            I => \N__49369\
        );

    \I__12253\ : InMux
    port map (
            O => \N__49435\,
            I => \N__49360\
        );

    \I__12252\ : InMux
    port map (
            O => \N__49434\,
            I => \N__49360\
        );

    \I__12251\ : InMux
    port map (
            O => \N__49433\,
            I => \N__49360\
        );

    \I__12250\ : InMux
    port map (
            O => \N__49432\,
            I => \N__49360\
        );

    \I__12249\ : Span4Mux_h
    port map (
            O => \N__49427\,
            I => \N__49357\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__49422\,
            I => \N__49348\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__49419\,
            I => \N__49348\
        );

    \I__12246\ : Sp12to4
    port map (
            O => \N__49416\,
            I => \N__49348\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__49407\,
            I => \N__49348\
        );

    \I__12244\ : InMux
    port map (
            O => \N__49406\,
            I => \N__49343\
        );

    \I__12243\ : InMux
    port map (
            O => \N__49405\,
            I => \N__49343\
        );

    \I__12242\ : InMux
    port map (
            O => \N__49404\,
            I => \N__49338\
        );

    \I__12241\ : InMux
    port map (
            O => \N__49403\,
            I => \N__49338\
        );

    \I__12240\ : InMux
    port map (
            O => \N__49402\,
            I => \N__49335\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__49399\,
            I => \N__49328\
        );

    \I__12238\ : Span4Mux_h
    port map (
            O => \N__49394\,
            I => \N__49328\
        );

    \I__12237\ : Span4Mux_h
    port map (
            O => \N__49389\,
            I => \N__49328\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__49386\,
            I => \N__49321\
        );

    \I__12235\ : LocalMux
    port map (
            O => \N__49383\,
            I => \N__49321\
        );

    \I__12234\ : Span12Mux_h
    port map (
            O => \N__49378\,
            I => \N__49321\
        );

    \I__12233\ : LocalMux
    port map (
            O => \N__49375\,
            I => comm_state_2
        );

    \I__12232\ : LocalMux
    port map (
            O => \N__49372\,
            I => comm_state_2
        );

    \I__12231\ : LocalMux
    port map (
            O => \N__49369\,
            I => comm_state_2
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__49360\,
            I => comm_state_2
        );

    \I__12229\ : Odrv4
    port map (
            O => \N__49357\,
            I => comm_state_2
        );

    \I__12228\ : Odrv12
    port map (
            O => \N__49348\,
            I => comm_state_2
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__49343\,
            I => comm_state_2
        );

    \I__12226\ : LocalMux
    port map (
            O => \N__49338\,
            I => comm_state_2
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__49335\,
            I => comm_state_2
        );

    \I__12224\ : Odrv4
    port map (
            O => \N__49328\,
            I => comm_state_2
        );

    \I__12223\ : Odrv12
    port map (
            O => \N__49321\,
            I => comm_state_2
        );

    \I__12222\ : CEMux
    port map (
            O => \N__49298\,
            I => \N__49295\
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__49295\,
            I => \N__49292\
        );

    \I__12220\ : Span4Mux_v
    port map (
            O => \N__49292\,
            I => \N__49289\
        );

    \I__12219\ : Odrv4
    port map (
            O => \N__49289\,
            I => n8129
        );

    \I__12218\ : CascadeMux
    port map (
            O => \N__49286\,
            I => \N__49282\
        );

    \I__12217\ : InMux
    port map (
            O => \N__49285\,
            I => \N__49278\
        );

    \I__12216\ : InMux
    port map (
            O => \N__49282\,
            I => \N__49273\
        );

    \I__12215\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49273\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__49278\,
            I => cmd_rdadctmp_19_adj_1093
        );

    \I__12213\ : LocalMux
    port map (
            O => \N__49273\,
            I => cmd_rdadctmp_19_adj_1093
        );

    \I__12212\ : InMux
    port map (
            O => \N__49268\,
            I => \N__49257\
        );

    \I__12211\ : InMux
    port map (
            O => \N__49267\,
            I => \N__49257\
        );

    \I__12210\ : CascadeMux
    port map (
            O => \N__49266\,
            I => \N__49253\
        );

    \I__12209\ : InMux
    port map (
            O => \N__49265\,
            I => \N__49244\
        );

    \I__12208\ : InMux
    port map (
            O => \N__49264\,
            I => \N__49244\
        );

    \I__12207\ : InMux
    port map (
            O => \N__49263\,
            I => \N__49244\
        );

    \I__12206\ : InMux
    port map (
            O => \N__49262\,
            I => \N__49244\
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__49257\,
            I => \N__49234\
        );

    \I__12204\ : CascadeMux
    port map (
            O => \N__49256\,
            I => \N__49228\
        );

    \I__12203\ : InMux
    port map (
            O => \N__49253\,
            I => \N__49222\
        );

    \I__12202\ : LocalMux
    port map (
            O => \N__49244\,
            I => \N__49217\
        );

    \I__12201\ : InMux
    port map (
            O => \N__49243\,
            I => \N__49214\
        );

    \I__12200\ : InMux
    port map (
            O => \N__49242\,
            I => \N__49209\
        );

    \I__12199\ : CascadeMux
    port map (
            O => \N__49241\,
            I => \N__49206\
        );

    \I__12198\ : InMux
    port map (
            O => \N__49240\,
            I => \N__49186\
        );

    \I__12197\ : InMux
    port map (
            O => \N__49239\,
            I => \N__49183\
        );

    \I__12196\ : InMux
    port map (
            O => \N__49238\,
            I => \N__49178\
        );

    \I__12195\ : InMux
    port map (
            O => \N__49237\,
            I => \N__49178\
        );

    \I__12194\ : Span4Mux_h
    port map (
            O => \N__49234\,
            I => \N__49175\
        );

    \I__12193\ : InMux
    port map (
            O => \N__49233\,
            I => \N__49170\
        );

    \I__12192\ : InMux
    port map (
            O => \N__49232\,
            I => \N__49170\
        );

    \I__12191\ : InMux
    port map (
            O => \N__49231\,
            I => \N__49167\
        );

    \I__12190\ : InMux
    port map (
            O => \N__49228\,
            I => \N__49158\
        );

    \I__12189\ : InMux
    port map (
            O => \N__49227\,
            I => \N__49158\
        );

    \I__12188\ : InMux
    port map (
            O => \N__49226\,
            I => \N__49158\
        );

    \I__12187\ : InMux
    port map (
            O => \N__49225\,
            I => \N__49158\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__49222\,
            I => \N__49155\
        );

    \I__12185\ : InMux
    port map (
            O => \N__49221\,
            I => \N__49150\
        );

    \I__12184\ : InMux
    port map (
            O => \N__49220\,
            I => \N__49150\
        );

    \I__12183\ : Span4Mux_h
    port map (
            O => \N__49217\,
            I => \N__49145\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__49214\,
            I => \N__49145\
        );

    \I__12181\ : InMux
    port map (
            O => \N__49213\,
            I => \N__49142\
        );

    \I__12180\ : InMux
    port map (
            O => \N__49212\,
            I => \N__49139\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__49209\,
            I => \N__49136\
        );

    \I__12178\ : InMux
    port map (
            O => \N__49206\,
            I => \N__49131\
        );

    \I__12177\ : InMux
    port map (
            O => \N__49205\,
            I => \N__49131\
        );

    \I__12176\ : CascadeMux
    port map (
            O => \N__49204\,
            I => \N__49125\
        );

    \I__12175\ : CascadeMux
    port map (
            O => \N__49203\,
            I => \N__49115\
        );

    \I__12174\ : CascadeMux
    port map (
            O => \N__49202\,
            I => \N__49112\
        );

    \I__12173\ : InMux
    port map (
            O => \N__49201\,
            I => \N__49102\
        );

    \I__12172\ : InMux
    port map (
            O => \N__49200\,
            I => \N__49102\
        );

    \I__12171\ : InMux
    port map (
            O => \N__49199\,
            I => \N__49095\
        );

    \I__12170\ : InMux
    port map (
            O => \N__49198\,
            I => \N__49095\
        );

    \I__12169\ : InMux
    port map (
            O => \N__49197\,
            I => \N__49095\
        );

    \I__12168\ : InMux
    port map (
            O => \N__49196\,
            I => \N__49090\
        );

    \I__12167\ : InMux
    port map (
            O => \N__49195\,
            I => \N__49090\
        );

    \I__12166\ : InMux
    port map (
            O => \N__49194\,
            I => \N__49079\
        );

    \I__12165\ : InMux
    port map (
            O => \N__49193\,
            I => \N__49079\
        );

    \I__12164\ : InMux
    port map (
            O => \N__49192\,
            I => \N__49079\
        );

    \I__12163\ : InMux
    port map (
            O => \N__49191\,
            I => \N__49079\
        );

    \I__12162\ : InMux
    port map (
            O => \N__49190\,
            I => \N__49079\
        );

    \I__12161\ : InMux
    port map (
            O => \N__49189\,
            I => \N__49074\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__49186\,
            I => \N__49071\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__49183\,
            I => \N__49066\
        );

    \I__12158\ : LocalMux
    port map (
            O => \N__49178\,
            I => \N__49066\
        );

    \I__12157\ : Span4Mux_h
    port map (
            O => \N__49175\,
            I => \N__49061\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__49170\,
            I => \N__49061\
        );

    \I__12155\ : LocalMux
    port map (
            O => \N__49167\,
            I => \N__49056\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__49158\,
            I => \N__49056\
        );

    \I__12153\ : Span4Mux_v
    port map (
            O => \N__49155\,
            I => \N__49049\
        );

    \I__12152\ : LocalMux
    port map (
            O => \N__49150\,
            I => \N__49049\
        );

    \I__12151\ : Span4Mux_v
    port map (
            O => \N__49145\,
            I => \N__49049\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__49142\,
            I => \N__49046\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__49139\,
            I => \N__49043\
        );

    \I__12148\ : Span4Mux_v
    port map (
            O => \N__49136\,
            I => \N__49040\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__49131\,
            I => \N__49037\
        );

    \I__12146\ : InMux
    port map (
            O => \N__49130\,
            I => \N__49030\
        );

    \I__12145\ : InMux
    port map (
            O => \N__49129\,
            I => \N__49030\
        );

    \I__12144\ : InMux
    port map (
            O => \N__49128\,
            I => \N__49030\
        );

    \I__12143\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49024\
        );

    \I__12142\ : InMux
    port map (
            O => \N__49124\,
            I => \N__49024\
        );

    \I__12141\ : InMux
    port map (
            O => \N__49123\,
            I => \N__49021\
        );

    \I__12140\ : InMux
    port map (
            O => \N__49122\,
            I => \N__49013\
        );

    \I__12139\ : InMux
    port map (
            O => \N__49121\,
            I => \N__49013\
        );

    \I__12138\ : InMux
    port map (
            O => \N__49120\,
            I => \N__49013\
        );

    \I__12137\ : CascadeMux
    port map (
            O => \N__49119\,
            I => \N__49008\
        );

    \I__12136\ : InMux
    port map (
            O => \N__49118\,
            I => \N__49004\
        );

    \I__12135\ : InMux
    port map (
            O => \N__49115\,
            I => \N__48993\
        );

    \I__12134\ : InMux
    port map (
            O => \N__49112\,
            I => \N__48993\
        );

    \I__12133\ : InMux
    port map (
            O => \N__49111\,
            I => \N__48993\
        );

    \I__12132\ : InMux
    port map (
            O => \N__49110\,
            I => \N__48993\
        );

    \I__12131\ : InMux
    port map (
            O => \N__49109\,
            I => \N__48993\
        );

    \I__12130\ : InMux
    port map (
            O => \N__49108\,
            I => \N__48988\
        );

    \I__12129\ : InMux
    port map (
            O => \N__49107\,
            I => \N__48988\
        );

    \I__12128\ : LocalMux
    port map (
            O => \N__49102\,
            I => \N__48979\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__49095\,
            I => \N__48979\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__49090\,
            I => \N__48979\
        );

    \I__12125\ : LocalMux
    port map (
            O => \N__49079\,
            I => \N__48979\
        );

    \I__12124\ : InMux
    port map (
            O => \N__49078\,
            I => \N__48972\
        );

    \I__12123\ : InMux
    port map (
            O => \N__49077\,
            I => \N__48972\
        );

    \I__12122\ : LocalMux
    port map (
            O => \N__49074\,
            I => \N__48961\
        );

    \I__12121\ : Span4Mux_v
    port map (
            O => \N__49071\,
            I => \N__48961\
        );

    \I__12120\ : Span4Mux_v
    port map (
            O => \N__49066\,
            I => \N__48961\
        );

    \I__12119\ : Span4Mux_v
    port map (
            O => \N__49061\,
            I => \N__48961\
        );

    \I__12118\ : Span4Mux_v
    port map (
            O => \N__49056\,
            I => \N__48961\
        );

    \I__12117\ : Span4Mux_h
    port map (
            O => \N__49049\,
            I => \N__48958\
        );

    \I__12116\ : Span4Mux_v
    port map (
            O => \N__49046\,
            I => \N__48955\
        );

    \I__12115\ : Span4Mux_v
    port map (
            O => \N__49043\,
            I => \N__48950\
        );

    \I__12114\ : Span4Mux_v
    port map (
            O => \N__49040\,
            I => \N__48950\
        );

    \I__12113\ : Span4Mux_v
    port map (
            O => \N__49037\,
            I => \N__48947\
        );

    \I__12112\ : LocalMux
    port map (
            O => \N__49030\,
            I => \N__48944\
        );

    \I__12111\ : InMux
    port map (
            O => \N__49029\,
            I => \N__48939\
        );

    \I__12110\ : LocalMux
    port map (
            O => \N__49024\,
            I => \N__48936\
        );

    \I__12109\ : LocalMux
    port map (
            O => \N__49021\,
            I => \N__48933\
        );

    \I__12108\ : InMux
    port map (
            O => \N__49020\,
            I => \N__48930\
        );

    \I__12107\ : LocalMux
    port map (
            O => \N__49013\,
            I => \N__48927\
        );

    \I__12106\ : InMux
    port map (
            O => \N__49012\,
            I => \N__48924\
        );

    \I__12105\ : InMux
    port map (
            O => \N__49011\,
            I => \N__48919\
        );

    \I__12104\ : InMux
    port map (
            O => \N__49008\,
            I => \N__48919\
        );

    \I__12103\ : InMux
    port map (
            O => \N__49007\,
            I => \N__48916\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__49004\,
            I => \N__48913\
        );

    \I__12101\ : LocalMux
    port map (
            O => \N__48993\,
            I => \N__48910\
        );

    \I__12100\ : LocalMux
    port map (
            O => \N__48988\,
            I => \N__48905\
        );

    \I__12099\ : Span4Mux_v
    port map (
            O => \N__48979\,
            I => \N__48905\
        );

    \I__12098\ : InMux
    port map (
            O => \N__48978\,
            I => \N__48900\
        );

    \I__12097\ : InMux
    port map (
            O => \N__48977\,
            I => \N__48900\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__48972\,
            I => \N__48889\
        );

    \I__12095\ : Sp12to4
    port map (
            O => \N__48961\,
            I => \N__48889\
        );

    \I__12094\ : Sp12to4
    port map (
            O => \N__48958\,
            I => \N__48889\
        );

    \I__12093\ : Sp12to4
    port map (
            O => \N__48955\,
            I => \N__48889\
        );

    \I__12092\ : Sp12to4
    port map (
            O => \N__48950\,
            I => \N__48889\
        );

    \I__12091\ : Span4Mux_h
    port map (
            O => \N__48947\,
            I => \N__48884\
        );

    \I__12090\ : Span4Mux_h
    port map (
            O => \N__48944\,
            I => \N__48884\
        );

    \I__12089\ : InMux
    port map (
            O => \N__48943\,
            I => \N__48879\
        );

    \I__12088\ : InMux
    port map (
            O => \N__48942\,
            I => \N__48879\
        );

    \I__12087\ : LocalMux
    port map (
            O => \N__48939\,
            I => \N__48868\
        );

    \I__12086\ : Span4Mux_h
    port map (
            O => \N__48936\,
            I => \N__48868\
        );

    \I__12085\ : Span4Mux_v
    port map (
            O => \N__48933\,
            I => \N__48868\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__48930\,
            I => \N__48868\
        );

    \I__12083\ : Span4Mux_h
    port map (
            O => \N__48927\,
            I => \N__48868\
        );

    \I__12082\ : LocalMux
    port map (
            O => \N__48924\,
            I => adc_state_0_adj_1080
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__48919\,
            I => adc_state_0_adj_1080
        );

    \I__12080\ : LocalMux
    port map (
            O => \N__48916\,
            I => adc_state_0_adj_1080
        );

    \I__12079\ : Odrv4
    port map (
            O => \N__48913\,
            I => adc_state_0_adj_1080
        );

    \I__12078\ : Odrv4
    port map (
            O => \N__48910\,
            I => adc_state_0_adj_1080
        );

    \I__12077\ : Odrv4
    port map (
            O => \N__48905\,
            I => adc_state_0_adj_1080
        );

    \I__12076\ : LocalMux
    port map (
            O => \N__48900\,
            I => adc_state_0_adj_1080
        );

    \I__12075\ : Odrv12
    port map (
            O => \N__48889\,
            I => adc_state_0_adj_1080
        );

    \I__12074\ : Odrv4
    port map (
            O => \N__48884\,
            I => adc_state_0_adj_1080
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__48879\,
            I => adc_state_0_adj_1080
        );

    \I__12072\ : Odrv4
    port map (
            O => \N__48868\,
            I => adc_state_0_adj_1080
        );

    \I__12071\ : CascadeMux
    port map (
            O => \N__48845\,
            I => \N__48842\
        );

    \I__12070\ : InMux
    port map (
            O => \N__48842\,
            I => \N__48836\
        );

    \I__12069\ : InMux
    port map (
            O => \N__48841\,
            I => \N__48833\
        );

    \I__12068\ : InMux
    port map (
            O => \N__48840\,
            I => \N__48825\
        );

    \I__12067\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48825\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__48836\,
            I => \N__48819\
        );

    \I__12065\ : LocalMux
    port map (
            O => \N__48833\,
            I => \N__48819\
        );

    \I__12064\ : InMux
    port map (
            O => \N__48832\,
            I => \N__48811\
        );

    \I__12063\ : CascadeMux
    port map (
            O => \N__48831\,
            I => \N__48806\
        );

    \I__12062\ : InMux
    port map (
            O => \N__48830\,
            I => \N__48800\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__48825\,
            I => \N__48797\
        );

    \I__12060\ : InMux
    port map (
            O => \N__48824\,
            I => \N__48794\
        );

    \I__12059\ : Span4Mux_v
    port map (
            O => \N__48819\,
            I => \N__48791\
        );

    \I__12058\ : InMux
    port map (
            O => \N__48818\,
            I => \N__48786\
        );

    \I__12057\ : InMux
    port map (
            O => \N__48817\,
            I => \N__48786\
        );

    \I__12056\ : InMux
    port map (
            O => \N__48816\,
            I => \N__48781\
        );

    \I__12055\ : InMux
    port map (
            O => \N__48815\,
            I => \N__48778\
        );

    \I__12054\ : InMux
    port map (
            O => \N__48814\,
            I => \N__48773\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__48811\,
            I => \N__48770\
        );

    \I__12052\ : InMux
    port map (
            O => \N__48810\,
            I => \N__48767\
        );

    \I__12051\ : InMux
    port map (
            O => \N__48809\,
            I => \N__48764\
        );

    \I__12050\ : InMux
    port map (
            O => \N__48806\,
            I => \N__48758\
        );

    \I__12049\ : InMux
    port map (
            O => \N__48805\,
            I => \N__48758\
        );

    \I__12048\ : InMux
    port map (
            O => \N__48804\,
            I => \N__48752\
        );

    \I__12047\ : InMux
    port map (
            O => \N__48803\,
            I => \N__48749\
        );

    \I__12046\ : LocalMux
    port map (
            O => \N__48800\,
            I => \N__48746\
        );

    \I__12045\ : Span4Mux_h
    port map (
            O => \N__48797\,
            I => \N__48741\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__48794\,
            I => \N__48741\
        );

    \I__12043\ : Span4Mux_h
    port map (
            O => \N__48791\,
            I => \N__48736\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__48786\,
            I => \N__48736\
        );

    \I__12041\ : InMux
    port map (
            O => \N__48785\,
            I => \N__48728\
        );

    \I__12040\ : InMux
    port map (
            O => \N__48784\,
            I => \N__48728\
        );

    \I__12039\ : LocalMux
    port map (
            O => \N__48781\,
            I => \N__48723\
        );

    \I__12038\ : LocalMux
    port map (
            O => \N__48778\,
            I => \N__48723\
        );

    \I__12037\ : InMux
    port map (
            O => \N__48777\,
            I => \N__48718\
        );

    \I__12036\ : InMux
    port map (
            O => \N__48776\,
            I => \N__48718\
        );

    \I__12035\ : LocalMux
    port map (
            O => \N__48773\,
            I => \N__48715\
        );

    \I__12034\ : Span4Mux_v
    port map (
            O => \N__48770\,
            I => \N__48712\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__48767\,
            I => \N__48707\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__48764\,
            I => \N__48707\
        );

    \I__12031\ : InMux
    port map (
            O => \N__48763\,
            I => \N__48704\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__48758\,
            I => \N__48701\
        );

    \I__12029\ : InMux
    port map (
            O => \N__48757\,
            I => \N__48698\
        );

    \I__12028\ : InMux
    port map (
            O => \N__48756\,
            I => \N__48693\
        );

    \I__12027\ : InMux
    port map (
            O => \N__48755\,
            I => \N__48693\
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__48752\,
            I => \N__48686\
        );

    \I__12025\ : LocalMux
    port map (
            O => \N__48749\,
            I => \N__48686\
        );

    \I__12024\ : Span4Mux_h
    port map (
            O => \N__48746\,
            I => \N__48686\
        );

    \I__12023\ : Span4Mux_h
    port map (
            O => \N__48741\,
            I => \N__48681\
        );

    \I__12022\ : Span4Mux_h
    port map (
            O => \N__48736\,
            I => \N__48681\
        );

    \I__12021\ : InMux
    port map (
            O => \N__48735\,
            I => \N__48671\
        );

    \I__12020\ : InMux
    port map (
            O => \N__48734\,
            I => \N__48671\
        );

    \I__12019\ : InMux
    port map (
            O => \N__48733\,
            I => \N__48671\
        );

    \I__12018\ : LocalMux
    port map (
            O => \N__48728\,
            I => \N__48668\
        );

    \I__12017\ : Span4Mux_v
    port map (
            O => \N__48723\,
            I => \N__48661\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__48718\,
            I => \N__48661\
        );

    \I__12015\ : Span4Mux_h
    port map (
            O => \N__48715\,
            I => \N__48661\
        );

    \I__12014\ : Sp12to4
    port map (
            O => \N__48712\,
            I => \N__48658\
        );

    \I__12013\ : Span4Mux_v
    port map (
            O => \N__48707\,
            I => \N__48655\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__48704\,
            I => \N__48652\
        );

    \I__12011\ : Span4Mux_h
    port map (
            O => \N__48701\,
            I => \N__48649\
        );

    \I__12010\ : LocalMux
    port map (
            O => \N__48698\,
            I => \N__48640\
        );

    \I__12009\ : LocalMux
    port map (
            O => \N__48693\,
            I => \N__48640\
        );

    \I__12008\ : Span4Mux_h
    port map (
            O => \N__48686\,
            I => \N__48640\
        );

    \I__12007\ : Span4Mux_v
    port map (
            O => \N__48681\,
            I => \N__48640\
        );

    \I__12006\ : InMux
    port map (
            O => \N__48680\,
            I => \N__48637\
        );

    \I__12005\ : InMux
    port map (
            O => \N__48679\,
            I => \N__48632\
        );

    \I__12004\ : InMux
    port map (
            O => \N__48678\,
            I => \N__48632\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__48671\,
            I => \N__48627\
        );

    \I__12002\ : Span4Mux_h
    port map (
            O => \N__48668\,
            I => \N__48627\
        );

    \I__12001\ : Span4Mux_v
    port map (
            O => \N__48661\,
            I => \N__48624\
        );

    \I__12000\ : Span12Mux_s9_v
    port map (
            O => \N__48658\,
            I => \N__48619\
        );

    \I__11999\ : Sp12to4
    port map (
            O => \N__48655\,
            I => \N__48619\
        );

    \I__11998\ : Span4Mux_v
    port map (
            O => \N__48652\,
            I => \N__48612\
        );

    \I__11997\ : Span4Mux_v
    port map (
            O => \N__48649\,
            I => \N__48612\
        );

    \I__11996\ : Span4Mux_h
    port map (
            O => \N__48640\,
            I => \N__48612\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__48637\,
            I => n8332
        );

    \I__11994\ : LocalMux
    port map (
            O => \N__48632\,
            I => n8332
        );

    \I__11993\ : Odrv4
    port map (
            O => \N__48627\,
            I => n8332
        );

    \I__11992\ : Odrv4
    port map (
            O => \N__48624\,
            I => n8332
        );

    \I__11991\ : Odrv12
    port map (
            O => \N__48619\,
            I => n8332
        );

    \I__11990\ : Odrv4
    port map (
            O => \N__48612\,
            I => n8332
        );

    \I__11989\ : CascadeMux
    port map (
            O => \N__48599\,
            I => \N__48595\
        );

    \I__11988\ : InMux
    port map (
            O => \N__48598\,
            I => \N__48590\
        );

    \I__11987\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48590\
        );

    \I__11986\ : LocalMux
    port map (
            O => \N__48590\,
            I => \N__48586\
        );

    \I__11985\ : CascadeMux
    port map (
            O => \N__48589\,
            I => \N__48583\
        );

    \I__11984\ : Span12Mux_h
    port map (
            O => \N__48586\,
            I => \N__48580\
        );

    \I__11983\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48577\
        );

    \I__11982\ : Odrv12
    port map (
            O => \N__48580\,
            I => cmd_rdadctmp_20_adj_1092
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__48577\,
            I => cmd_rdadctmp_20_adj_1092
        );

    \I__11980\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48569\
        );

    \I__11979\ : LocalMux
    port map (
            O => \N__48569\,
            I => \N__48566\
        );

    \I__11978\ : Odrv12
    port map (
            O => \N__48566\,
            I => n15640
        );

    \I__11977\ : CascadeMux
    port map (
            O => \N__48563\,
            I => \N__48560\
        );

    \I__11976\ : InMux
    port map (
            O => \N__48560\,
            I => \N__48557\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__48557\,
            I => \N__48554\
        );

    \I__11974\ : Span12Mux_v
    port map (
            O => \N__48554\,
            I => \N__48551\
        );

    \I__11973\ : Odrv12
    port map (
            O => \N__48551\,
            I => n10_adj_1172
        );

    \I__11972\ : CEMux
    port map (
            O => \N__48548\,
            I => \N__48539\
        );

    \I__11971\ : CascadeMux
    port map (
            O => \N__48547\,
            I => \N__48533\
        );

    \I__11970\ : CascadeMux
    port map (
            O => \N__48546\,
            I => \N__48530\
        );

    \I__11969\ : InMux
    port map (
            O => \N__48545\,
            I => \N__48510\
        );

    \I__11968\ : InMux
    port map (
            O => \N__48544\,
            I => \N__48510\
        );

    \I__11967\ : InMux
    port map (
            O => \N__48543\,
            I => \N__48510\
        );

    \I__11966\ : InMux
    port map (
            O => \N__48542\,
            I => \N__48507\
        );

    \I__11965\ : LocalMux
    port map (
            O => \N__48539\,
            I => \N__48500\
        );

    \I__11964\ : SRMux
    port map (
            O => \N__48538\,
            I => \N__48497\
        );

    \I__11963\ : InMux
    port map (
            O => \N__48537\,
            I => \N__48494\
        );

    \I__11962\ : InMux
    port map (
            O => \N__48536\,
            I => \N__48477\
        );

    \I__11961\ : InMux
    port map (
            O => \N__48533\,
            I => \N__48477\
        );

    \I__11960\ : InMux
    port map (
            O => \N__48530\,
            I => \N__48477\
        );

    \I__11959\ : InMux
    port map (
            O => \N__48529\,
            I => \N__48477\
        );

    \I__11958\ : InMux
    port map (
            O => \N__48528\,
            I => \N__48477\
        );

    \I__11957\ : InMux
    port map (
            O => \N__48527\,
            I => \N__48477\
        );

    \I__11956\ : InMux
    port map (
            O => \N__48526\,
            I => \N__48477\
        );

    \I__11955\ : InMux
    port map (
            O => \N__48525\,
            I => \N__48477\
        );

    \I__11954\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48460\
        );

    \I__11953\ : InMux
    port map (
            O => \N__48523\,
            I => \N__48460\
        );

    \I__11952\ : InMux
    port map (
            O => \N__48522\,
            I => \N__48460\
        );

    \I__11951\ : InMux
    port map (
            O => \N__48521\,
            I => \N__48460\
        );

    \I__11950\ : InMux
    port map (
            O => \N__48520\,
            I => \N__48460\
        );

    \I__11949\ : InMux
    port map (
            O => \N__48519\,
            I => \N__48460\
        );

    \I__11948\ : InMux
    port map (
            O => \N__48518\,
            I => \N__48460\
        );

    \I__11947\ : InMux
    port map (
            O => \N__48517\,
            I => \N__48460\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__48510\,
            I => \N__48457\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__48507\,
            I => \N__48454\
        );

    \I__11944\ : InMux
    port map (
            O => \N__48506\,
            I => \N__48445\
        );

    \I__11943\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48445\
        );

    \I__11942\ : InMux
    port map (
            O => \N__48504\,
            I => \N__48445\
        );

    \I__11941\ : InMux
    port map (
            O => \N__48503\,
            I => \N__48445\
        );

    \I__11940\ : Span4Mux_v
    port map (
            O => \N__48500\,
            I => \N__48442\
        );

    \I__11939\ : LocalMux
    port map (
            O => \N__48497\,
            I => \N__48439\
        );

    \I__11938\ : LocalMux
    port map (
            O => \N__48494\,
            I => \N__48436\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__48477\,
            I => \N__48431\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__48460\,
            I => \N__48431\
        );

    \I__11935\ : Span4Mux_h
    port map (
            O => \N__48457\,
            I => \N__48424\
        );

    \I__11934\ : Span4Mux_h
    port map (
            O => \N__48454\,
            I => \N__48424\
        );

    \I__11933\ : LocalMux
    port map (
            O => \N__48445\,
            I => \N__48424\
        );

    \I__11932\ : Span4Mux_h
    port map (
            O => \N__48442\,
            I => \N__48421\
        );

    \I__11931\ : Span4Mux_v
    port map (
            O => \N__48439\,
            I => \N__48413\
        );

    \I__11930\ : Span4Mux_h
    port map (
            O => \N__48436\,
            I => \N__48413\
        );

    \I__11929\ : Span4Mux_h
    port map (
            O => \N__48431\,
            I => \N__48413\
        );

    \I__11928\ : Span4Mux_h
    port map (
            O => \N__48424\,
            I => \N__48410\
        );

    \I__11927\ : Span4Mux_v
    port map (
            O => \N__48421\,
            I => \N__48407\
        );

    \I__11926\ : InMux
    port map (
            O => \N__48420\,
            I => \N__48404\
        );

    \I__11925\ : Span4Mux_v
    port map (
            O => \N__48413\,
            I => \N__48401\
        );

    \I__11924\ : Span4Mux_v
    port map (
            O => \N__48410\,
            I => \N__48398\
        );

    \I__11923\ : Odrv4
    port map (
            O => \N__48407\,
            I => dds_state_1
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__48404\,
            I => dds_state_1
        );

    \I__11921\ : Odrv4
    port map (
            O => \N__48401\,
            I => dds_state_1
        );

    \I__11920\ : Odrv4
    port map (
            O => \N__48398\,
            I => dds_state_1
        );

    \I__11919\ : CascadeMux
    port map (
            O => \N__48389\,
            I => \N__48384\
        );

    \I__11918\ : InMux
    port map (
            O => \N__48388\,
            I => \N__48377\
        );

    \I__11917\ : InMux
    port map (
            O => \N__48387\,
            I => \N__48374\
        );

    \I__11916\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48367\
        );

    \I__11915\ : InMux
    port map (
            O => \N__48383\,
            I => \N__48367\
        );

    \I__11914\ : InMux
    port map (
            O => \N__48382\,
            I => \N__48367\
        );

    \I__11913\ : InMux
    port map (
            O => \N__48381\,
            I => \N__48364\
        );

    \I__11912\ : InMux
    port map (
            O => \N__48380\,
            I => \N__48360\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__48377\,
            I => \N__48357\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__48374\,
            I => \N__48352\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48352\
        );

    \I__11908\ : LocalMux
    port map (
            O => \N__48364\,
            I => \N__48349\
        );

    \I__11907\ : InMux
    port map (
            O => \N__48363\,
            I => \N__48346\
        );

    \I__11906\ : LocalMux
    port map (
            O => \N__48360\,
            I => \N__48343\
        );

    \I__11905\ : Span4Mux_v
    port map (
            O => \N__48357\,
            I => \N__48340\
        );

    \I__11904\ : Span4Mux_v
    port map (
            O => \N__48352\,
            I => \N__48335\
        );

    \I__11903\ : Span4Mux_h
    port map (
            O => \N__48349\,
            I => \N__48335\
        );

    \I__11902\ : LocalMux
    port map (
            O => \N__48346\,
            I => \N__48331\
        );

    \I__11901\ : Span4Mux_h
    port map (
            O => \N__48343\,
            I => \N__48328\
        );

    \I__11900\ : Span4Mux_h
    port map (
            O => \N__48340\,
            I => \N__48325\
        );

    \I__11899\ : Span4Mux_h
    port map (
            O => \N__48335\,
            I => \N__48322\
        );

    \I__11898\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48319\
        );

    \I__11897\ : Span12Mux_h
    port map (
            O => \N__48331\,
            I => \N__48316\
        );

    \I__11896\ : Span4Mux_v
    port map (
            O => \N__48328\,
            I => \N__48311\
        );

    \I__11895\ : Span4Mux_h
    port map (
            O => \N__48325\,
            I => \N__48311\
        );

    \I__11894\ : Span4Mux_h
    port map (
            O => \N__48322\,
            I => \N__48308\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__48319\,
            I => dds_state_0
        );

    \I__11892\ : Odrv12
    port map (
            O => \N__48316\,
            I => dds_state_0
        );

    \I__11891\ : Odrv4
    port map (
            O => \N__48311\,
            I => dds_state_0
        );

    \I__11890\ : Odrv4
    port map (
            O => \N__48308\,
            I => dds_state_0
        );

    \I__11889\ : CEMux
    port map (
            O => \N__48299\,
            I => \N__48295\
        );

    \I__11888\ : CEMux
    port map (
            O => \N__48298\,
            I => \N__48292\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__48295\,
            I => \N__48289\
        );

    \I__11886\ : LocalMux
    port map (
            O => \N__48292\,
            I => \N__48286\
        );

    \I__11885\ : Span4Mux_h
    port map (
            O => \N__48289\,
            I => \N__48283\
        );

    \I__11884\ : Span4Mux_h
    port map (
            O => \N__48286\,
            I => \N__48280\
        );

    \I__11883\ : Sp12to4
    port map (
            O => \N__48283\,
            I => \N__48277\
        );

    \I__11882\ : Odrv4
    port map (
            O => \N__48280\,
            I => \CLOCK_DDS.n9\
        );

    \I__11881\ : Odrv12
    port map (
            O => \N__48277\,
            I => \CLOCK_DDS.n9\
        );

    \I__11880\ : CascadeMux
    port map (
            O => \N__48272\,
            I => \N__48269\
        );

    \I__11879\ : InMux
    port map (
            O => \N__48269\,
            I => \N__48266\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__48266\,
            I => \N__48263\
        );

    \I__11877\ : Span4Mux_v
    port map (
            O => \N__48263\,
            I => \N__48260\
        );

    \I__11876\ : Span4Mux_h
    port map (
            O => \N__48260\,
            I => \N__48256\
        );

    \I__11875\ : InMux
    port map (
            O => \N__48259\,
            I => \N__48253\
        );

    \I__11874\ : Span4Mux_h
    port map (
            O => \N__48256\,
            I => \N__48249\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__48253\,
            I => \N__48246\
        );

    \I__11872\ : CascadeMux
    port map (
            O => \N__48252\,
            I => \N__48243\
        );

    \I__11871\ : Span4Mux_h
    port map (
            O => \N__48249\,
            I => \N__48240\
        );

    \I__11870\ : Span4Mux_h
    port map (
            O => \N__48246\,
            I => \N__48237\
        );

    \I__11869\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48234\
        );

    \I__11868\ : Odrv4
    port map (
            O => \N__48240\,
            I => cmd_rdadctmp_24
        );

    \I__11867\ : Odrv4
    port map (
            O => \N__48237\,
            I => cmd_rdadctmp_24
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__48234\,
            I => cmd_rdadctmp_24
        );

    \I__11865\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48223\
        );

    \I__11864\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48220\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__48223\,
            I => \N__48217\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__48220\,
            I => buf_adcdata1_16
        );

    \I__11861\ : Odrv4
    port map (
            O => \N__48217\,
            I => buf_adcdata1_16
        );

    \I__11860\ : InMux
    port map (
            O => \N__48212\,
            I => \N__48209\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__48209\,
            I => \N__48206\
        );

    \I__11858\ : Span4Mux_v
    port map (
            O => \N__48206\,
            I => \N__48203\
        );

    \I__11857\ : Span4Mux_h
    port map (
            O => \N__48203\,
            I => \N__48198\
        );

    \I__11856\ : CascadeMux
    port map (
            O => \N__48202\,
            I => \N__48195\
        );

    \I__11855\ : InMux
    port map (
            O => \N__48201\,
            I => \N__48192\
        );

    \I__11854\ : Span4Mux_h
    port map (
            O => \N__48198\,
            I => \N__48189\
        );

    \I__11853\ : InMux
    port map (
            O => \N__48195\,
            I => \N__48186\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__48192\,
            I => cmd_rdadctmp_30_adj_1046
        );

    \I__11851\ : Odrv4
    port map (
            O => \N__48189\,
            I => cmd_rdadctmp_30_adj_1046
        );

    \I__11850\ : LocalMux
    port map (
            O => \N__48186\,
            I => cmd_rdadctmp_30_adj_1046
        );

    \I__11849\ : InMux
    port map (
            O => \N__48179\,
            I => \N__48176\
        );

    \I__11848\ : LocalMux
    port map (
            O => \N__48176\,
            I => \N__48173\
        );

    \I__11847\ : Span4Mux_v
    port map (
            O => \N__48173\,
            I => \N__48169\
        );

    \I__11846\ : InMux
    port map (
            O => \N__48172\,
            I => \N__48166\
        );

    \I__11845\ : Span4Mux_v
    port map (
            O => \N__48169\,
            I => \N__48163\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__48166\,
            I => buf_adcdata2_22
        );

    \I__11843\ : Odrv4
    port map (
            O => \N__48163\,
            I => buf_adcdata2_22
        );

    \I__11842\ : CascadeMux
    port map (
            O => \N__48158\,
            I => \N__48155\
        );

    \I__11841\ : InMux
    port map (
            O => \N__48155\,
            I => \N__48152\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__48152\,
            I => \N__48149\
        );

    \I__11839\ : Span4Mux_h
    port map (
            O => \N__48149\,
            I => \N__48146\
        );

    \I__11838\ : Span4Mux_h
    port map (
            O => \N__48146\,
            I => \N__48143\
        );

    \I__11837\ : Span4Mux_v
    port map (
            O => \N__48143\,
            I => \N__48140\
        );

    \I__11836\ : Span4Mux_h
    port map (
            O => \N__48140\,
            I => \N__48136\
        );

    \I__11835\ : CascadeMux
    port map (
            O => \N__48139\,
            I => \N__48133\
        );

    \I__11834\ : Span4Mux_h
    port map (
            O => \N__48136\,
            I => \N__48130\
        );

    \I__11833\ : InMux
    port map (
            O => \N__48133\,
            I => \N__48127\
        );

    \I__11832\ : Odrv4
    port map (
            O => \N__48130\,
            I => cmd_rdadctmp_31_adj_1045
        );

    \I__11831\ : LocalMux
    port map (
            O => \N__48127\,
            I => cmd_rdadctmp_31_adj_1045
        );

    \I__11830\ : InMux
    port map (
            O => \N__48122\,
            I => \N__48119\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__48119\,
            I => \N__48115\
        );

    \I__11828\ : InMux
    port map (
            O => \N__48118\,
            I => \N__48112\
        );

    \I__11827\ : Span4Mux_v
    port map (
            O => \N__48115\,
            I => \N__48109\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__48112\,
            I => buf_adcdata2_23
        );

    \I__11825\ : Odrv4
    port map (
            O => \N__48109\,
            I => buf_adcdata2_23
        );

    \I__11824\ : InMux
    port map (
            O => \N__48104\,
            I => \N__48101\
        );

    \I__11823\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__48098\
        );

    \I__11822\ : Span4Mux_v
    port map (
            O => \N__48098\,
            I => \N__48095\
        );

    \I__11821\ : Odrv4
    port map (
            O => \N__48095\,
            I => buf_data2_16
        );

    \I__11820\ : CascadeMux
    port map (
            O => \N__48092\,
            I => \N__48088\
        );

    \I__11819\ : InMux
    port map (
            O => \N__48091\,
            I => \N__48080\
        );

    \I__11818\ : InMux
    port map (
            O => \N__48088\,
            I => \N__48075\
        );

    \I__11817\ : InMux
    port map (
            O => \N__48087\,
            I => \N__48075\
        );

    \I__11816\ : CascadeMux
    port map (
            O => \N__48086\,
            I => \N__48064\
        );

    \I__11815\ : CascadeMux
    port map (
            O => \N__48085\,
            I => \N__48061\
        );

    \I__11814\ : InMux
    port map (
            O => \N__48084\,
            I => \N__48057\
        );

    \I__11813\ : InMux
    port map (
            O => \N__48083\,
            I => \N__48054\
        );

    \I__11812\ : LocalMux
    port map (
            O => \N__48080\,
            I => \N__48049\
        );

    \I__11811\ : LocalMux
    port map (
            O => \N__48075\,
            I => \N__48049\
        );

    \I__11810\ : InMux
    port map (
            O => \N__48074\,
            I => \N__48043\
        );

    \I__11809\ : InMux
    port map (
            O => \N__48073\,
            I => \N__48030\
        );

    \I__11808\ : InMux
    port map (
            O => \N__48072\,
            I => \N__48030\
        );

    \I__11807\ : InMux
    port map (
            O => \N__48071\,
            I => \N__48023\
        );

    \I__11806\ : InMux
    port map (
            O => \N__48070\,
            I => \N__48023\
        );

    \I__11805\ : InMux
    port map (
            O => \N__48069\,
            I => \N__48023\
        );

    \I__11804\ : InMux
    port map (
            O => \N__48068\,
            I => \N__48020\
        );

    \I__11803\ : InMux
    port map (
            O => \N__48067\,
            I => \N__48015\
        );

    \I__11802\ : InMux
    port map (
            O => \N__48064\,
            I => \N__48015\
        );

    \I__11801\ : InMux
    port map (
            O => \N__48061\,
            I => \N__48007\
        );

    \I__11800\ : InMux
    port map (
            O => \N__48060\,
            I => \N__48007\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__48057\,
            I => \N__48001\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__48054\,
            I => \N__47996\
        );

    \I__11797\ : Span4Mux_h
    port map (
            O => \N__48049\,
            I => \N__47996\
        );

    \I__11796\ : InMux
    port map (
            O => \N__48048\,
            I => \N__47993\
        );

    \I__11795\ : CascadeMux
    port map (
            O => \N__48047\,
            I => \N__47990\
        );

    \I__11794\ : CascadeMux
    port map (
            O => \N__48046\,
            I => \N__47986\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__48043\,
            I => \N__47980\
        );

    \I__11792\ : InMux
    port map (
            O => \N__48042\,
            I => \N__47977\
        );

    \I__11791\ : InMux
    port map (
            O => \N__48041\,
            I => \N__47974\
        );

    \I__11790\ : InMux
    port map (
            O => \N__48040\,
            I => \N__47971\
        );

    \I__11789\ : InMux
    port map (
            O => \N__48039\,
            I => \N__47966\
        );

    \I__11788\ : InMux
    port map (
            O => \N__48038\,
            I => \N__47966\
        );

    \I__11787\ : InMux
    port map (
            O => \N__48037\,
            I => \N__47963\
        );

    \I__11786\ : InMux
    port map (
            O => \N__48036\,
            I => \N__47958\
        );

    \I__11785\ : InMux
    port map (
            O => \N__48035\,
            I => \N__47958\
        );

    \I__11784\ : LocalMux
    port map (
            O => \N__48030\,
            I => \N__47955\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__48023\,
            I => \N__47948\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__48020\,
            I => \N__47948\
        );

    \I__11781\ : LocalMux
    port map (
            O => \N__48015\,
            I => \N__47948\
        );

    \I__11780\ : InMux
    port map (
            O => \N__48014\,
            I => \N__47945\
        );

    \I__11779\ : InMux
    port map (
            O => \N__48013\,
            I => \N__47941\
        );

    \I__11778\ : InMux
    port map (
            O => \N__48012\,
            I => \N__47938\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__48007\,
            I => \N__47935\
        );

    \I__11776\ : InMux
    port map (
            O => \N__48006\,
            I => \N__47930\
        );

    \I__11775\ : InMux
    port map (
            O => \N__48005\,
            I => \N__47930\
        );

    \I__11774\ : InMux
    port map (
            O => \N__48004\,
            I => \N__47925\
        );

    \I__11773\ : Span4Mux_v
    port map (
            O => \N__48001\,
            I => \N__47902\
        );

    \I__11772\ : Span4Mux_h
    port map (
            O => \N__47996\,
            I => \N__47902\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__47993\,
            I => \N__47902\
        );

    \I__11770\ : InMux
    port map (
            O => \N__47990\,
            I => \N__47895\
        );

    \I__11769\ : InMux
    port map (
            O => \N__47989\,
            I => \N__47895\
        );

    \I__11768\ : InMux
    port map (
            O => \N__47986\,
            I => \N__47895\
        );

    \I__11767\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47888\
        );

    \I__11766\ : InMux
    port map (
            O => \N__47984\,
            I => \N__47888\
        );

    \I__11765\ : InMux
    port map (
            O => \N__47983\,
            I => \N__47888\
        );

    \I__11764\ : Span4Mux_h
    port map (
            O => \N__47980\,
            I => \N__47877\
        );

    \I__11763\ : LocalMux
    port map (
            O => \N__47977\,
            I => \N__47877\
        );

    \I__11762\ : LocalMux
    port map (
            O => \N__47974\,
            I => \N__47877\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__47971\,
            I => \N__47877\
        );

    \I__11760\ : LocalMux
    port map (
            O => \N__47966\,
            I => \N__47877\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__47963\,
            I => \N__47866\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__47958\,
            I => \N__47866\
        );

    \I__11757\ : Span4Mux_v
    port map (
            O => \N__47955\,
            I => \N__47866\
        );

    \I__11756\ : Span4Mux_v
    port map (
            O => \N__47948\,
            I => \N__47866\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__47945\,
            I => \N__47866\
        );

    \I__11754\ : InMux
    port map (
            O => \N__47944\,
            I => \N__47861\
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__47941\,
            I => \N__47856\
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__47938\,
            I => \N__47849\
        );

    \I__11751\ : Span4Mux_v
    port map (
            O => \N__47935\,
            I => \N__47844\
        );

    \I__11750\ : LocalMux
    port map (
            O => \N__47930\,
            I => \N__47844\
        );

    \I__11749\ : InMux
    port map (
            O => \N__47929\,
            I => \N__47841\
        );

    \I__11748\ : InMux
    port map (
            O => \N__47928\,
            I => \N__47838\
        );

    \I__11747\ : LocalMux
    port map (
            O => \N__47925\,
            I => \N__47835\
        );

    \I__11746\ : InMux
    port map (
            O => \N__47924\,
            I => \N__47828\
        );

    \I__11745\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47828\
        );

    \I__11744\ : InMux
    port map (
            O => \N__47922\,
            I => \N__47828\
        );

    \I__11743\ : InMux
    port map (
            O => \N__47921\,
            I => \N__47825\
        );

    \I__11742\ : InMux
    port map (
            O => \N__47920\,
            I => \N__47817\
        );

    \I__11741\ : InMux
    port map (
            O => \N__47919\,
            I => \N__47817\
        );

    \I__11740\ : CascadeMux
    port map (
            O => \N__47918\,
            I => \N__47812\
        );

    \I__11739\ : InMux
    port map (
            O => \N__47917\,
            I => \N__47807\
        );

    \I__11738\ : InMux
    port map (
            O => \N__47916\,
            I => \N__47787\
        );

    \I__11737\ : InMux
    port map (
            O => \N__47915\,
            I => \N__47776\
        );

    \I__11736\ : InMux
    port map (
            O => \N__47914\,
            I => \N__47776\
        );

    \I__11735\ : InMux
    port map (
            O => \N__47913\,
            I => \N__47776\
        );

    \I__11734\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47776\
        );

    \I__11733\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47776\
        );

    \I__11732\ : InMux
    port map (
            O => \N__47910\,
            I => \N__47771\
        );

    \I__11731\ : InMux
    port map (
            O => \N__47909\,
            I => \N__47771\
        );

    \I__11730\ : Span4Mux_h
    port map (
            O => \N__47902\,
            I => \N__47764\
        );

    \I__11729\ : LocalMux
    port map (
            O => \N__47895\,
            I => \N__47764\
        );

    \I__11728\ : LocalMux
    port map (
            O => \N__47888\,
            I => \N__47764\
        );

    \I__11727\ : Span4Mux_v
    port map (
            O => \N__47877\,
            I => \N__47759\
        );

    \I__11726\ : Span4Mux_h
    port map (
            O => \N__47866\,
            I => \N__47759\
        );

    \I__11725\ : InMux
    port map (
            O => \N__47865\,
            I => \N__47754\
        );

    \I__11724\ : InMux
    port map (
            O => \N__47864\,
            I => \N__47754\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__47861\,
            I => \N__47751\
        );

    \I__11722\ : InMux
    port map (
            O => \N__47860\,
            I => \N__47746\
        );

    \I__11721\ : InMux
    port map (
            O => \N__47859\,
            I => \N__47746\
        );

    \I__11720\ : Span4Mux_h
    port map (
            O => \N__47856\,
            I => \N__47738\
        );

    \I__11719\ : InMux
    port map (
            O => \N__47855\,
            I => \N__47735\
        );

    \I__11718\ : InMux
    port map (
            O => \N__47854\,
            I => \N__47732\
        );

    \I__11717\ : InMux
    port map (
            O => \N__47853\,
            I => \N__47727\
        );

    \I__11716\ : InMux
    port map (
            O => \N__47852\,
            I => \N__47727\
        );

    \I__11715\ : Span4Mux_v
    port map (
            O => \N__47849\,
            I => \N__47722\
        );

    \I__11714\ : Span4Mux_h
    port map (
            O => \N__47844\,
            I => \N__47722\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__47841\,
            I => \N__47719\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__47838\,
            I => \N__47716\
        );

    \I__11711\ : Span4Mux_h
    port map (
            O => \N__47835\,
            I => \N__47711\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__47828\,
            I => \N__47711\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__47825\,
            I => \N__47708\
        );

    \I__11708\ : InMux
    port map (
            O => \N__47824\,
            I => \N__47703\
        );

    \I__11707\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47703\
        );

    \I__11706\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47697\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__47817\,
            I => \N__47694\
        );

    \I__11704\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47687\
        );

    \I__11703\ : InMux
    port map (
            O => \N__47815\,
            I => \N__47687\
        );

    \I__11702\ : InMux
    port map (
            O => \N__47812\,
            I => \N__47687\
        );

    \I__11701\ : InMux
    port map (
            O => \N__47811\,
            I => \N__47684\
        );

    \I__11700\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47681\
        );

    \I__11699\ : LocalMux
    port map (
            O => \N__47807\,
            I => \N__47678\
        );

    \I__11698\ : InMux
    port map (
            O => \N__47806\,
            I => \N__47671\
        );

    \I__11697\ : InMux
    port map (
            O => \N__47805\,
            I => \N__47671\
        );

    \I__11696\ : InMux
    port map (
            O => \N__47804\,
            I => \N__47671\
        );

    \I__11695\ : InMux
    port map (
            O => \N__47803\,
            I => \N__47667\
        );

    \I__11694\ : InMux
    port map (
            O => \N__47802\,
            I => \N__47664\
        );

    \I__11693\ : InMux
    port map (
            O => \N__47801\,
            I => \N__47659\
        );

    \I__11692\ : InMux
    port map (
            O => \N__47800\,
            I => \N__47659\
        );

    \I__11691\ : InMux
    port map (
            O => \N__47799\,
            I => \N__47654\
        );

    \I__11690\ : InMux
    port map (
            O => \N__47798\,
            I => \N__47654\
        );

    \I__11689\ : InMux
    port map (
            O => \N__47797\,
            I => \N__47647\
        );

    \I__11688\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47647\
        );

    \I__11687\ : InMux
    port map (
            O => \N__47795\,
            I => \N__47647\
        );

    \I__11686\ : InMux
    port map (
            O => \N__47794\,
            I => \N__47640\
        );

    \I__11685\ : InMux
    port map (
            O => \N__47793\,
            I => \N__47640\
        );

    \I__11684\ : InMux
    port map (
            O => \N__47792\,
            I => \N__47640\
        );

    \I__11683\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47637\
        );

    \I__11682\ : CascadeMux
    port map (
            O => \N__47790\,
            I => \N__47633\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__47787\,
            I => \N__47620\
        );

    \I__11680\ : LocalMux
    port map (
            O => \N__47776\,
            I => \N__47620\
        );

    \I__11679\ : LocalMux
    port map (
            O => \N__47771\,
            I => \N__47620\
        );

    \I__11678\ : Span4Mux_v
    port map (
            O => \N__47764\,
            I => \N__47620\
        );

    \I__11677\ : Span4Mux_h
    port map (
            O => \N__47759\,
            I => \N__47620\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__47754\,
            I => \N__47620\
        );

    \I__11675\ : Span4Mux_h
    port map (
            O => \N__47751\,
            I => \N__47615\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__47746\,
            I => \N__47615\
        );

    \I__11673\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47606\
        );

    \I__11672\ : InMux
    port map (
            O => \N__47744\,
            I => \N__47606\
        );

    \I__11671\ : InMux
    port map (
            O => \N__47743\,
            I => \N__47606\
        );

    \I__11670\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47606\
        );

    \I__11669\ : CascadeMux
    port map (
            O => \N__47741\,
            I => \N__47596\
        );

    \I__11668\ : Span4Mux_h
    port map (
            O => \N__47738\,
            I => \N__47588\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__47735\,
            I => \N__47588\
        );

    \I__11666\ : LocalMux
    port map (
            O => \N__47732\,
            I => \N__47585\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__47727\,
            I => \N__47580\
        );

    \I__11664\ : Span4Mux_h
    port map (
            O => \N__47722\,
            I => \N__47580\
        );

    \I__11663\ : Span4Mux_h
    port map (
            O => \N__47719\,
            I => \N__47577\
        );

    \I__11662\ : Span4Mux_v
    port map (
            O => \N__47716\,
            I => \N__47572\
        );

    \I__11661\ : Span4Mux_h
    port map (
            O => \N__47711\,
            I => \N__47572\
        );

    \I__11660\ : Span4Mux_h
    port map (
            O => \N__47708\,
            I => \N__47567\
        );

    \I__11659\ : LocalMux
    port map (
            O => \N__47703\,
            I => \N__47567\
        );

    \I__11658\ : InMux
    port map (
            O => \N__47702\,
            I => \N__47564\
        );

    \I__11657\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47559\
        );

    \I__11656\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47559\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__47697\,
            I => \N__47544\
        );

    \I__11654\ : Span4Mux_h
    port map (
            O => \N__47694\,
            I => \N__47544\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__47687\,
            I => \N__47544\
        );

    \I__11652\ : LocalMux
    port map (
            O => \N__47684\,
            I => \N__47544\
        );

    \I__11651\ : LocalMux
    port map (
            O => \N__47681\,
            I => \N__47544\
        );

    \I__11650\ : Span4Mux_h
    port map (
            O => \N__47678\,
            I => \N__47544\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__47671\,
            I => \N__47544\
        );

    \I__11648\ : CascadeMux
    port map (
            O => \N__47670\,
            I => \N__47537\
        );

    \I__11647\ : LocalMux
    port map (
            O => \N__47667\,
            I => \N__47522\
        );

    \I__11646\ : LocalMux
    port map (
            O => \N__47664\,
            I => \N__47522\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__47659\,
            I => \N__47522\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__47654\,
            I => \N__47522\
        );

    \I__11643\ : LocalMux
    port map (
            O => \N__47647\,
            I => \N__47522\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__47640\,
            I => \N__47522\
        );

    \I__11641\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47522\
        );

    \I__11640\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47517\
        );

    \I__11639\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47517\
        );

    \I__11638\ : Span4Mux_v
    port map (
            O => \N__47620\,
            I => \N__47510\
        );

    \I__11637\ : Span4Mux_v
    port map (
            O => \N__47615\,
            I => \N__47510\
        );

    \I__11636\ : LocalMux
    port map (
            O => \N__47606\,
            I => \N__47510\
        );

    \I__11635\ : InMux
    port map (
            O => \N__47605\,
            I => \N__47504\
        );

    \I__11634\ : InMux
    port map (
            O => \N__47604\,
            I => \N__47497\
        );

    \I__11633\ : InMux
    port map (
            O => \N__47603\,
            I => \N__47497\
        );

    \I__11632\ : InMux
    port map (
            O => \N__47602\,
            I => \N__47497\
        );

    \I__11631\ : CascadeMux
    port map (
            O => \N__47601\,
            I => \N__47492\
        );

    \I__11630\ : InMux
    port map (
            O => \N__47600\,
            I => \N__47485\
        );

    \I__11629\ : InMux
    port map (
            O => \N__47599\,
            I => \N__47480\
        );

    \I__11628\ : InMux
    port map (
            O => \N__47596\,
            I => \N__47480\
        );

    \I__11627\ : InMux
    port map (
            O => \N__47595\,
            I => \N__47473\
        );

    \I__11626\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47473\
        );

    \I__11625\ : InMux
    port map (
            O => \N__47593\,
            I => \N__47473\
        );

    \I__11624\ : Span4Mux_h
    port map (
            O => \N__47588\,
            I => \N__47470\
        );

    \I__11623\ : Span4Mux_h
    port map (
            O => \N__47585\,
            I => \N__47459\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__47580\,
            I => \N__47459\
        );

    \I__11621\ : Span4Mux_v
    port map (
            O => \N__47577\,
            I => \N__47459\
        );

    \I__11620\ : Span4Mux_v
    port map (
            O => \N__47572\,
            I => \N__47459\
        );

    \I__11619\ : Span4Mux_h
    port map (
            O => \N__47567\,
            I => \N__47459\
        );

    \I__11618\ : LocalMux
    port map (
            O => \N__47564\,
            I => \N__47452\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__47559\,
            I => \N__47452\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__47544\,
            I => \N__47452\
        );

    \I__11615\ : InMux
    port map (
            O => \N__47543\,
            I => \N__47447\
        );

    \I__11614\ : InMux
    port map (
            O => \N__47542\,
            I => \N__47447\
        );

    \I__11613\ : InMux
    port map (
            O => \N__47541\,
            I => \N__47440\
        );

    \I__11612\ : InMux
    port map (
            O => \N__47540\,
            I => \N__47440\
        );

    \I__11611\ : InMux
    port map (
            O => \N__47537\,
            I => \N__47440\
        );

    \I__11610\ : Span4Mux_v
    port map (
            O => \N__47522\,
            I => \N__47433\
        );

    \I__11609\ : LocalMux
    port map (
            O => \N__47517\,
            I => \N__47433\
        );

    \I__11608\ : Span4Mux_h
    port map (
            O => \N__47510\,
            I => \N__47433\
        );

    \I__11607\ : InMux
    port map (
            O => \N__47509\,
            I => \N__47426\
        );

    \I__11606\ : InMux
    port map (
            O => \N__47508\,
            I => \N__47426\
        );

    \I__11605\ : InMux
    port map (
            O => \N__47507\,
            I => \N__47426\
        );

    \I__11604\ : LocalMux
    port map (
            O => \N__47504\,
            I => \N__47421\
        );

    \I__11603\ : LocalMux
    port map (
            O => \N__47497\,
            I => \N__47421\
        );

    \I__11602\ : InMux
    port map (
            O => \N__47496\,
            I => \N__47412\
        );

    \I__11601\ : InMux
    port map (
            O => \N__47495\,
            I => \N__47412\
        );

    \I__11600\ : InMux
    port map (
            O => \N__47492\,
            I => \N__47412\
        );

    \I__11599\ : InMux
    port map (
            O => \N__47491\,
            I => \N__47412\
        );

    \I__11598\ : InMux
    port map (
            O => \N__47490\,
            I => \N__47405\
        );

    \I__11597\ : InMux
    port map (
            O => \N__47489\,
            I => \N__47405\
        );

    \I__11596\ : InMux
    port map (
            O => \N__47488\,
            I => \N__47405\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__47485\,
            I => comm_cmd_0
        );

    \I__11594\ : LocalMux
    port map (
            O => \N__47480\,
            I => comm_cmd_0
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__47473\,
            I => comm_cmd_0
        );

    \I__11592\ : Odrv4
    port map (
            O => \N__47470\,
            I => comm_cmd_0
        );

    \I__11591\ : Odrv4
    port map (
            O => \N__47459\,
            I => comm_cmd_0
        );

    \I__11590\ : Odrv4
    port map (
            O => \N__47452\,
            I => comm_cmd_0
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__47447\,
            I => comm_cmd_0
        );

    \I__11588\ : LocalMux
    port map (
            O => \N__47440\,
            I => comm_cmd_0
        );

    \I__11587\ : Odrv4
    port map (
            O => \N__47433\,
            I => comm_cmd_0
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__47426\,
            I => comm_cmd_0
        );

    \I__11585\ : Odrv4
    port map (
            O => \N__47421\,
            I => comm_cmd_0
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__47412\,
            I => comm_cmd_0
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__47405\,
            I => comm_cmd_0
        );

    \I__11582\ : CascadeMux
    port map (
            O => \N__47378\,
            I => \N__47375\
        );

    \I__11581\ : InMux
    port map (
            O => \N__47375\,
            I => \N__47372\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__47372\,
            I => \N__47368\
        );

    \I__11579\ : InMux
    port map (
            O => \N__47371\,
            I => \N__47365\
        );

    \I__11578\ : Span4Mux_v
    port map (
            O => \N__47368\,
            I => \N__47360\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__47365\,
            I => \N__47360\
        );

    \I__11576\ : Span4Mux_v
    port map (
            O => \N__47360\,
            I => \N__47356\
        );

    \I__11575\ : CascadeMux
    port map (
            O => \N__47359\,
            I => \N__47353\
        );

    \I__11574\ : Span4Mux_h
    port map (
            O => \N__47356\,
            I => \N__47350\
        );

    \I__11573\ : InMux
    port map (
            O => \N__47353\,
            I => \N__47347\
        );

    \I__11572\ : Span4Mux_h
    port map (
            O => \N__47350\,
            I => \N__47344\
        );

    \I__11571\ : LocalMux
    port map (
            O => \N__47347\,
            I => buf_adcdata4_16
        );

    \I__11570\ : Odrv4
    port map (
            O => \N__47344\,
            I => buf_adcdata4_16
        );

    \I__11569\ : InMux
    port map (
            O => \N__47339\,
            I => \N__47330\
        );

    \I__11568\ : InMux
    port map (
            O => \N__47338\,
            I => \N__47330\
        );

    \I__11567\ : InMux
    port map (
            O => \N__47337\,
            I => \N__47327\
        );

    \I__11566\ : CascadeMux
    port map (
            O => \N__47336\,
            I => \N__47316\
        );

    \I__11565\ : InMux
    port map (
            O => \N__47335\,
            I => \N__47312\
        );

    \I__11564\ : LocalMux
    port map (
            O => \N__47330\,
            I => \N__47304\
        );

    \I__11563\ : LocalMux
    port map (
            O => \N__47327\,
            I => \N__47301\
        );

    \I__11562\ : InMux
    port map (
            O => \N__47326\,
            I => \N__47294\
        );

    \I__11561\ : InMux
    port map (
            O => \N__47325\,
            I => \N__47294\
        );

    \I__11560\ : InMux
    port map (
            O => \N__47324\,
            I => \N__47294\
        );

    \I__11559\ : InMux
    port map (
            O => \N__47323\,
            I => \N__47285\
        );

    \I__11558\ : InMux
    port map (
            O => \N__47322\,
            I => \N__47285\
        );

    \I__11557\ : InMux
    port map (
            O => \N__47321\,
            I => \N__47278\
        );

    \I__11556\ : InMux
    port map (
            O => \N__47320\,
            I => \N__47278\
        );

    \I__11555\ : InMux
    port map (
            O => \N__47319\,
            I => \N__47278\
        );

    \I__11554\ : InMux
    port map (
            O => \N__47316\,
            I => \N__47275\
        );

    \I__11553\ : CascadeMux
    port map (
            O => \N__47315\,
            I => \N__47269\
        );

    \I__11552\ : LocalMux
    port map (
            O => \N__47312\,
            I => \N__47263\
        );

    \I__11551\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47257\
        );

    \I__11550\ : InMux
    port map (
            O => \N__47310\,
            I => \N__47240\
        );

    \I__11549\ : CascadeMux
    port map (
            O => \N__47309\,
            I => \N__47233\
        );

    \I__11548\ : InMux
    port map (
            O => \N__47308\,
            I => \N__47227\
        );

    \I__11547\ : CascadeMux
    port map (
            O => \N__47307\,
            I => \N__47224\
        );

    \I__11546\ : Span4Mux_h
    port map (
            O => \N__47304\,
            I => \N__47217\
        );

    \I__11545\ : Span4Mux_v
    port map (
            O => \N__47301\,
            I => \N__47217\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__47294\,
            I => \N__47217\
        );

    \I__11543\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47214\
        );

    \I__11542\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47209\
        );

    \I__11541\ : InMux
    port map (
            O => \N__47291\,
            I => \N__47209\
        );

    \I__11540\ : InMux
    port map (
            O => \N__47290\,
            I => \N__47206\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__47285\,
            I => \N__47199\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__47278\,
            I => \N__47199\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__47275\,
            I => \N__47199\
        );

    \I__11536\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47196\
        );

    \I__11535\ : InMux
    port map (
            O => \N__47273\,
            I => \N__47191\
        );

    \I__11534\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47191\
        );

    \I__11533\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47188\
        );

    \I__11532\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47185\
        );

    \I__11531\ : InMux
    port map (
            O => \N__47267\,
            I => \N__47178\
        );

    \I__11530\ : InMux
    port map (
            O => \N__47266\,
            I => \N__47175\
        );

    \I__11529\ : Span4Mux_v
    port map (
            O => \N__47263\,
            I => \N__47170\
        );

    \I__11528\ : InMux
    port map (
            O => \N__47262\,
            I => \N__47163\
        );

    \I__11527\ : InMux
    port map (
            O => \N__47261\,
            I => \N__47163\
        );

    \I__11526\ : InMux
    port map (
            O => \N__47260\,
            I => \N__47163\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__47257\,
            I => \N__47160\
        );

    \I__11524\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47153\
        );

    \I__11523\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47153\
        );

    \I__11522\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47153\
        );

    \I__11521\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47143\
        );

    \I__11520\ : InMux
    port map (
            O => \N__47252\,
            I => \N__47143\
        );

    \I__11519\ : InMux
    port map (
            O => \N__47251\,
            I => \N__47143\
        );

    \I__11518\ : InMux
    port map (
            O => \N__47250\,
            I => \N__47134\
        );

    \I__11517\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47127\
        );

    \I__11516\ : InMux
    port map (
            O => \N__47248\,
            I => \N__47127\
        );

    \I__11515\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47127\
        );

    \I__11514\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47124\
        );

    \I__11513\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47121\
        );

    \I__11512\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47116\
        );

    \I__11511\ : InMux
    port map (
            O => \N__47243\,
            I => \N__47116\
        );

    \I__11510\ : LocalMux
    port map (
            O => \N__47240\,
            I => \N__47113\
        );

    \I__11509\ : InMux
    port map (
            O => \N__47239\,
            I => \N__47110\
        );

    \I__11508\ : InMux
    port map (
            O => \N__47238\,
            I => \N__47107\
        );

    \I__11507\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47102\
        );

    \I__11506\ : InMux
    port map (
            O => \N__47236\,
            I => \N__47102\
        );

    \I__11505\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47099\
        );

    \I__11504\ : CascadeMux
    port map (
            O => \N__47232\,
            I => \N__47096\
        );

    \I__11503\ : InMux
    port map (
            O => \N__47231\,
            I => \N__47089\
        );

    \I__11502\ : InMux
    port map (
            O => \N__47230\,
            I => \N__47089\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__47227\,
            I => \N__47081\
        );

    \I__11500\ : InMux
    port map (
            O => \N__47224\,
            I => \N__47078\
        );

    \I__11499\ : Span4Mux_h
    port map (
            O => \N__47217\,
            I => \N__47072\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__47214\,
            I => \N__47072\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__47209\,
            I => \N__47065\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__47206\,
            I => \N__47065\
        );

    \I__11495\ : Span4Mux_v
    port map (
            O => \N__47199\,
            I => \N__47065\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__47196\,
            I => \N__47060\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__47191\,
            I => \N__47060\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__47188\,
            I => \N__47055\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__47185\,
            I => \N__47055\
        );

    \I__11490\ : CascadeMux
    port map (
            O => \N__47184\,
            I => \N__47052\
        );

    \I__11489\ : CascadeMux
    port map (
            O => \N__47183\,
            I => \N__47049\
        );

    \I__11488\ : CascadeMux
    port map (
            O => \N__47182\,
            I => \N__47043\
        );

    \I__11487\ : CascadeMux
    port map (
            O => \N__47181\,
            I => \N__47040\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__47178\,
            I => \N__47037\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__47175\,
            I => \N__47034\
        );

    \I__11484\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47031\
        );

    \I__11483\ : InMux
    port map (
            O => \N__47173\,
            I => \N__47028\
        );

    \I__11482\ : Span4Mux_v
    port map (
            O => \N__47170\,
            I => \N__47018\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__47163\,
            I => \N__47018\
        );

    \I__11480\ : Span4Mux_v
    port map (
            O => \N__47160\,
            I => \N__47018\
        );

    \I__11479\ : LocalMux
    port map (
            O => \N__47153\,
            I => \N__47018\
        );

    \I__11478\ : InMux
    port map (
            O => \N__47152\,
            I => \N__47011\
        );

    \I__11477\ : InMux
    port map (
            O => \N__47151\,
            I => \N__47011\
        );

    \I__11476\ : InMux
    port map (
            O => \N__47150\,
            I => \N__47011\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__47143\,
            I => \N__47008\
        );

    \I__11474\ : InMux
    port map (
            O => \N__47142\,
            I => \N__47001\
        );

    \I__11473\ : InMux
    port map (
            O => \N__47141\,
            I => \N__47001\
        );

    \I__11472\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47001\
        );

    \I__11471\ : InMux
    port map (
            O => \N__47139\,
            I => \N__46994\
        );

    \I__11470\ : InMux
    port map (
            O => \N__47138\,
            I => \N__46994\
        );

    \I__11469\ : InMux
    port map (
            O => \N__47137\,
            I => \N__46994\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__47134\,
            I => \N__46977\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__47127\,
            I => \N__46977\
        );

    \I__11466\ : LocalMux
    port map (
            O => \N__47124\,
            I => \N__46977\
        );

    \I__11465\ : LocalMux
    port map (
            O => \N__47121\,
            I => \N__46977\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__47116\,
            I => \N__46977\
        );

    \I__11463\ : Span4Mux_v
    port map (
            O => \N__47113\,
            I => \N__46977\
        );

    \I__11462\ : LocalMux
    port map (
            O => \N__47110\,
            I => \N__46977\
        );

    \I__11461\ : LocalMux
    port map (
            O => \N__47107\,
            I => \N__46977\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__47102\,
            I => \N__46972\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__46972\
        );

    \I__11458\ : InMux
    port map (
            O => \N__47096\,
            I => \N__46967\
        );

    \I__11457\ : InMux
    port map (
            O => \N__47095\,
            I => \N__46967\
        );

    \I__11456\ : InMux
    port map (
            O => \N__47094\,
            I => \N__46960\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__47089\,
            I => \N__46957\
        );

    \I__11454\ : InMux
    port map (
            O => \N__47088\,
            I => \N__46952\
        );

    \I__11453\ : InMux
    port map (
            O => \N__47087\,
            I => \N__46952\
        );

    \I__11452\ : InMux
    port map (
            O => \N__47086\,
            I => \N__46947\
        );

    \I__11451\ : InMux
    port map (
            O => \N__47085\,
            I => \N__46947\
        );

    \I__11450\ : InMux
    port map (
            O => \N__47084\,
            I => \N__46943\
        );

    \I__11449\ : Span4Mux_v
    port map (
            O => \N__47081\,
            I => \N__46938\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__47078\,
            I => \N__46938\
        );

    \I__11447\ : InMux
    port map (
            O => \N__47077\,
            I => \N__46935\
        );

    \I__11446\ : Span4Mux_h
    port map (
            O => \N__47072\,
            I => \N__46932\
        );

    \I__11445\ : Span4Mux_h
    port map (
            O => \N__47065\,
            I => \N__46924\
        );

    \I__11444\ : Span4Mux_v
    port map (
            O => \N__47060\,
            I => \N__46924\
        );

    \I__11443\ : Span4Mux_v
    port map (
            O => \N__47055\,
            I => \N__46924\
        );

    \I__11442\ : InMux
    port map (
            O => \N__47052\,
            I => \N__46917\
        );

    \I__11441\ : InMux
    port map (
            O => \N__47049\,
            I => \N__46917\
        );

    \I__11440\ : InMux
    port map (
            O => \N__47048\,
            I => \N__46917\
        );

    \I__11439\ : InMux
    port map (
            O => \N__47047\,
            I => \N__46912\
        );

    \I__11438\ : InMux
    port map (
            O => \N__47046\,
            I => \N__46912\
        );

    \I__11437\ : InMux
    port map (
            O => \N__47043\,
            I => \N__46905\
        );

    \I__11436\ : InMux
    port map (
            O => \N__47040\,
            I => \N__46902\
        );

    \I__11435\ : Span4Mux_h
    port map (
            O => \N__47037\,
            I => \N__46899\
        );

    \I__11434\ : Span4Mux_h
    port map (
            O => \N__47034\,
            I => \N__46891\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__47031\,
            I => \N__46891\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__47028\,
            I => \N__46891\
        );

    \I__11431\ : InMux
    port map (
            O => \N__47027\,
            I => \N__46888\
        );

    \I__11430\ : Span4Mux_h
    port map (
            O => \N__47018\,
            I => \N__46875\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__47011\,
            I => \N__46875\
        );

    \I__11428\ : Span4Mux_v
    port map (
            O => \N__47008\,
            I => \N__46875\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__47001\,
            I => \N__46875\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__46994\,
            I => \N__46875\
        );

    \I__11425\ : Span4Mux_v
    port map (
            O => \N__46977\,
            I => \N__46875\
        );

    \I__11424\ : Span4Mux_v
    port map (
            O => \N__46972\,
            I => \N__46870\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__46967\,
            I => \N__46870\
        );

    \I__11422\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46867\
        );

    \I__11421\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46864\
        );

    \I__11420\ : InMux
    port map (
            O => \N__46964\,
            I => \N__46861\
        );

    \I__11419\ : InMux
    port map (
            O => \N__46963\,
            I => \N__46858\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__46960\,
            I => \N__46855\
        );

    \I__11417\ : Sp12to4
    port map (
            O => \N__46957\,
            I => \N__46848\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__46952\,
            I => \N__46848\
        );

    \I__11415\ : LocalMux
    port map (
            O => \N__46947\,
            I => \N__46848\
        );

    \I__11414\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46845\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__46943\,
            I => \N__46842\
        );

    \I__11412\ : Sp12to4
    port map (
            O => \N__46938\,
            I => \N__46839\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__46935\,
            I => \N__46836\
        );

    \I__11410\ : Span4Mux_h
    port map (
            O => \N__46932\,
            I => \N__46830\
        );

    \I__11409\ : InMux
    port map (
            O => \N__46931\,
            I => \N__46827\
        );

    \I__11408\ : Span4Mux_h
    port map (
            O => \N__46924\,
            I => \N__46820\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__46917\,
            I => \N__46820\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__46912\,
            I => \N__46820\
        );

    \I__11405\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46814\
        );

    \I__11404\ : InMux
    port map (
            O => \N__46910\,
            I => \N__46811\
        );

    \I__11403\ : InMux
    port map (
            O => \N__46909\,
            I => \N__46806\
        );

    \I__11402\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46806\
        );

    \I__11401\ : LocalMux
    port map (
            O => \N__46905\,
            I => \N__46799\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__46902\,
            I => \N__46799\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__46899\,
            I => \N__46799\
        );

    \I__11398\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46796\
        );

    \I__11397\ : Span4Mux_v
    port map (
            O => \N__46891\,
            I => \N__46787\
        );

    \I__11396\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46787\
        );

    \I__11395\ : Span4Mux_h
    port map (
            O => \N__46875\,
            I => \N__46787\
        );

    \I__11394\ : Span4Mux_v
    port map (
            O => \N__46870\,
            I => \N__46787\
        );

    \I__11393\ : LocalMux
    port map (
            O => \N__46867\,
            I => \N__46772\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__46864\,
            I => \N__46772\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__46861\,
            I => \N__46772\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__46858\,
            I => \N__46772\
        );

    \I__11389\ : Span12Mux_s10_h
    port map (
            O => \N__46855\,
            I => \N__46772\
        );

    \I__11388\ : Span12Mux_h
    port map (
            O => \N__46848\,
            I => \N__46772\
        );

    \I__11387\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46772\
        );

    \I__11386\ : Span12Mux_v
    port map (
            O => \N__46842\,
            I => \N__46765\
        );

    \I__11385\ : Span12Mux_v
    port map (
            O => \N__46839\,
            I => \N__46765\
        );

    \I__11384\ : Span12Mux_h
    port map (
            O => \N__46836\,
            I => \N__46765\
        );

    \I__11383\ : InMux
    port map (
            O => \N__46835\,
            I => \N__46758\
        );

    \I__11382\ : InMux
    port map (
            O => \N__46834\,
            I => \N__46758\
        );

    \I__11381\ : InMux
    port map (
            O => \N__46833\,
            I => \N__46758\
        );

    \I__11380\ : Span4Mux_v
    port map (
            O => \N__46830\,
            I => \N__46751\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__46827\,
            I => \N__46751\
        );

    \I__11378\ : Span4Mux_h
    port map (
            O => \N__46820\,
            I => \N__46751\
        );

    \I__11377\ : InMux
    port map (
            O => \N__46819\,
            I => \N__46748\
        );

    \I__11376\ : InMux
    port map (
            O => \N__46818\,
            I => \N__46743\
        );

    \I__11375\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46743\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__46814\,
            I => comm_cmd_3
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__46811\,
            I => comm_cmd_3
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__46806\,
            I => comm_cmd_3
        );

    \I__11371\ : Odrv4
    port map (
            O => \N__46799\,
            I => comm_cmd_3
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__46796\,
            I => comm_cmd_3
        );

    \I__11369\ : Odrv4
    port map (
            O => \N__46787\,
            I => comm_cmd_3
        );

    \I__11368\ : Odrv12
    port map (
            O => \N__46772\,
            I => comm_cmd_3
        );

    \I__11367\ : Odrv12
    port map (
            O => \N__46765\,
            I => comm_cmd_3
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__46758\,
            I => comm_cmd_3
        );

    \I__11365\ : Odrv4
    port map (
            O => \N__46751\,
            I => comm_cmd_3
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__46748\,
            I => comm_cmd_3
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__46743\,
            I => comm_cmd_3
        );

    \I__11362\ : InMux
    port map (
            O => \N__46718\,
            I => \N__46715\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__46715\,
            I => \N__46712\
        );

    \I__11360\ : Span12Mux_h
    port map (
            O => \N__46712\,
            I => \N__46709\
        );

    \I__11359\ : Odrv12
    port map (
            O => \N__46709\,
            I => n4108
        );

    \I__11358\ : CascadeMux
    port map (
            O => \N__46706\,
            I => \N__46703\
        );

    \I__11357\ : InMux
    port map (
            O => \N__46703\,
            I => \N__46700\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__46700\,
            I => \N__46697\
        );

    \I__11355\ : Span4Mux_v
    port map (
            O => \N__46697\,
            I => \N__46692\
        );

    \I__11354\ : CascadeMux
    port map (
            O => \N__46696\,
            I => \N__46689\
        );

    \I__11353\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46686\
        );

    \I__11352\ : Sp12to4
    port map (
            O => \N__46692\,
            I => \N__46683\
        );

    \I__11351\ : InMux
    port map (
            O => \N__46689\,
            I => \N__46680\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__46686\,
            I => \N__46677\
        );

    \I__11349\ : Span12Mux_h
    port map (
            O => \N__46683\,
            I => \N__46674\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__46680\,
            I => cmd_rdadctmp_10_adj_1066
        );

    \I__11347\ : Odrv4
    port map (
            O => \N__46677\,
            I => cmd_rdadctmp_10_adj_1066
        );

    \I__11346\ : Odrv12
    port map (
            O => \N__46674\,
            I => cmd_rdadctmp_10_adj_1066
        );

    \I__11345\ : InMux
    port map (
            O => \N__46667\,
            I => \N__46663\
        );

    \I__11344\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46660\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__46663\,
            I => buf_adcdata2_2
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__46660\,
            I => buf_adcdata2_2
        );

    \I__11341\ : SRMux
    port map (
            O => \N__46655\,
            I => \N__46652\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__46652\,
            I => \N__46649\
        );

    \I__11339\ : Span4Mux_h
    port map (
            O => \N__46649\,
            I => \N__46646\
        );

    \I__11338\ : Span4Mux_v
    port map (
            O => \N__46646\,
            I => \N__46643\
        );

    \I__11337\ : Odrv4
    port map (
            O => \N__46643\,
            I => \comm_spi.data_tx_7__N_808\
        );

    \I__11336\ : InMux
    port map (
            O => \N__46640\,
            I => \N__46635\
        );

    \I__11335\ : InMux
    port map (
            O => \N__46639\,
            I => \N__46630\
        );

    \I__11334\ : InMux
    port map (
            O => \N__46638\,
            I => \N__46630\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__46635\,
            I => \N__46627\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__46630\,
            I => \N__46624\
        );

    \I__11331\ : Span4Mux_v
    port map (
            O => \N__46627\,
            I => \N__46621\
        );

    \I__11330\ : Span12Mux_h
    port map (
            O => \N__46624\,
            I => \N__46618\
        );

    \I__11329\ : Span4Mux_v
    port map (
            O => \N__46621\,
            I => \N__46615\
        );

    \I__11328\ : Odrv12
    port map (
            O => \N__46618\,
            I => comm_tx_buf_4
        );

    \I__11327\ : Odrv4
    port map (
            O => \N__46615\,
            I => comm_tx_buf_4
        );

    \I__11326\ : InMux
    port map (
            O => \N__46610\,
            I => \N__46588\
        );

    \I__11325\ : InMux
    port map (
            O => \N__46609\,
            I => \N__46588\
        );

    \I__11324\ : InMux
    port map (
            O => \N__46608\,
            I => \N__46588\
        );

    \I__11323\ : InMux
    port map (
            O => \N__46607\,
            I => \N__46588\
        );

    \I__11322\ : InMux
    port map (
            O => \N__46606\,
            I => \N__46588\
        );

    \I__11321\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46585\
        );

    \I__11320\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46571\
        );

    \I__11319\ : InMux
    port map (
            O => \N__46603\,
            I => \N__46562\
        );

    \I__11318\ : InMux
    port map (
            O => \N__46602\,
            I => \N__46562\
        );

    \I__11317\ : InMux
    port map (
            O => \N__46601\,
            I => \N__46562\
        );

    \I__11316\ : InMux
    port map (
            O => \N__46600\,
            I => \N__46562\
        );

    \I__11315\ : InMux
    port map (
            O => \N__46599\,
            I => \N__46557\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__46588\,
            I => \N__46550\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__46585\,
            I => \N__46550\
        );

    \I__11312\ : SRMux
    port map (
            O => \N__46584\,
            I => \N__46547\
        );

    \I__11311\ : InMux
    port map (
            O => \N__46583\,
            I => \N__46540\
        );

    \I__11310\ : InMux
    port map (
            O => \N__46582\,
            I => \N__46540\
        );

    \I__11309\ : InMux
    port map (
            O => \N__46581\,
            I => \N__46540\
        );

    \I__11308\ : SRMux
    port map (
            O => \N__46580\,
            I => \N__46537\
        );

    \I__11307\ : InMux
    port map (
            O => \N__46579\,
            I => \N__46524\
        );

    \I__11306\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46524\
        );

    \I__11305\ : InMux
    port map (
            O => \N__46577\,
            I => \N__46524\
        );

    \I__11304\ : InMux
    port map (
            O => \N__46576\,
            I => \N__46524\
        );

    \I__11303\ : InMux
    port map (
            O => \N__46575\,
            I => \N__46524\
        );

    \I__11302\ : InMux
    port map (
            O => \N__46574\,
            I => \N__46524\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__46571\,
            I => \N__46519\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__46562\,
            I => \N__46519\
        );

    \I__11299\ : InMux
    port map (
            O => \N__46561\,
            I => \N__46516\
        );

    \I__11298\ : InMux
    port map (
            O => \N__46560\,
            I => \N__46513\
        );

    \I__11297\ : LocalMux
    port map (
            O => \N__46557\,
            I => \N__46510\
        );

    \I__11296\ : InMux
    port map (
            O => \N__46556\,
            I => \N__46507\
        );

    \I__11295\ : SRMux
    port map (
            O => \N__46555\,
            I => \N__46504\
        );

    \I__11294\ : Span4Mux_v
    port map (
            O => \N__46550\,
            I => \N__46498\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__46547\,
            I => \N__46495\
        );

    \I__11292\ : LocalMux
    port map (
            O => \N__46540\,
            I => \N__46490\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__46537\,
            I => \N__46490\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__46524\,
            I => \N__46487\
        );

    \I__11289\ : Span4Mux_v
    port map (
            O => \N__46519\,
            I => \N__46484\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__46516\,
            I => \N__46481\
        );

    \I__11287\ : LocalMux
    port map (
            O => \N__46513\,
            I => \N__46478\
        );

    \I__11286\ : Span4Mux_v
    port map (
            O => \N__46510\,
            I => \N__46471\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__46507\,
            I => \N__46471\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__46504\,
            I => \N__46471\
        );

    \I__11283\ : InMux
    port map (
            O => \N__46503\,
            I => \N__46466\
        );

    \I__11282\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46457\
        );

    \I__11281\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46457\
        );

    \I__11280\ : Span4Mux_h
    port map (
            O => \N__46498\,
            I => \N__46450\
        );

    \I__11279\ : Span4Mux_v
    port map (
            O => \N__46495\,
            I => \N__46450\
        );

    \I__11278\ : Span4Mux_v
    port map (
            O => \N__46490\,
            I => \N__46450\
        );

    \I__11277\ : Span4Mux_v
    port map (
            O => \N__46487\,
            I => \N__46447\
        );

    \I__11276\ : Span4Mux_h
    port map (
            O => \N__46484\,
            I => \N__46442\
        );

    \I__11275\ : Span4Mux_v
    port map (
            O => \N__46481\,
            I => \N__46442\
        );

    \I__11274\ : Span4Mux_v
    port map (
            O => \N__46478\,
            I => \N__46437\
        );

    \I__11273\ : Span4Mux_h
    port map (
            O => \N__46471\,
            I => \N__46437\
        );

    \I__11272\ : InMux
    port map (
            O => \N__46470\,
            I => \N__46434\
        );

    \I__11271\ : InMux
    port map (
            O => \N__46469\,
            I => \N__46431\
        );

    \I__11270\ : LocalMux
    port map (
            O => \N__46466\,
            I => \N__46428\
        );

    \I__11269\ : InMux
    port map (
            O => \N__46465\,
            I => \N__46419\
        );

    \I__11268\ : InMux
    port map (
            O => \N__46464\,
            I => \N__46419\
        );

    \I__11267\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46419\
        );

    \I__11266\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46419\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__46457\,
            I => \N__46412\
        );

    \I__11264\ : Span4Mux_h
    port map (
            O => \N__46450\,
            I => \N__46412\
        );

    \I__11263\ : Span4Mux_h
    port map (
            O => \N__46447\,
            I => \N__46412\
        );

    \I__11262\ : Odrv4
    port map (
            O => \N__46442\,
            I => comm_clear
        );

    \I__11261\ : Odrv4
    port map (
            O => \N__46437\,
            I => comm_clear
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__46434\,
            I => comm_clear
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__46431\,
            I => comm_clear
        );

    \I__11258\ : Odrv4
    port map (
            O => \N__46428\,
            I => comm_clear
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__46419\,
            I => comm_clear
        );

    \I__11256\ : Odrv4
    port map (
            O => \N__46412\,
            I => comm_clear
        );

    \I__11255\ : InMux
    port map (
            O => \N__46397\,
            I => \N__46393\
        );

    \I__11254\ : InMux
    port map (
            O => \N__46396\,
            I => \N__46390\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__46393\,
            I => \N__46387\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__46390\,
            I => \N__46384\
        );

    \I__11251\ : Span4Mux_h
    port map (
            O => \N__46387\,
            I => \N__46381\
        );

    \I__11250\ : Span4Mux_h
    port map (
            O => \N__46384\,
            I => \N__46378\
        );

    \I__11249\ : Span4Mux_h
    port map (
            O => \N__46381\,
            I => \N__46374\
        );

    \I__11248\ : Span4Mux_h
    port map (
            O => \N__46378\,
            I => \N__46371\
        );

    \I__11247\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46368\
        );

    \I__11246\ : Odrv4
    port map (
            O => \N__46374\,
            I => \comm_spi.n16899\
        );

    \I__11245\ : Odrv4
    port map (
            O => \N__46371\,
            I => \comm_spi.n16899\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__46368\,
            I => \comm_spi.n16899\
        );

    \I__11243\ : CascadeMux
    port map (
            O => \N__46361\,
            I => \N__46358\
        );

    \I__11242\ : InMux
    port map (
            O => \N__46358\,
            I => \N__46354\
        );

    \I__11241\ : CascadeMux
    port map (
            O => \N__46357\,
            I => \N__46350\
        );

    \I__11240\ : LocalMux
    port map (
            O => \N__46354\,
            I => \N__46347\
        );

    \I__11239\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46344\
        );

    \I__11238\ : InMux
    port map (
            O => \N__46350\,
            I => \N__46341\
        );

    \I__11237\ : Span4Mux_v
    port map (
            O => \N__46347\,
            I => \N__46338\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__46344\,
            I => cmd_rdadctmp_29_adj_1047
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__46341\,
            I => cmd_rdadctmp_29_adj_1047
        );

    \I__11234\ : Odrv4
    port map (
            O => \N__46338\,
            I => cmd_rdadctmp_29_adj_1047
        );

    \I__11233\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46328\
        );

    \I__11232\ : LocalMux
    port map (
            O => \N__46328\,
            I => \N__46324\
        );

    \I__11231\ : InMux
    port map (
            O => \N__46327\,
            I => \N__46321\
        );

    \I__11230\ : Span4Mux_v
    port map (
            O => \N__46324\,
            I => \N__46318\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__46321\,
            I => buf_adcdata2_21
        );

    \I__11228\ : Odrv4
    port map (
            O => \N__46318\,
            I => buf_adcdata2_21
        );

    \I__11227\ : IoInMux
    port map (
            O => \N__46313\,
            I => \N__46310\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__46310\,
            I => \N__46307\
        );

    \I__11225\ : IoSpan4Mux
    port map (
            O => \N__46307\,
            I => \N__46304\
        );

    \I__11224\ : IoSpan4Mux
    port map (
            O => \N__46304\,
            I => \N__46301\
        );

    \I__11223\ : Span4Mux_s3_h
    port map (
            O => \N__46301\,
            I => \N__46298\
        );

    \I__11222\ : Span4Mux_h
    port map (
            O => \N__46298\,
            I => \N__46295\
        );

    \I__11221\ : Odrv4
    port map (
            O => \N__46295\,
            I => \ICE_GPMI_0\
        );

    \I__11220\ : CascadeMux
    port map (
            O => \N__46292\,
            I => \N__46289\
        );

    \I__11219\ : InMux
    port map (
            O => \N__46289\,
            I => \N__46286\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__46286\,
            I => \N__46282\
        );

    \I__11217\ : CascadeMux
    port map (
            O => \N__46285\,
            I => \N__46279\
        );

    \I__11216\ : Span4Mux_v
    port map (
            O => \N__46282\,
            I => \N__46276\
        );

    \I__11215\ : InMux
    port map (
            O => \N__46279\,
            I => \N__46273\
        );

    \I__11214\ : Span4Mux_h
    port map (
            O => \N__46276\,
            I => \N__46269\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__46273\,
            I => \N__46266\
        );

    \I__11212\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46263\
        );

    \I__11211\ : Odrv4
    port map (
            O => \N__46269\,
            I => cmd_rdadctmp_20
        );

    \I__11210\ : Odrv4
    port map (
            O => \N__46266\,
            I => cmd_rdadctmp_20
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__46263\,
            I => cmd_rdadctmp_20
        );

    \I__11208\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46253\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__46253\,
            I => \N__46249\
        );

    \I__11206\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46246\
        );

    \I__11205\ : Span4Mux_h
    port map (
            O => \N__46249\,
            I => \N__46243\
        );

    \I__11204\ : LocalMux
    port map (
            O => \N__46246\,
            I => buf_adcdata1_12
        );

    \I__11203\ : Odrv4
    port map (
            O => \N__46243\,
            I => buf_adcdata1_12
        );

    \I__11202\ : CascadeMux
    port map (
            O => \N__46238\,
            I => \N__46235\
        );

    \I__11201\ : InMux
    port map (
            O => \N__46235\,
            I => \N__46232\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__46232\,
            I => \N__46229\
        );

    \I__11199\ : Span12Mux_s11_v
    port map (
            O => \N__46229\,
            I => \N__46224\
        );

    \I__11198\ : InMux
    port map (
            O => \N__46228\,
            I => \N__46221\
        );

    \I__11197\ : CascadeMux
    port map (
            O => \N__46227\,
            I => \N__46218\
        );

    \I__11196\ : Span12Mux_h
    port map (
            O => \N__46224\,
            I => \N__46215\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__46221\,
            I => \N__46212\
        );

    \I__11194\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46209\
        );

    \I__11193\ : Odrv12
    port map (
            O => \N__46215\,
            I => cmd_rdadctmp_17_adj_1059
        );

    \I__11192\ : Odrv12
    port map (
            O => \N__46212\,
            I => cmd_rdadctmp_17_adj_1059
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__46209\,
            I => cmd_rdadctmp_17_adj_1059
        );

    \I__11190\ : InMux
    port map (
            O => \N__46202\,
            I => \N__46199\
        );

    \I__11189\ : LocalMux
    port map (
            O => \N__46199\,
            I => \N__46196\
        );

    \I__11188\ : Span4Mux_v
    port map (
            O => \N__46196\,
            I => \N__46192\
        );

    \I__11187\ : InMux
    port map (
            O => \N__46195\,
            I => \N__46189\
        );

    \I__11186\ : Span4Mux_h
    port map (
            O => \N__46192\,
            I => \N__46186\
        );

    \I__11185\ : LocalMux
    port map (
            O => \N__46189\,
            I => buf_adcdata2_9
        );

    \I__11184\ : Odrv4
    port map (
            O => \N__46186\,
            I => buf_adcdata2_9
        );

    \I__11183\ : CascadeMux
    port map (
            O => \N__46181\,
            I => \N__46178\
        );

    \I__11182\ : InMux
    port map (
            O => \N__46178\,
            I => \N__46174\
        );

    \I__11181\ : InMux
    port map (
            O => \N__46177\,
            I => \N__46171\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__46174\,
            I => \N__46168\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__46171\,
            I => \N__46165\
        );

    \I__11178\ : Span4Mux_v
    port map (
            O => \N__46168\,
            I => \N__46159\
        );

    \I__11177\ : Span4Mux_h
    port map (
            O => \N__46165\,
            I => \N__46159\
        );

    \I__11176\ : CascadeMux
    port map (
            O => \N__46164\,
            I => \N__46156\
        );

    \I__11175\ : Span4Mux_h
    port map (
            O => \N__46159\,
            I => \N__46153\
        );

    \I__11174\ : InMux
    port map (
            O => \N__46156\,
            I => \N__46150\
        );

    \I__11173\ : Odrv4
    port map (
            O => \N__46153\,
            I => cmd_rdadctmp_19_adj_1057
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__46150\,
            I => cmd_rdadctmp_19_adj_1057
        );

    \I__11171\ : CascadeMux
    port map (
            O => \N__46145\,
            I => \N__46142\
        );

    \I__11170\ : InMux
    port map (
            O => \N__46142\,
            I => \N__46138\
        );

    \I__11169\ : CascadeMux
    port map (
            O => \N__46141\,
            I => \N__46134\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__46138\,
            I => \N__46131\
        );

    \I__11167\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46126\
        );

    \I__11166\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46126\
        );

    \I__11165\ : Odrv4
    port map (
            O => \N__46131\,
            I => cmd_rdadctmp_20_adj_1056
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__46126\,
            I => cmd_rdadctmp_20_adj_1056
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__46121\,
            I => \N__46112\
        );

    \I__11162\ : CascadeMux
    port map (
            O => \N__46120\,
            I => \N__46109\
        );

    \I__11161\ : InMux
    port map (
            O => \N__46119\,
            I => \N__46097\
        );

    \I__11160\ : InMux
    port map (
            O => \N__46118\,
            I => \N__46097\
        );

    \I__11159\ : InMux
    port map (
            O => \N__46117\,
            I => \N__46097\
        );

    \I__11158\ : InMux
    port map (
            O => \N__46116\,
            I => \N__46097\
        );

    \I__11157\ : InMux
    port map (
            O => \N__46115\,
            I => \N__46097\
        );

    \I__11156\ : InMux
    port map (
            O => \N__46112\,
            I => \N__46090\
        );

    \I__11155\ : InMux
    port map (
            O => \N__46109\,
            I => \N__46090\
        );

    \I__11154\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46090\
        );

    \I__11153\ : LocalMux
    port map (
            O => \N__46097\,
            I => \N__46086\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__46090\,
            I => \N__46083\
        );

    \I__11151\ : InMux
    port map (
            O => \N__46089\,
            I => \N__46073\
        );

    \I__11150\ : Span4Mux_v
    port map (
            O => \N__46086\,
            I => \N__46067\
        );

    \I__11149\ : Span4Mux_v
    port map (
            O => \N__46083\,
            I => \N__46067\
        );

    \I__11148\ : InMux
    port map (
            O => \N__46082\,
            I => \N__46064\
        );

    \I__11147\ : InMux
    port map (
            O => \N__46081\,
            I => \N__46059\
        );

    \I__11146\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46053\
        );

    \I__11145\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46053\
        );

    \I__11144\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46046\
        );

    \I__11143\ : InMux
    port map (
            O => \N__46077\,
            I => \N__46046\
        );

    \I__11142\ : InMux
    port map (
            O => \N__46076\,
            I => \N__46046\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__46073\,
            I => \N__46043\
        );

    \I__11140\ : InMux
    port map (
            O => \N__46072\,
            I => \N__46040\
        );

    \I__11139\ : Span4Mux_h
    port map (
            O => \N__46067\,
            I => \N__46034\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__46064\,
            I => \N__46031\
        );

    \I__11137\ : InMux
    port map (
            O => \N__46063\,
            I => \N__46028\
        );

    \I__11136\ : InMux
    port map (
            O => \N__46062\,
            I => \N__46025\
        );

    \I__11135\ : LocalMux
    port map (
            O => \N__46059\,
            I => \N__46022\
        );

    \I__11134\ : InMux
    port map (
            O => \N__46058\,
            I => \N__46019\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__46053\,
            I => \N__46014\
        );

    \I__11132\ : LocalMux
    port map (
            O => \N__46046\,
            I => \N__46014\
        );

    \I__11131\ : Span4Mux_v
    port map (
            O => \N__46043\,
            I => \N__46011\
        );

    \I__11130\ : LocalMux
    port map (
            O => \N__46040\,
            I => \N__46008\
        );

    \I__11129\ : InMux
    port map (
            O => \N__46039\,
            I => \N__46005\
        );

    \I__11128\ : CascadeMux
    port map (
            O => \N__46038\,
            I => \N__45998\
        );

    \I__11127\ : CascadeMux
    port map (
            O => \N__46037\,
            I => \N__45994\
        );

    \I__11126\ : Sp12to4
    port map (
            O => \N__46034\,
            I => \N__45986\
        );

    \I__11125\ : Span12Mux_v
    port map (
            O => \N__46031\,
            I => \N__45986\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__46028\,
            I => \N__45986\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__46025\,
            I => \N__45983\
        );

    \I__11122\ : Span4Mux_h
    port map (
            O => \N__46022\,
            I => \N__45978\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__46019\,
            I => \N__45978\
        );

    \I__11120\ : Span4Mux_v
    port map (
            O => \N__46014\,
            I => \N__45975\
        );

    \I__11119\ : Span4Mux_h
    port map (
            O => \N__46011\,
            I => \N__45968\
        );

    \I__11118\ : Span4Mux_v
    port map (
            O => \N__46008\,
            I => \N__45968\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__46005\,
            I => \N__45968\
        );

    \I__11116\ : InMux
    port map (
            O => \N__46004\,
            I => \N__45959\
        );

    \I__11115\ : InMux
    port map (
            O => \N__46003\,
            I => \N__45959\
        );

    \I__11114\ : InMux
    port map (
            O => \N__46002\,
            I => \N__45959\
        );

    \I__11113\ : InMux
    port map (
            O => \N__46001\,
            I => \N__45959\
        );

    \I__11112\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45950\
        );

    \I__11111\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45950\
        );

    \I__11110\ : InMux
    port map (
            O => \N__45994\,
            I => \N__45950\
        );

    \I__11109\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45950\
        );

    \I__11108\ : Span12Mux_h
    port map (
            O => \N__45986\,
            I => \N__45945\
        );

    \I__11107\ : Span4Mux_v
    port map (
            O => \N__45983\,
            I => \N__45942\
        );

    \I__11106\ : Span4Mux_h
    port map (
            O => \N__45978\,
            I => \N__45939\
        );

    \I__11105\ : Span4Mux_v
    port map (
            O => \N__45975\,
            I => \N__45934\
        );

    \I__11104\ : Span4Mux_h
    port map (
            O => \N__45968\,
            I => \N__45934\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__45959\,
            I => \N__45931\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__45950\,
            I => \N__45928\
        );

    \I__11101\ : InMux
    port map (
            O => \N__45949\,
            I => \N__45923\
        );

    \I__11100\ : InMux
    port map (
            O => \N__45948\,
            I => \N__45923\
        );

    \I__11099\ : Odrv12
    port map (
            O => \N__45945\,
            I => n8302
        );

    \I__11098\ : Odrv4
    port map (
            O => \N__45942\,
            I => n8302
        );

    \I__11097\ : Odrv4
    port map (
            O => \N__45939\,
            I => n8302
        );

    \I__11096\ : Odrv4
    port map (
            O => \N__45934\,
            I => n8302
        );

    \I__11095\ : Odrv12
    port map (
            O => \N__45931\,
            I => n8302
        );

    \I__11094\ : Odrv4
    port map (
            O => \N__45928\,
            I => n8302
        );

    \I__11093\ : LocalMux
    port map (
            O => \N__45923\,
            I => n8302
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__45908\,
            I => \N__45905\
        );

    \I__11091\ : InMux
    port map (
            O => \N__45905\,
            I => \N__45900\
        );

    \I__11090\ : InMux
    port map (
            O => \N__45904\,
            I => \N__45895\
        );

    \I__11089\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45895\
        );

    \I__11088\ : LocalMux
    port map (
            O => \N__45900\,
            I => cmd_rdadctmp_21_adj_1055
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__45895\,
            I => cmd_rdadctmp_21_adj_1055
        );

    \I__11086\ : InMux
    port map (
            O => \N__45890\,
            I => \N__45887\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__45887\,
            I => \N__45884\
        );

    \I__11084\ : Span4Mux_h
    port map (
            O => \N__45884\,
            I => \N__45881\
        );

    \I__11083\ : Odrv4
    port map (
            O => \N__45881\,
            I => buf_data2_23
        );

    \I__11082\ : InMux
    port map (
            O => \N__45878\,
            I => \N__45874\
        );

    \I__11081\ : CascadeMux
    port map (
            O => \N__45877\,
            I => \N__45871\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__45874\,
            I => \N__45868\
        );

    \I__11079\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45864\
        );

    \I__11078\ : Span4Mux_h
    port map (
            O => \N__45868\,
            I => \N__45861\
        );

    \I__11077\ : CascadeMux
    port map (
            O => \N__45867\,
            I => \N__45858\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__45864\,
            I => \N__45855\
        );

    \I__11075\ : Span4Mux_v
    port map (
            O => \N__45861\,
            I => \N__45852\
        );

    \I__11074\ : InMux
    port map (
            O => \N__45858\,
            I => \N__45849\
        );

    \I__11073\ : Span12Mux_s10_v
    port map (
            O => \N__45855\,
            I => \N__45846\
        );

    \I__11072\ : Span4Mux_h
    port map (
            O => \N__45852\,
            I => \N__45843\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__45849\,
            I => buf_adcdata4_23
        );

    \I__11070\ : Odrv12
    port map (
            O => \N__45846\,
            I => buf_adcdata4_23
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__45843\,
            I => buf_adcdata4_23
        );

    \I__11068\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45833\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__45833\,
            I => \N__45830\
        );

    \I__11066\ : Span4Mux_v
    port map (
            O => \N__45830\,
            I => \N__45827\
        );

    \I__11065\ : Span4Mux_h
    port map (
            O => \N__45827\,
            I => \N__45824\
        );

    \I__11064\ : Sp12to4
    port map (
            O => \N__45824\,
            I => \N__45821\
        );

    \I__11063\ : Odrv12
    port map (
            O => \N__45821\,
            I => n4101
        );

    \I__11062\ : InMux
    port map (
            O => \N__45818\,
            I => \N__45815\
        );

    \I__11061\ : LocalMux
    port map (
            O => \N__45815\,
            I => \N__45810\
        );

    \I__11060\ : InMux
    port map (
            O => \N__45814\,
            I => \N__45807\
        );

    \I__11059\ : InMux
    port map (
            O => \N__45813\,
            I => \N__45804\
        );

    \I__11058\ : Odrv12
    port map (
            O => \N__45810\,
            I => \comm_spi.n10442\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__45807\,
            I => \comm_spi.n10442\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__45804\,
            I => \comm_spi.n10442\
        );

    \I__11055\ : InMux
    port map (
            O => \N__45797\,
            I => \N__45789\
        );

    \I__11054\ : InMux
    port map (
            O => \N__45796\,
            I => \N__45789\
        );

    \I__11053\ : InMux
    port map (
            O => \N__45795\,
            I => \N__45786\
        );

    \I__11052\ : InMux
    port map (
            O => \N__45794\,
            I => \N__45783\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__45789\,
            I => \N__45778\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__45786\,
            I => \N__45778\
        );

    \I__11049\ : LocalMux
    port map (
            O => \N__45783\,
            I => \N__45774\
        );

    \I__11048\ : Span4Mux_v
    port map (
            O => \N__45778\,
            I => \N__45771\
        );

    \I__11047\ : InMux
    port map (
            O => \N__45777\,
            I => \N__45768\
        );

    \I__11046\ : Span4Mux_v
    port map (
            O => \N__45774\,
            I => \N__45765\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__45771\,
            I => \N__45762\
        );

    \I__11044\ : LocalMux
    port map (
            O => \N__45768\,
            I => \N__45759\
        );

    \I__11043\ : Sp12to4
    port map (
            O => \N__45765\,
            I => \N__45754\
        );

    \I__11042\ : Sp12to4
    port map (
            O => \N__45762\,
            I => \N__45754\
        );

    \I__11041\ : Span4Mux_h
    port map (
            O => \N__45759\,
            I => \N__45751\
        );

    \I__11040\ : Span12Mux_s6_h
    port map (
            O => \N__45754\,
            I => \N__45746\
        );

    \I__11039\ : Sp12to4
    port map (
            O => \N__45751\,
            I => \N__45746\
        );

    \I__11038\ : Span12Mux_v
    port map (
            O => \N__45746\,
            I => \N__45743\
        );

    \I__11037\ : Odrv12
    port map (
            O => \N__45743\,
            I => \ICE_SPI_MOSI\
        );

    \I__11036\ : SRMux
    port map (
            O => \N__45740\,
            I => \N__45737\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__45737\,
            I => \comm_spi.imosi_N_792\
        );

    \I__11034\ : CascadeMux
    port map (
            O => \N__45734\,
            I => \N__45731\
        );

    \I__11033\ : InMux
    port map (
            O => \N__45731\,
            I => \N__45727\
        );

    \I__11032\ : CascadeMux
    port map (
            O => \N__45730\,
            I => \N__45723\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__45727\,
            I => \N__45720\
        );

    \I__11030\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45715\
        );

    \I__11029\ : InMux
    port map (
            O => \N__45723\,
            I => \N__45715\
        );

    \I__11028\ : Span4Mux_v
    port map (
            O => \N__45720\,
            I => \N__45712\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__45715\,
            I => cmd_rdadctmp_28_adj_1048
        );

    \I__11026\ : Odrv4
    port map (
            O => \N__45712\,
            I => cmd_rdadctmp_28_adj_1048
        );

    \I__11025\ : InMux
    port map (
            O => \N__45707\,
            I => \N__45704\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__45704\,
            I => \N__45700\
        );

    \I__11023\ : InMux
    port map (
            O => \N__45703\,
            I => \N__45697\
        );

    \I__11022\ : Span4Mux_h
    port map (
            O => \N__45700\,
            I => \N__45694\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__45697\,
            I => buf_adcdata2_20
        );

    \I__11020\ : Odrv4
    port map (
            O => \N__45694\,
            I => buf_adcdata2_20
        );

    \I__11019\ : InMux
    port map (
            O => \N__45689\,
            I => \N__45686\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__45686\,
            I => \N__45683\
        );

    \I__11017\ : Odrv12
    port map (
            O => \N__45683\,
            I => n4_adj_1250
        );

    \I__11016\ : InMux
    port map (
            O => \N__45680\,
            I => \N__45677\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__45677\,
            I => \N__45673\
        );

    \I__11014\ : InMux
    port map (
            O => \N__45676\,
            I => \N__45670\
        );

    \I__11013\ : Span4Mux_h
    port map (
            O => \N__45673\,
            I => \N__45667\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__45670\,
            I => buf_adcdata2_12
        );

    \I__11011\ : Odrv4
    port map (
            O => \N__45667\,
            I => buf_adcdata2_12
        );

    \I__11010\ : InMux
    port map (
            O => \N__45662\,
            I => \N__45640\
        );

    \I__11009\ : InMux
    port map (
            O => \N__45661\,
            I => \N__45640\
        );

    \I__11008\ : InMux
    port map (
            O => \N__45660\,
            I => \N__45636\
        );

    \I__11007\ : InMux
    port map (
            O => \N__45659\,
            I => \N__45633\
        );

    \I__11006\ : InMux
    port map (
            O => \N__45658\,
            I => \N__45630\
        );

    \I__11005\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45627\
        );

    \I__11004\ : InMux
    port map (
            O => \N__45656\,
            I => \N__45622\
        );

    \I__11003\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45622\
        );

    \I__11002\ : InMux
    port map (
            O => \N__45654\,
            I => \N__45619\
        );

    \I__11001\ : CascadeMux
    port map (
            O => \N__45653\,
            I => \N__45616\
        );

    \I__11000\ : InMux
    port map (
            O => \N__45652\,
            I => \N__45613\
        );

    \I__10999\ : InMux
    port map (
            O => \N__45651\,
            I => \N__45608\
        );

    \I__10998\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45608\
        );

    \I__10997\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45599\
        );

    \I__10996\ : InMux
    port map (
            O => \N__45648\,
            I => \N__45592\
        );

    \I__10995\ : InMux
    port map (
            O => \N__45647\,
            I => \N__45592\
        );

    \I__10994\ : InMux
    port map (
            O => \N__45646\,
            I => \N__45589\
        );

    \I__10993\ : InMux
    port map (
            O => \N__45645\,
            I => \N__45586\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45583\
        );

    \I__10991\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45580\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__45636\,
            I => \N__45575\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__45633\,
            I => \N__45575\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__45630\,
            I => \N__45572\
        );

    \I__10987\ : LocalMux
    port map (
            O => \N__45627\,
            I => \N__45569\
        );

    \I__10986\ : LocalMux
    port map (
            O => \N__45622\,
            I => \N__45566\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__45619\,
            I => \N__45563\
        );

    \I__10984\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45560\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__45613\,
            I => \N__45557\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__45608\,
            I => \N__45554\
        );

    \I__10981\ : InMux
    port map (
            O => \N__45607\,
            I => \N__45551\
        );

    \I__10980\ : InMux
    port map (
            O => \N__45606\,
            I => \N__45546\
        );

    \I__10979\ : InMux
    port map (
            O => \N__45605\,
            I => \N__45546\
        );

    \I__10978\ : InMux
    port map (
            O => \N__45604\,
            I => \N__45531\
        );

    \I__10977\ : InMux
    port map (
            O => \N__45603\,
            I => \N__45531\
        );

    \I__10976\ : InMux
    port map (
            O => \N__45602\,
            I => \N__45528\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__45599\,
            I => \N__45525\
        );

    \I__10974\ : InMux
    port map (
            O => \N__45598\,
            I => \N__45522\
        );

    \I__10973\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45519\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__45592\,
            I => \N__45506\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__45589\,
            I => \N__45506\
        );

    \I__10970\ : LocalMux
    port map (
            O => \N__45586\,
            I => \N__45506\
        );

    \I__10969\ : Span4Mux_v
    port map (
            O => \N__45583\,
            I => \N__45506\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__45580\,
            I => \N__45506\
        );

    \I__10967\ : Span4Mux_h
    port map (
            O => \N__45575\,
            I => \N__45506\
        );

    \I__10966\ : Span4Mux_v
    port map (
            O => \N__45572\,
            I => \N__45501\
        );

    \I__10965\ : Span4Mux_v
    port map (
            O => \N__45569\,
            I => \N__45501\
        );

    \I__10964\ : Span4Mux_h
    port map (
            O => \N__45566\,
            I => \N__45497\
        );

    \I__10963\ : Span4Mux_h
    port map (
            O => \N__45563\,
            I => \N__45488\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__45560\,
            I => \N__45488\
        );

    \I__10961\ : Span4Mux_v
    port map (
            O => \N__45557\,
            I => \N__45488\
        );

    \I__10960\ : Span4Mux_v
    port map (
            O => \N__45554\,
            I => \N__45488\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__45551\,
            I => \N__45483\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__45546\,
            I => \N__45483\
        );

    \I__10957\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45478\
        );

    \I__10956\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45478\
        );

    \I__10955\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45471\
        );

    \I__10954\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45471\
        );

    \I__10953\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45471\
        );

    \I__10952\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45466\
        );

    \I__10951\ : InMux
    port map (
            O => \N__45539\,
            I => \N__45466\
        );

    \I__10950\ : InMux
    port map (
            O => \N__45538\,
            I => \N__45461\
        );

    \I__10949\ : InMux
    port map (
            O => \N__45537\,
            I => \N__45456\
        );

    \I__10948\ : InMux
    port map (
            O => \N__45536\,
            I => \N__45456\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__45531\,
            I => \N__45451\
        );

    \I__10946\ : LocalMux
    port map (
            O => \N__45528\,
            I => \N__45446\
        );

    \I__10945\ : Span4Mux_h
    port map (
            O => \N__45525\,
            I => \N__45446\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__45522\,
            I => \N__45441\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__45519\,
            I => \N__45441\
        );

    \I__10942\ : Span4Mux_h
    port map (
            O => \N__45506\,
            I => \N__45438\
        );

    \I__10941\ : Span4Mux_h
    port map (
            O => \N__45501\,
            I => \N__45432\
        );

    \I__10940\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45429\
        );

    \I__10939\ : Span4Mux_h
    port map (
            O => \N__45497\,
            I => \N__45416\
        );

    \I__10938\ : Span4Mux_h
    port map (
            O => \N__45488\,
            I => \N__45416\
        );

    \I__10937\ : Span4Mux_v
    port map (
            O => \N__45483\,
            I => \N__45416\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__45478\,
            I => \N__45416\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45416\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45416\
        );

    \I__10933\ : CascadeMux
    port map (
            O => \N__45465\,
            I => \N__45406\
        );

    \I__10932\ : InMux
    port map (
            O => \N__45464\,
            I => \N__45402\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__45461\,
            I => \N__45397\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__45456\,
            I => \N__45397\
        );

    \I__10929\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45394\
        );

    \I__10928\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45391\
        );

    \I__10927\ : Span4Mux_h
    port map (
            O => \N__45451\,
            I => \N__45382\
        );

    \I__10926\ : Span4Mux_v
    port map (
            O => \N__45446\,
            I => \N__45382\
        );

    \I__10925\ : Span4Mux_h
    port map (
            O => \N__45441\,
            I => \N__45382\
        );

    \I__10924\ : Span4Mux_h
    port map (
            O => \N__45438\,
            I => \N__45382\
        );

    \I__10923\ : InMux
    port map (
            O => \N__45437\,
            I => \N__45379\
        );

    \I__10922\ : InMux
    port map (
            O => \N__45436\,
            I => \N__45374\
        );

    \I__10921\ : InMux
    port map (
            O => \N__45435\,
            I => \N__45374\
        );

    \I__10920\ : Span4Mux_h
    port map (
            O => \N__45432\,
            I => \N__45369\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__45429\,
            I => \N__45369\
        );

    \I__10918\ : Span4Mux_v
    port map (
            O => \N__45416\,
            I => \N__45366\
        );

    \I__10917\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45361\
        );

    \I__10916\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45361\
        );

    \I__10915\ : InMux
    port map (
            O => \N__45413\,
            I => \N__45352\
        );

    \I__10914\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45352\
        );

    \I__10913\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45352\
        );

    \I__10912\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45352\
        );

    \I__10911\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45349\
        );

    \I__10910\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45344\
        );

    \I__10909\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45344\
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__45402\,
            I => comm_cmd_2
        );

    \I__10907\ : Odrv12
    port map (
            O => \N__45397\,
            I => comm_cmd_2
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__45394\,
            I => comm_cmd_2
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__45391\,
            I => comm_cmd_2
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__45382\,
            I => comm_cmd_2
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__45379\,
            I => comm_cmd_2
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__45374\,
            I => comm_cmd_2
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__45369\,
            I => comm_cmd_2
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__45366\,
            I => comm_cmd_2
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__45361\,
            I => comm_cmd_2
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__45352\,
            I => comm_cmd_2
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__45349\,
            I => comm_cmd_2
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__45344\,
            I => comm_cmd_2
        );

    \I__10895\ : CascadeMux
    port map (
            O => \N__45317\,
            I => \N__45314\
        );

    \I__10894\ : InMux
    port map (
            O => \N__45314\,
            I => \N__45310\
        );

    \I__10893\ : CascadeMux
    port map (
            O => \N__45313\,
            I => \N__45303\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__45310\,
            I => \N__45299\
        );

    \I__10891\ : InMux
    port map (
            O => \N__45309\,
            I => \N__45290\
        );

    \I__10890\ : InMux
    port map (
            O => \N__45308\,
            I => \N__45286\
        );

    \I__10889\ : InMux
    port map (
            O => \N__45307\,
            I => \N__45280\
        );

    \I__10888\ : InMux
    port map (
            O => \N__45306\,
            I => \N__45280\
        );

    \I__10887\ : InMux
    port map (
            O => \N__45303\,
            I => \N__45273\
        );

    \I__10886\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45273\
        );

    \I__10885\ : Span4Mux_v
    port map (
            O => \N__45299\,
            I => \N__45270\
        );

    \I__10884\ : InMux
    port map (
            O => \N__45298\,
            I => \N__45265\
        );

    \I__10883\ : InMux
    port map (
            O => \N__45297\,
            I => \N__45265\
        );

    \I__10882\ : InMux
    port map (
            O => \N__45296\,
            I => \N__45256\
        );

    \I__10881\ : InMux
    port map (
            O => \N__45295\,
            I => \N__45256\
        );

    \I__10880\ : InMux
    port map (
            O => \N__45294\,
            I => \N__45253\
        );

    \I__10879\ : InMux
    port map (
            O => \N__45293\,
            I => \N__45250\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__45290\,
            I => \N__45247\
        );

    \I__10877\ : InMux
    port map (
            O => \N__45289\,
            I => \N__45244\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__45286\,
            I => \N__45241\
        );

    \I__10875\ : InMux
    port map (
            O => \N__45285\,
            I => \N__45226\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__45280\,
            I => \N__45212\
        );

    \I__10873\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45207\
        );

    \I__10872\ : InMux
    port map (
            O => \N__45278\,
            I => \N__45207\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__45273\,
            I => \N__45200\
        );

    \I__10870\ : Span4Mux_h
    port map (
            O => \N__45270\,
            I => \N__45200\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__45265\,
            I => \N__45200\
        );

    \I__10868\ : InMux
    port map (
            O => \N__45264\,
            I => \N__45197\
        );

    \I__10867\ : InMux
    port map (
            O => \N__45263\,
            I => \N__45190\
        );

    \I__10866\ : InMux
    port map (
            O => \N__45262\,
            I => \N__45190\
        );

    \I__10865\ : InMux
    port map (
            O => \N__45261\,
            I => \N__45190\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__45256\,
            I => \N__45185\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__45253\,
            I => \N__45185\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__45250\,
            I => \N__45173\
        );

    \I__10861\ : Span4Mux_h
    port map (
            O => \N__45247\,
            I => \N__45173\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__45244\,
            I => \N__45173\
        );

    \I__10859\ : Span4Mux_v
    port map (
            O => \N__45241\,
            I => \N__45173\
        );

    \I__10858\ : InMux
    port map (
            O => \N__45240\,
            I => \N__45170\
        );

    \I__10857\ : InMux
    port map (
            O => \N__45239\,
            I => \N__45167\
        );

    \I__10856\ : InMux
    port map (
            O => \N__45238\,
            I => \N__45160\
        );

    \I__10855\ : InMux
    port map (
            O => \N__45237\,
            I => \N__45160\
        );

    \I__10854\ : InMux
    port map (
            O => \N__45236\,
            I => \N__45160\
        );

    \I__10853\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45155\
        );

    \I__10852\ : InMux
    port map (
            O => \N__45234\,
            I => \N__45155\
        );

    \I__10851\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45142\
        );

    \I__10850\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45142\
        );

    \I__10849\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45142\
        );

    \I__10848\ : InMux
    port map (
            O => \N__45230\,
            I => \N__45142\
        );

    \I__10847\ : InMux
    port map (
            O => \N__45229\,
            I => \N__45139\
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__45226\,
            I => \N__45136\
        );

    \I__10845\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45133\
        );

    \I__10844\ : InMux
    port map (
            O => \N__45224\,
            I => \N__45128\
        );

    \I__10843\ : InMux
    port map (
            O => \N__45223\,
            I => \N__45128\
        );

    \I__10842\ : InMux
    port map (
            O => \N__45222\,
            I => \N__45123\
        );

    \I__10841\ : InMux
    port map (
            O => \N__45221\,
            I => \N__45123\
        );

    \I__10840\ : InMux
    port map (
            O => \N__45220\,
            I => \N__45120\
        );

    \I__10839\ : InMux
    port map (
            O => \N__45219\,
            I => \N__45117\
        );

    \I__10838\ : InMux
    port map (
            O => \N__45218\,
            I => \N__45114\
        );

    \I__10837\ : InMux
    port map (
            O => \N__45217\,
            I => \N__45109\
        );

    \I__10836\ : InMux
    port map (
            O => \N__45216\,
            I => \N__45109\
        );

    \I__10835\ : CascadeMux
    port map (
            O => \N__45215\,
            I => \N__45106\
        );

    \I__10834\ : Span4Mux_h
    port map (
            O => \N__45212\,
            I => \N__45096\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__45207\,
            I => \N__45096\
        );

    \I__10832\ : Span4Mux_h
    port map (
            O => \N__45200\,
            I => \N__45096\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__45197\,
            I => \N__45096\
        );

    \I__10830\ : LocalMux
    port map (
            O => \N__45190\,
            I => \N__45091\
        );

    \I__10829\ : Span4Mux_h
    port map (
            O => \N__45185\,
            I => \N__45091\
        );

    \I__10828\ : InMux
    port map (
            O => \N__45184\,
            I => \N__45084\
        );

    \I__10827\ : InMux
    port map (
            O => \N__45183\,
            I => \N__45084\
        );

    \I__10826\ : InMux
    port map (
            O => \N__45182\,
            I => \N__45084\
        );

    \I__10825\ : Span4Mux_h
    port map (
            O => \N__45173\,
            I => \N__45079\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__45170\,
            I => \N__45079\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__45167\,
            I => \N__45076\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__45160\,
            I => \N__45071\
        );

    \I__10821\ : LocalMux
    port map (
            O => \N__45155\,
            I => \N__45071\
        );

    \I__10820\ : InMux
    port map (
            O => \N__45154\,
            I => \N__45066\
        );

    \I__10819\ : InMux
    port map (
            O => \N__45153\,
            I => \N__45066\
        );

    \I__10818\ : InMux
    port map (
            O => \N__45152\,
            I => \N__45063\
        );

    \I__10817\ : InMux
    port map (
            O => \N__45151\,
            I => \N__45060\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__45142\,
            I => \N__45055\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__45139\,
            I => \N__45044\
        );

    \I__10814\ : Span4Mux_v
    port map (
            O => \N__45136\,
            I => \N__45044\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__45133\,
            I => \N__45044\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__45128\,
            I => \N__45044\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__45123\,
            I => \N__45044\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__45120\,
            I => \N__45031\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__45117\,
            I => \N__45031\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__45114\,
            I => \N__45031\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__45109\,
            I => \N__45031\
        );

    \I__10806\ : InMux
    port map (
            O => \N__45106\,
            I => \N__45026\
        );

    \I__10805\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45026\
        );

    \I__10804\ : Span4Mux_v
    port map (
            O => \N__45096\,
            I => \N__45019\
        );

    \I__10803\ : Span4Mux_v
    port map (
            O => \N__45091\,
            I => \N__45019\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__45084\,
            I => \N__45019\
        );

    \I__10801\ : Span4Mux_h
    port map (
            O => \N__45079\,
            I => \N__45006\
        );

    \I__10800\ : Span4Mux_h
    port map (
            O => \N__45076\,
            I => \N__45006\
        );

    \I__10799\ : Span4Mux_v
    port map (
            O => \N__45071\,
            I => \N__45006\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__45066\,
            I => \N__45006\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__45063\,
            I => \N__45006\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__45060\,
            I => \N__45006\
        );

    \I__10795\ : InMux
    port map (
            O => \N__45059\,
            I => \N__45001\
        );

    \I__10794\ : InMux
    port map (
            O => \N__45058\,
            I => \N__45001\
        );

    \I__10793\ : Span4Mux_h
    port map (
            O => \N__45055\,
            I => \N__44996\
        );

    \I__10792\ : Span4Mux_h
    port map (
            O => \N__45044\,
            I => \N__44996\
        );

    \I__10791\ : InMux
    port map (
            O => \N__45043\,
            I => \N__44991\
        );

    \I__10790\ : InMux
    port map (
            O => \N__45042\,
            I => \N__44991\
        );

    \I__10789\ : InMux
    port map (
            O => \N__45041\,
            I => \N__44986\
        );

    \I__10788\ : InMux
    port map (
            O => \N__45040\,
            I => \N__44986\
        );

    \I__10787\ : Odrv12
    port map (
            O => \N__45031\,
            I => comm_cmd_1
        );

    \I__10786\ : LocalMux
    port map (
            O => \N__45026\,
            I => comm_cmd_1
        );

    \I__10785\ : Odrv4
    port map (
            O => \N__45019\,
            I => comm_cmd_1
        );

    \I__10784\ : Odrv4
    port map (
            O => \N__45006\,
            I => comm_cmd_1
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__45001\,
            I => comm_cmd_1
        );

    \I__10782\ : Odrv4
    port map (
            O => \N__44996\,
            I => comm_cmd_1
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__44991\,
            I => comm_cmd_1
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__44986\,
            I => comm_cmd_1
        );

    \I__10779\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44964\
        );

    \I__10778\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44960\
        );

    \I__10777\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44957\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__44964\,
            I => \N__44954\
        );

    \I__10775\ : InMux
    port map (
            O => \N__44963\,
            I => \N__44951\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__44960\,
            I => \N__44948\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__44957\,
            I => \N__44945\
        );

    \I__10772\ : Span4Mux_h
    port map (
            O => \N__44954\,
            I => \N__44942\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__44951\,
            I => \N__44939\
        );

    \I__10770\ : Span4Mux_h
    port map (
            O => \N__44948\,
            I => \N__44934\
        );

    \I__10769\ : Span4Mux_h
    port map (
            O => \N__44945\,
            I => \N__44934\
        );

    \I__10768\ : Span4Mux_v
    port map (
            O => \N__44942\,
            I => \N__44931\
        );

    \I__10767\ : Span4Mux_h
    port map (
            O => \N__44939\,
            I => \N__44926\
        );

    \I__10766\ : Span4Mux_v
    port map (
            O => \N__44934\,
            I => \N__44926\
        );

    \I__10765\ : Odrv4
    port map (
            O => \N__44931\,
            I => n9
        );

    \I__10764\ : Odrv4
    port map (
            O => \N__44926\,
            I => n9
        );

    \I__10763\ : InMux
    port map (
            O => \N__44921\,
            I => \N__44918\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__44918\,
            I => \N__44914\
        );

    \I__10761\ : InMux
    port map (
            O => \N__44917\,
            I => \N__44911\
        );

    \I__10760\ : Span4Mux_v
    port map (
            O => \N__44914\,
            I => \N__44904\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__44911\,
            I => \N__44901\
        );

    \I__10758\ : InMux
    port map (
            O => \N__44910\,
            I => \N__44898\
        );

    \I__10757\ : InMux
    port map (
            O => \N__44909\,
            I => \N__44895\
        );

    \I__10756\ : InMux
    port map (
            O => \N__44908\,
            I => \N__44892\
        );

    \I__10755\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44889\
        );

    \I__10754\ : Span4Mux_h
    port map (
            O => \N__44904\,
            I => \N__44874\
        );

    \I__10753\ : Span4Mux_v
    port map (
            O => \N__44901\,
            I => \N__44874\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__44898\,
            I => \N__44874\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44874\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__44892\,
            I => \N__44869\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__44889\,
            I => \N__44869\
        );

    \I__10748\ : InMux
    port map (
            O => \N__44888\,
            I => \N__44866\
        );

    \I__10747\ : InMux
    port map (
            O => \N__44887\,
            I => \N__44863\
        );

    \I__10746\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44860\
        );

    \I__10745\ : InMux
    port map (
            O => \N__44885\,
            I => \N__44857\
        );

    \I__10744\ : InMux
    port map (
            O => \N__44884\,
            I => \N__44853\
        );

    \I__10743\ : CascadeMux
    port map (
            O => \N__44883\,
            I => \N__44850\
        );

    \I__10742\ : Span4Mux_v
    port map (
            O => \N__44874\,
            I => \N__44847\
        );

    \I__10741\ : Span4Mux_v
    port map (
            O => \N__44869\,
            I => \N__44844\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__44866\,
            I => \N__44839\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__44863\,
            I => \N__44839\
        );

    \I__10738\ : LocalMux
    port map (
            O => \N__44860\,
            I => \N__44834\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__44857\,
            I => \N__44834\
        );

    \I__10736\ : InMux
    port map (
            O => \N__44856\,
            I => \N__44831\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__44853\,
            I => \N__44828\
        );

    \I__10734\ : InMux
    port map (
            O => \N__44850\,
            I => \N__44825\
        );

    \I__10733\ : Span4Mux_h
    port map (
            O => \N__44847\,
            I => \N__44822\
        );

    \I__10732\ : Span4Mux_h
    port map (
            O => \N__44844\,
            I => \N__44813\
        );

    \I__10731\ : Span4Mux_v
    port map (
            O => \N__44839\,
            I => \N__44813\
        );

    \I__10730\ : Span4Mux_v
    port map (
            O => \N__44834\,
            I => \N__44813\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__44831\,
            I => \N__44813\
        );

    \I__10728\ : Span4Mux_v
    port map (
            O => \N__44828\,
            I => \N__44808\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__44825\,
            I => \N__44808\
        );

    \I__10726\ : Span4Mux_h
    port map (
            O => \N__44822\,
            I => \N__44804\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__44813\,
            I => \N__44801\
        );

    \I__10724\ : Span4Mux_v
    port map (
            O => \N__44808\,
            I => \N__44798\
        );

    \I__10723\ : InMux
    port map (
            O => \N__44807\,
            I => \N__44795\
        );

    \I__10722\ : Odrv4
    port map (
            O => \N__44804\,
            I => comm_rx_buf_3
        );

    \I__10721\ : Odrv4
    port map (
            O => \N__44801\,
            I => comm_rx_buf_3
        );

    \I__10720\ : Odrv4
    port map (
            O => \N__44798\,
            I => comm_rx_buf_3
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__44795\,
            I => comm_rx_buf_3
        );

    \I__10718\ : InMux
    port map (
            O => \N__44786\,
            I => \N__44783\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__44783\,
            I => \N__44780\
        );

    \I__10716\ : Odrv4
    port map (
            O => \N__44780\,
            I => n4261
        );

    \I__10715\ : CascadeMux
    port map (
            O => \N__44777\,
            I => \N__44771\
        );

    \I__10714\ : InMux
    port map (
            O => \N__44776\,
            I => \N__44768\
        );

    \I__10713\ : CascadeMux
    port map (
            O => \N__44775\,
            I => \N__44765\
        );

    \I__10712\ : InMux
    port map (
            O => \N__44774\,
            I => \N__44761\
        );

    \I__10711\ : InMux
    port map (
            O => \N__44771\,
            I => \N__44758\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__44768\,
            I => \N__44755\
        );

    \I__10709\ : InMux
    port map (
            O => \N__44765\,
            I => \N__44752\
        );

    \I__10708\ : InMux
    port map (
            O => \N__44764\,
            I => \N__44749\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__44761\,
            I => \N__44746\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__44758\,
            I => \N__44743\
        );

    \I__10705\ : Span4Mux_h
    port map (
            O => \N__44755\,
            I => \N__44740\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__44752\,
            I => \N__44737\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__44749\,
            I => \N__44732\
        );

    \I__10702\ : Span4Mux_h
    port map (
            O => \N__44746\,
            I => \N__44732\
        );

    \I__10701\ : Span4Mux_h
    port map (
            O => \N__44743\,
            I => \N__44727\
        );

    \I__10700\ : Span4Mux_h
    port map (
            O => \N__44740\,
            I => \N__44727\
        );

    \I__10699\ : Span4Mux_h
    port map (
            O => \N__44737\,
            I => \N__44722\
        );

    \I__10698\ : Span4Mux_v
    port map (
            O => \N__44732\,
            I => \N__44722\
        );

    \I__10697\ : Odrv4
    port map (
            O => \N__44727\,
            I => comm_buf_1_3
        );

    \I__10696\ : Odrv4
    port map (
            O => \N__44722\,
            I => comm_buf_1_3
        );

    \I__10695\ : CEMux
    port map (
            O => \N__44717\,
            I => \N__44713\
        );

    \I__10694\ : CEMux
    port map (
            O => \N__44716\,
            I => \N__44708\
        );

    \I__10693\ : LocalMux
    port map (
            O => \N__44713\,
            I => \N__44705\
        );

    \I__10692\ : CEMux
    port map (
            O => \N__44712\,
            I => \N__44702\
        );

    \I__10691\ : CEMux
    port map (
            O => \N__44711\,
            I => \N__44699\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__44708\,
            I => \N__44695\
        );

    \I__10689\ : Span4Mux_v
    port map (
            O => \N__44705\,
            I => \N__44690\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__44702\,
            I => \N__44690\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__44699\,
            I => \N__44687\
        );

    \I__10686\ : CEMux
    port map (
            O => \N__44698\,
            I => \N__44684\
        );

    \I__10685\ : Span4Mux_v
    port map (
            O => \N__44695\,
            I => \N__44681\
        );

    \I__10684\ : Span4Mux_h
    port map (
            O => \N__44690\,
            I => \N__44678\
        );

    \I__10683\ : Span4Mux_h
    port map (
            O => \N__44687\,
            I => \N__44673\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__44684\,
            I => \N__44673\
        );

    \I__10681\ : Span4Mux_h
    port map (
            O => \N__44681\,
            I => \N__44670\
        );

    \I__10680\ : Span4Mux_h
    port map (
            O => \N__44678\,
            I => \N__44667\
        );

    \I__10679\ : Span4Mux_v
    port map (
            O => \N__44673\,
            I => \N__44664\
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__44670\,
            I => n8702
        );

    \I__10677\ : Odrv4
    port map (
            O => \N__44667\,
            I => n8702
        );

    \I__10676\ : Odrv4
    port map (
            O => \N__44664\,
            I => n8702
        );

    \I__10675\ : SRMux
    port map (
            O => \N__44657\,
            I => \N__44654\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__44654\,
            I => \N__44649\
        );

    \I__10673\ : SRMux
    port map (
            O => \N__44653\,
            I => \N__44646\
        );

    \I__10672\ : SRMux
    port map (
            O => \N__44652\,
            I => \N__44642\
        );

    \I__10671\ : Span4Mux_v
    port map (
            O => \N__44649\,
            I => \N__44636\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__44646\,
            I => \N__44636\
        );

    \I__10669\ : SRMux
    port map (
            O => \N__44645\,
            I => \N__44633\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__44642\,
            I => \N__44630\
        );

    \I__10667\ : SRMux
    port map (
            O => \N__44641\,
            I => \N__44627\
        );

    \I__10666\ : Span4Mux_h
    port map (
            O => \N__44636\,
            I => \N__44622\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__44633\,
            I => \N__44622\
        );

    \I__10664\ : Span4Mux_v
    port map (
            O => \N__44630\,
            I => \N__44617\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__44627\,
            I => \N__44617\
        );

    \I__10662\ : Span4Mux_h
    port map (
            O => \N__44622\,
            I => \N__44614\
        );

    \I__10661\ : Span4Mux_h
    port map (
            O => \N__44617\,
            I => \N__44611\
        );

    \I__10660\ : Span4Mux_h
    port map (
            O => \N__44614\,
            I => \N__44608\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__44611\,
            I => n10583
        );

    \I__10658\ : Odrv4
    port map (
            O => \N__44608\,
            I => n10583
        );

    \I__10657\ : InMux
    port map (
            O => \N__44603\,
            I => \N__44599\
        );

    \I__10656\ : CascadeMux
    port map (
            O => \N__44602\,
            I => \N__44596\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__44599\,
            I => \N__44593\
        );

    \I__10654\ : InMux
    port map (
            O => \N__44596\,
            I => \N__44590\
        );

    \I__10653\ : Span4Mux_h
    port map (
            O => \N__44593\,
            I => \N__44587\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__44590\,
            I => \N__44584\
        );

    \I__10651\ : Span4Mux_h
    port map (
            O => \N__44587\,
            I => \N__44580\
        );

    \I__10650\ : Span4Mux_v
    port map (
            O => \N__44584\,
            I => \N__44577\
        );

    \I__10649\ : InMux
    port map (
            O => \N__44583\,
            I => \N__44574\
        );

    \I__10648\ : Odrv4
    port map (
            O => \N__44580\,
            I => cmd_rdadctmp_21
        );

    \I__10647\ : Odrv4
    port map (
            O => \N__44577\,
            I => cmd_rdadctmp_21
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__44574\,
            I => cmd_rdadctmp_21
        );

    \I__10645\ : CascadeMux
    port map (
            O => \N__44567\,
            I => \N__44564\
        );

    \I__10644\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44560\
        );

    \I__10643\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44557\
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__44560\,
            I => \N__44552\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__44557\,
            I => \N__44552\
        );

    \I__10640\ : Odrv4
    port map (
            O => \N__44552\,
            I => buf_adcdata1_13
        );

    \I__10639\ : CascadeMux
    port map (
            O => \N__44549\,
            I => \N__44546\
        );

    \I__10638\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44543\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__44543\,
            I => \N__44539\
        );

    \I__10636\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44536\
        );

    \I__10635\ : Span4Mux_h
    port map (
            O => \N__44539\,
            I => \N__44532\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__44536\,
            I => \N__44529\
        );

    \I__10633\ : CascadeMux
    port map (
            O => \N__44535\,
            I => \N__44526\
        );

    \I__10632\ : Span4Mux_h
    port map (
            O => \N__44532\,
            I => \N__44523\
        );

    \I__10631\ : Span4Mux_h
    port map (
            O => \N__44529\,
            I => \N__44520\
        );

    \I__10630\ : InMux
    port map (
            O => \N__44526\,
            I => \N__44517\
        );

    \I__10629\ : Odrv4
    port map (
            O => \N__44523\,
            I => cmd_rdadctmp_17_adj_1095
        );

    \I__10628\ : Odrv4
    port map (
            O => \N__44520\,
            I => cmd_rdadctmp_17_adj_1095
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__44517\,
            I => cmd_rdadctmp_17_adj_1095
        );

    \I__10626\ : InMux
    port map (
            O => \N__44510\,
            I => \N__44505\
        );

    \I__10625\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44502\
        );

    \I__10624\ : CascadeMux
    port map (
            O => \N__44508\,
            I => \N__44499\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__44505\,
            I => \N__44494\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__44502\,
            I => \N__44494\
        );

    \I__10621\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44491\
        );

    \I__10620\ : Odrv12
    port map (
            O => \N__44494\,
            I => cmd_rdadctmp_18_adj_1094
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__44491\,
            I => cmd_rdadctmp_18_adj_1094
        );

    \I__10618\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44482\
        );

    \I__10617\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44479\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__44482\,
            I => \N__44476\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__44479\,
            I => buf_adcdata2_13
        );

    \I__10614\ : Odrv4
    port map (
            O => \N__44476\,
            I => buf_adcdata2_13
        );

    \I__10613\ : CascadeMux
    port map (
            O => \N__44471\,
            I => \N__44468\
        );

    \I__10612\ : InMux
    port map (
            O => \N__44468\,
            I => \N__44465\
        );

    \I__10611\ : LocalMux
    port map (
            O => \N__44465\,
            I => \N__44461\
        );

    \I__10610\ : InMux
    port map (
            O => \N__44464\,
            I => \N__44458\
        );

    \I__10609\ : Span4Mux_v
    port map (
            O => \N__44461\,
            I => \N__44455\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__44458\,
            I => \N__44452\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__44455\,
            I => \N__44448\
        );

    \I__10606\ : Span4Mux_v
    port map (
            O => \N__44452\,
            I => \N__44445\
        );

    \I__10605\ : CascadeMux
    port map (
            O => \N__44451\,
            I => \N__44442\
        );

    \I__10604\ : Sp12to4
    port map (
            O => \N__44448\,
            I => \N__44439\
        );

    \I__10603\ : Span4Mux_h
    port map (
            O => \N__44445\,
            I => \N__44436\
        );

    \I__10602\ : InMux
    port map (
            O => \N__44442\,
            I => \N__44433\
        );

    \I__10601\ : Odrv12
    port map (
            O => \N__44439\,
            I => cmd_rdadctmp_10
        );

    \I__10600\ : Odrv4
    port map (
            O => \N__44436\,
            I => cmd_rdadctmp_10
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__44433\,
            I => cmd_rdadctmp_10
        );

    \I__10598\ : InMux
    port map (
            O => \N__44426\,
            I => \N__44423\
        );

    \I__10597\ : LocalMux
    port map (
            O => \N__44423\,
            I => \N__44420\
        );

    \I__10596\ : Span4Mux_h
    port map (
            O => \N__44420\,
            I => \N__44416\
        );

    \I__10595\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44413\
        );

    \I__10594\ : Span4Mux_v
    port map (
            O => \N__44416\,
            I => \N__44410\
        );

    \I__10593\ : LocalMux
    port map (
            O => \N__44413\,
            I => buf_adcdata1_2
        );

    \I__10592\ : Odrv4
    port map (
            O => \N__44410\,
            I => buf_adcdata1_2
        );

    \I__10591\ : InMux
    port map (
            O => \N__44405\,
            I => \N__44395\
        );

    \I__10590\ : InMux
    port map (
            O => \N__44404\,
            I => \N__44390\
        );

    \I__10589\ : InMux
    port map (
            O => \N__44403\,
            I => \N__44390\
        );

    \I__10588\ : InMux
    port map (
            O => \N__44402\,
            I => \N__44383\
        );

    \I__10587\ : InMux
    port map (
            O => \N__44401\,
            I => \N__44383\
        );

    \I__10586\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44383\
        );

    \I__10585\ : InMux
    port map (
            O => \N__44399\,
            I => \N__44379\
        );

    \I__10584\ : InMux
    port map (
            O => \N__44398\,
            I => \N__44376\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__44395\,
            I => \N__44373\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__44390\,
            I => \N__44370\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__44383\,
            I => \N__44364\
        );

    \I__10580\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44361\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44348\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__44376\,
            I => \N__44345\
        );

    \I__10577\ : Span4Mux_h
    port map (
            O => \N__44373\,
            I => \N__44340\
        );

    \I__10576\ : Span4Mux_v
    port map (
            O => \N__44370\,
            I => \N__44340\
        );

    \I__10575\ : InMux
    port map (
            O => \N__44369\,
            I => \N__44337\
        );

    \I__10574\ : InMux
    port map (
            O => \N__44368\,
            I => \N__44332\
        );

    \I__10573\ : InMux
    port map (
            O => \N__44367\,
            I => \N__44332\
        );

    \I__10572\ : Span4Mux_v
    port map (
            O => \N__44364\,
            I => \N__44326\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__44361\,
            I => \N__44326\
        );

    \I__10570\ : InMux
    port map (
            O => \N__44360\,
            I => \N__44321\
        );

    \I__10569\ : InMux
    port map (
            O => \N__44359\,
            I => \N__44321\
        );

    \I__10568\ : InMux
    port map (
            O => \N__44358\,
            I => \N__44314\
        );

    \I__10567\ : InMux
    port map (
            O => \N__44357\,
            I => \N__44314\
        );

    \I__10566\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44314\
        );

    \I__10565\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44311\
        );

    \I__10564\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44308\
        );

    \I__10563\ : InMux
    port map (
            O => \N__44353\,
            I => \N__44303\
        );

    \I__10562\ : InMux
    port map (
            O => \N__44352\,
            I => \N__44303\
        );

    \I__10561\ : InMux
    port map (
            O => \N__44351\,
            I => \N__44299\
        );

    \I__10560\ : Span4Mux_h
    port map (
            O => \N__44348\,
            I => \N__44294\
        );

    \I__10559\ : Span4Mux_v
    port map (
            O => \N__44345\,
            I => \N__44294\
        );

    \I__10558\ : Span4Mux_h
    port map (
            O => \N__44340\,
            I => \N__44289\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__44337\,
            I => \N__44289\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__44332\,
            I => \N__44286\
        );

    \I__10555\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44283\
        );

    \I__10554\ : Span4Mux_v
    port map (
            O => \N__44326\,
            I => \N__44280\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__44321\,
            I => \N__44277\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44274\
        );

    \I__10551\ : LocalMux
    port map (
            O => \N__44311\,
            I => \N__44269\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__44308\,
            I => \N__44269\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__44303\,
            I => \N__44266\
        );

    \I__10548\ : InMux
    port map (
            O => \N__44302\,
            I => \N__44263\
        );

    \I__10547\ : LocalMux
    port map (
            O => \N__44299\,
            I => \N__44260\
        );

    \I__10546\ : Span4Mux_h
    port map (
            O => \N__44294\,
            I => \N__44255\
        );

    \I__10545\ : Span4Mux_v
    port map (
            O => \N__44289\,
            I => \N__44255\
        );

    \I__10544\ : Span4Mux_v
    port map (
            O => \N__44286\,
            I => \N__44250\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__44283\,
            I => \N__44250\
        );

    \I__10542\ : Span4Mux_h
    port map (
            O => \N__44280\,
            I => \N__44247\
        );

    \I__10541\ : Span4Mux_v
    port map (
            O => \N__44277\,
            I => \N__44244\
        );

    \I__10540\ : Span4Mux_v
    port map (
            O => \N__44274\,
            I => \N__44241\
        );

    \I__10539\ : Span4Mux_v
    port map (
            O => \N__44269\,
            I => \N__44236\
        );

    \I__10538\ : Span4Mux_h
    port map (
            O => \N__44266\,
            I => \N__44236\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__44263\,
            I => \N__44233\
        );

    \I__10536\ : Span4Mux_v
    port map (
            O => \N__44260\,
            I => \N__44230\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__44255\,
            I => \N__44225\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__44250\,
            I => \N__44225\
        );

    \I__10533\ : Span4Mux_h
    port map (
            O => \N__44247\,
            I => \N__44214\
        );

    \I__10532\ : Span4Mux_v
    port map (
            O => \N__44244\,
            I => \N__44214\
        );

    \I__10531\ : Span4Mux_v
    port map (
            O => \N__44241\,
            I => \N__44214\
        );

    \I__10530\ : Span4Mux_v
    port map (
            O => \N__44236\,
            I => \N__44214\
        );

    \I__10529\ : Span4Mux_h
    port map (
            O => \N__44233\,
            I => \N__44214\
        );

    \I__10528\ : Odrv4
    port map (
            O => \N__44230\,
            I => n15147
        );

    \I__10527\ : Odrv4
    port map (
            O => \N__44225\,
            I => n15147
        );

    \I__10526\ : Odrv4
    port map (
            O => \N__44214\,
            I => n15147
        );

    \I__10525\ : InMux
    port map (
            O => \N__44207\,
            I => \N__44203\
        );

    \I__10524\ : CascadeMux
    port map (
            O => \N__44206\,
            I => \N__44200\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__44203\,
            I => \N__44196\
        );

    \I__10522\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44193\
        );

    \I__10521\ : InMux
    port map (
            O => \N__44199\,
            I => \N__44190\
        );

    \I__10520\ : Span12Mux_v
    port map (
            O => \N__44196\,
            I => \N__44187\
        );

    \I__10519\ : LocalMux
    port map (
            O => \N__44193\,
            I => buf_adcdata3_10
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__44190\,
            I => buf_adcdata3_10
        );

    \I__10517\ : Odrv12
    port map (
            O => \N__44187\,
            I => buf_adcdata3_10
        );

    \I__10516\ : InMux
    port map (
            O => \N__44180\,
            I => \N__44175\
        );

    \I__10515\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44172\
        );

    \I__10514\ : InMux
    port map (
            O => \N__44178\,
            I => \N__44168\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__44175\,
            I => \N__44163\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__44172\,
            I => \N__44163\
        );

    \I__10511\ : InMux
    port map (
            O => \N__44171\,
            I => \N__44160\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__44168\,
            I => \N__44152\
        );

    \I__10509\ : Span4Mux_v
    port map (
            O => \N__44163\,
            I => \N__44146\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__44160\,
            I => \N__44146\
        );

    \I__10507\ : InMux
    port map (
            O => \N__44159\,
            I => \N__44143\
        );

    \I__10506\ : InMux
    port map (
            O => \N__44158\,
            I => \N__44140\
        );

    \I__10505\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44136\
        );

    \I__10504\ : InMux
    port map (
            O => \N__44156\,
            I => \N__44133\
        );

    \I__10503\ : InMux
    port map (
            O => \N__44155\,
            I => \N__44130\
        );

    \I__10502\ : Span4Mux_v
    port map (
            O => \N__44152\,
            I => \N__44127\
        );

    \I__10501\ : InMux
    port map (
            O => \N__44151\,
            I => \N__44124\
        );

    \I__10500\ : Span4Mux_h
    port map (
            O => \N__44146\,
            I => \N__44119\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__44143\,
            I => \N__44119\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__44140\,
            I => \N__44116\
        );

    \I__10497\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44113\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__44136\,
            I => \N__44108\
        );

    \I__10495\ : LocalMux
    port map (
            O => \N__44133\,
            I => \N__44108\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__44130\,
            I => \N__44105\
        );

    \I__10493\ : Span4Mux_h
    port map (
            O => \N__44127\,
            I => \N__44100\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__44124\,
            I => \N__44100\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__44119\,
            I => \N__44095\
        );

    \I__10490\ : Span4Mux_h
    port map (
            O => \N__44116\,
            I => \N__44092\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__44113\,
            I => \N__44089\
        );

    \I__10488\ : Span4Mux_v
    port map (
            O => \N__44108\,
            I => \N__44086\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__44105\,
            I => \N__44081\
        );

    \I__10486\ : Span4Mux_v
    port map (
            O => \N__44100\,
            I => \N__44081\
        );

    \I__10485\ : InMux
    port map (
            O => \N__44099\,
            I => \N__44078\
        );

    \I__10484\ : InMux
    port map (
            O => \N__44098\,
            I => \N__44075\
        );

    \I__10483\ : Span4Mux_h
    port map (
            O => \N__44095\,
            I => \N__44071\
        );

    \I__10482\ : Sp12to4
    port map (
            O => \N__44092\,
            I => \N__44068\
        );

    \I__10481\ : Span4Mux_v
    port map (
            O => \N__44089\,
            I => \N__44065\
        );

    \I__10480\ : Sp12to4
    port map (
            O => \N__44086\,
            I => \N__44056\
        );

    \I__10479\ : Sp12to4
    port map (
            O => \N__44081\,
            I => \N__44056\
        );

    \I__10478\ : LocalMux
    port map (
            O => \N__44078\,
            I => \N__44056\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__44075\,
            I => \N__44056\
        );

    \I__10476\ : InMux
    port map (
            O => \N__44074\,
            I => \N__44053\
        );

    \I__10475\ : Odrv4
    port map (
            O => \N__44071\,
            I => comm_rx_buf_1
        );

    \I__10474\ : Odrv12
    port map (
            O => \N__44068\,
            I => comm_rx_buf_1
        );

    \I__10473\ : Odrv4
    port map (
            O => \N__44065\,
            I => comm_rx_buf_1
        );

    \I__10472\ : Odrv12
    port map (
            O => \N__44056\,
            I => comm_rx_buf_1
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__44053\,
            I => comm_rx_buf_1
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__44042\,
            I => \N__44036\
        );

    \I__10469\ : InMux
    port map (
            O => \N__44041\,
            I => \N__44029\
        );

    \I__10468\ : InMux
    port map (
            O => \N__44040\,
            I => \N__44024\
        );

    \I__10467\ : InMux
    port map (
            O => \N__44039\,
            I => \N__44024\
        );

    \I__10466\ : InMux
    port map (
            O => \N__44036\,
            I => \N__44021\
        );

    \I__10465\ : InMux
    port map (
            O => \N__44035\,
            I => \N__44012\
        );

    \I__10464\ : InMux
    port map (
            O => \N__44034\,
            I => \N__44012\
        );

    \I__10463\ : InMux
    port map (
            O => \N__44033\,
            I => \N__44012\
        );

    \I__10462\ : InMux
    port map (
            O => \N__44032\,
            I => \N__44012\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__44029\,
            I => n8618
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__44024\,
            I => n8618
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__44021\,
            I => n8618
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__44012\,
            I => n8618
        );

    \I__10457\ : CascadeMux
    port map (
            O => \N__44003\,
            I => \N__43998\
        );

    \I__10456\ : CascadeMux
    port map (
            O => \N__44002\,
            I => \N__43991\
        );

    \I__10455\ : InMux
    port map (
            O => \N__44001\,
            I => \N__43988\
        );

    \I__10454\ : InMux
    port map (
            O => \N__43998\,
            I => \N__43981\
        );

    \I__10453\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43981\
        );

    \I__10452\ : InMux
    port map (
            O => \N__43996\,
            I => \N__43981\
        );

    \I__10451\ : InMux
    port map (
            O => \N__43995\,
            I => \N__43974\
        );

    \I__10450\ : InMux
    port map (
            O => \N__43994\,
            I => \N__43974\
        );

    \I__10449\ : InMux
    port map (
            O => \N__43991\,
            I => \N__43974\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__43988\,
            I => n10363
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__43981\,
            I => n10363
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__43974\,
            I => n10363
        );

    \I__10445\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43963\
        );

    \I__10444\ : CascadeMux
    port map (
            O => \N__43966\,
            I => \N__43959\
        );

    \I__10443\ : LocalMux
    port map (
            O => \N__43963\,
            I => \N__43956\
        );

    \I__10442\ : CascadeMux
    port map (
            O => \N__43962\,
            I => \N__43953\
        );

    \I__10441\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43950\
        );

    \I__10440\ : Span12Mux_v
    port map (
            O => \N__43956\,
            I => \N__43947\
        );

    \I__10439\ : InMux
    port map (
            O => \N__43953\,
            I => \N__43944\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__43950\,
            I => cmd_rdadctmp_25_adj_1051
        );

    \I__10437\ : Odrv12
    port map (
            O => \N__43947\,
            I => cmd_rdadctmp_25_adj_1051
        );

    \I__10436\ : LocalMux
    port map (
            O => \N__43944\,
            I => cmd_rdadctmp_25_adj_1051
        );

    \I__10435\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43933\
        );

    \I__10434\ : CascadeMux
    port map (
            O => \N__43936\,
            I => \N__43930\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43927\
        );

    \I__10432\ : InMux
    port map (
            O => \N__43930\,
            I => \N__43924\
        );

    \I__10431\ : Span4Mux_h
    port map (
            O => \N__43927\,
            I => \N__43921\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__43924\,
            I => buf_adcdata2_18
        );

    \I__10429\ : Odrv4
    port map (
            O => \N__43921\,
            I => buf_adcdata2_18
        );

    \I__10428\ : CascadeMux
    port map (
            O => \N__43916\,
            I => \N__43913\
        );

    \I__10427\ : InMux
    port map (
            O => \N__43913\,
            I => \N__43910\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__43910\,
            I => \N__43906\
        );

    \I__10425\ : InMux
    port map (
            O => \N__43909\,
            I => \N__43903\
        );

    \I__10424\ : Span4Mux_h
    port map (
            O => \N__43906\,
            I => \N__43900\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__43903\,
            I => \N__43897\
        );

    \I__10422\ : Odrv4
    port map (
            O => \N__43900\,
            I => n14_adj_1215
        );

    \I__10421\ : Odrv12
    port map (
            O => \N__43897\,
            I => n14_adj_1215
        );

    \I__10420\ : CascadeMux
    port map (
            O => \N__43892\,
            I => \N__43887\
        );

    \I__10419\ : InMux
    port map (
            O => \N__43891\,
            I => \N__43880\
        );

    \I__10418\ : InMux
    port map (
            O => \N__43890\,
            I => \N__43880\
        );

    \I__10417\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43880\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__43880\,
            I => cmd_rdadctmp_26_adj_1050
        );

    \I__10415\ : CascadeMux
    port map (
            O => \N__43877\,
            I => \N__43874\
        );

    \I__10414\ : InMux
    port map (
            O => \N__43874\,
            I => \N__43870\
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__43873\,
            I => \N__43866\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43863\
        );

    \I__10411\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43858\
        );

    \I__10410\ : InMux
    port map (
            O => \N__43866\,
            I => \N__43858\
        );

    \I__10409\ : Odrv4
    port map (
            O => \N__43863\,
            I => cmd_rdadctmp_27_adj_1049
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__43858\,
            I => cmd_rdadctmp_27_adj_1049
        );

    \I__10407\ : CascadeMux
    port map (
            O => \N__43853\,
            I => \N__43850\
        );

    \I__10406\ : InMux
    port map (
            O => \N__43850\,
            I => \N__43847\
        );

    \I__10405\ : LocalMux
    port map (
            O => \N__43847\,
            I => \N__43844\
        );

    \I__10404\ : Span4Mux_v
    port map (
            O => \N__43844\,
            I => \N__43841\
        );

    \I__10403\ : Span4Mux_h
    port map (
            O => \N__43841\,
            I => \N__43837\
        );

    \I__10402\ : CascadeMux
    port map (
            O => \N__43840\,
            I => \N__43834\
        );

    \I__10401\ : Span4Mux_h
    port map (
            O => \N__43837\,
            I => \N__43831\
        );

    \I__10400\ : InMux
    port map (
            O => \N__43834\,
            I => \N__43828\
        );

    \I__10399\ : Span4Mux_h
    port map (
            O => \N__43831\,
            I => \N__43822\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__43828\,
            I => \N__43822\
        );

    \I__10397\ : InMux
    port map (
            O => \N__43827\,
            I => \N__43819\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__43822\,
            I => cmd_rdadctmp_8_adj_1104
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__43819\,
            I => cmd_rdadctmp_8_adj_1104
        );

    \I__10394\ : InMux
    port map (
            O => \N__43814\,
            I => \N__43811\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__43811\,
            I => \N__43807\
        );

    \I__10392\ : InMux
    port map (
            O => \N__43810\,
            I => \N__43804\
        );

    \I__10391\ : Sp12to4
    port map (
            O => \N__43807\,
            I => \N__43801\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__43804\,
            I => \N__43797\
        );

    \I__10389\ : Span12Mux_v
    port map (
            O => \N__43801\,
            I => \N__43794\
        );

    \I__10388\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43791\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__43797\,
            I => \N__43788\
        );

    \I__10386\ : Span12Mux_h
    port map (
            O => \N__43794\,
            I => \N__43785\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__43791\,
            I => buf_adcdata3_0
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__43788\,
            I => buf_adcdata3_0
        );

    \I__10383\ : Odrv12
    port map (
            O => \N__43785\,
            I => buf_adcdata3_0
        );

    \I__10382\ : InMux
    port map (
            O => \N__43778\,
            I => \N__43775\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__43775\,
            I => \N__43771\
        );

    \I__10380\ : InMux
    port map (
            O => \N__43774\,
            I => \N__43768\
        );

    \I__10379\ : Span4Mux_h
    port map (
            O => \N__43771\,
            I => \N__43764\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__43768\,
            I => \N__43761\
        );

    \I__10377\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43758\
        );

    \I__10376\ : Span4Mux_v
    port map (
            O => \N__43764\,
            I => \N__43753\
        );

    \I__10375\ : Span4Mux_h
    port map (
            O => \N__43761\,
            I => \N__43753\
        );

    \I__10374\ : LocalMux
    port map (
            O => \N__43758\,
            I => buf_adcdata3_11
        );

    \I__10373\ : Odrv4
    port map (
            O => \N__43753\,
            I => buf_adcdata3_11
        );

    \I__10372\ : CascadeMux
    port map (
            O => \N__43748\,
            I => \N__43745\
        );

    \I__10371\ : InMux
    port map (
            O => \N__43745\,
            I => \N__43742\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__43742\,
            I => \N__43739\
        );

    \I__10369\ : Span4Mux_v
    port map (
            O => \N__43739\,
            I => \N__43735\
        );

    \I__10368\ : CascadeMux
    port map (
            O => \N__43738\,
            I => \N__43731\
        );

    \I__10367\ : Span4Mux_h
    port map (
            O => \N__43735\,
            I => \N__43728\
        );

    \I__10366\ : InMux
    port map (
            O => \N__43734\,
            I => \N__43723\
        );

    \I__10365\ : InMux
    port map (
            O => \N__43731\,
            I => \N__43723\
        );

    \I__10364\ : Odrv4
    port map (
            O => \N__43728\,
            I => cmd_rdadctmp_30_adj_1082
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__43723\,
            I => cmd_rdadctmp_30_adj_1082
        );

    \I__10362\ : InMux
    port map (
            O => \N__43718\,
            I => \N__43715\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__43715\,
            I => \N__43712\
        );

    \I__10360\ : Span4Mux_h
    port map (
            O => \N__43712\,
            I => \N__43709\
        );

    \I__10359\ : Span4Mux_v
    port map (
            O => \N__43709\,
            I => \N__43704\
        );

    \I__10358\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43699\
        );

    \I__10357\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43699\
        );

    \I__10356\ : Odrv4
    port map (
            O => \N__43704\,
            I => buf_adcdata3_22
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__43699\,
            I => buf_adcdata3_22
        );

    \I__10354\ : InMux
    port map (
            O => \N__43694\,
            I => \N__43691\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__43691\,
            I => \N__43688\
        );

    \I__10352\ : Odrv4
    port map (
            O => \N__43688\,
            I => n7_adj_1190
        );

    \I__10351\ : InMux
    port map (
            O => \N__43685\,
            I => \N__43682\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__43682\,
            I => \N__43678\
        );

    \I__10349\ : InMux
    port map (
            O => \N__43681\,
            I => \N__43674\
        );

    \I__10348\ : Span4Mux_h
    port map (
            O => \N__43678\,
            I => \N__43671\
        );

    \I__10347\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43668\
        );

    \I__10346\ : LocalMux
    port map (
            O => \N__43674\,
            I => buf_dds_2
        );

    \I__10345\ : Odrv4
    port map (
            O => \N__43671\,
            I => buf_dds_2
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__43668\,
            I => buf_dds_2
        );

    \I__10343\ : CascadeMux
    port map (
            O => \N__43661\,
            I => \N__43658\
        );

    \I__10342\ : InMux
    port map (
            O => \N__43658\,
            I => \N__43655\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__43655\,
            I => \N__43652\
        );

    \I__10340\ : Span4Mux_v
    port map (
            O => \N__43652\,
            I => \N__43649\
        );

    \I__10339\ : Span4Mux_h
    port map (
            O => \N__43649\,
            I => \N__43646\
        );

    \I__10338\ : Odrv4
    port map (
            O => \N__43646\,
            I => n4207
        );

    \I__10337\ : InMux
    port map (
            O => \N__43643\,
            I => \N__43640\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__43640\,
            I => \N__43637\
        );

    \I__10335\ : Span4Mux_v
    port map (
            O => \N__43637\,
            I => \N__43632\
        );

    \I__10334\ : InMux
    port map (
            O => \N__43636\,
            I => \N__43629\
        );

    \I__10333\ : InMux
    port map (
            O => \N__43635\,
            I => \N__43626\
        );

    \I__10332\ : Span4Mux_h
    port map (
            O => \N__43632\,
            I => \N__43621\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__43629\,
            I => \N__43621\
        );

    \I__10330\ : LocalMux
    port map (
            O => \N__43626\,
            I => n8094
        );

    \I__10329\ : Odrv4
    port map (
            O => \N__43621\,
            I => n8094
        );

    \I__10328\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43611\
        );

    \I__10327\ : InMux
    port map (
            O => \N__43615\,
            I => \N__43608\
        );

    \I__10326\ : InMux
    port map (
            O => \N__43614\,
            I => \N__43605\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__43611\,
            I => \N__43602\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__43608\,
            I => \N__43599\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__43605\,
            I => \N__43596\
        );

    \I__10322\ : Span4Mux_v
    port map (
            O => \N__43602\,
            I => \N__43593\
        );

    \I__10321\ : Span4Mux_h
    port map (
            O => \N__43599\,
            I => \N__43590\
        );

    \I__10320\ : Span4Mux_v
    port map (
            O => \N__43596\,
            I => \N__43585\
        );

    \I__10319\ : Span4Mux_h
    port map (
            O => \N__43593\,
            I => \N__43585\
        );

    \I__10318\ : Odrv4
    port map (
            O => \N__43590\,
            I => n729
        );

    \I__10317\ : Odrv4
    port map (
            O => \N__43585\,
            I => n729
        );

    \I__10316\ : InMux
    port map (
            O => \N__43580\,
            I => \N__43577\
        );

    \I__10315\ : LocalMux
    port map (
            O => \N__43577\,
            I => \N__43573\
        );

    \I__10314\ : InMux
    port map (
            O => \N__43576\,
            I => \N__43570\
        );

    \I__10313\ : Span4Mux_h
    port map (
            O => \N__43573\,
            I => \N__43567\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__43570\,
            I => buf_adcdata2_19
        );

    \I__10311\ : Odrv4
    port map (
            O => \N__43567\,
            I => buf_adcdata2_19
        );

    \I__10310\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43555\
        );

    \I__10309\ : CascadeMux
    port map (
            O => \N__43561\,
            I => \N__43552\
        );

    \I__10308\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43549\
        );

    \I__10307\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43546\
        );

    \I__10306\ : InMux
    port map (
            O => \N__43558\,
            I => \N__43543\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__43555\,
            I => \N__43540\
        );

    \I__10304\ : InMux
    port map (
            O => \N__43552\,
            I => \N__43537\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__43549\,
            I => \N__43534\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__43546\,
            I => \N__43529\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__43543\,
            I => \N__43526\
        );

    \I__10300\ : Span4Mux_h
    port map (
            O => \N__43540\,
            I => \N__43523\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__43537\,
            I => \N__43518\
        );

    \I__10298\ : Span4Mux_v
    port map (
            O => \N__43534\,
            I => \N__43518\
        );

    \I__10297\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43515\
        );

    \I__10296\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43512\
        );

    \I__10295\ : Span12Mux_v
    port map (
            O => \N__43529\,
            I => \N__43509\
        );

    \I__10294\ : Span4Mux_h
    port map (
            O => \N__43526\,
            I => \N__43502\
        );

    \I__10293\ : Span4Mux_h
    port map (
            O => \N__43523\,
            I => \N__43502\
        );

    \I__10292\ : Span4Mux_h
    port map (
            O => \N__43518\,
            I => \N__43502\
        );

    \I__10291\ : LocalMux
    port map (
            O => \N__43515\,
            I => comm_buf_0_3
        );

    \I__10290\ : LocalMux
    port map (
            O => \N__43512\,
            I => comm_buf_0_3
        );

    \I__10289\ : Odrv12
    port map (
            O => \N__43509\,
            I => comm_buf_0_3
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__43502\,
            I => comm_buf_0_3
        );

    \I__10287\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43489\
        );

    \I__10286\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43486\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__43489\,
            I => \N__43481\
        );

    \I__10284\ : LocalMux
    port map (
            O => \N__43486\,
            I => \N__43481\
        );

    \I__10283\ : Span4Mux_v
    port map (
            O => \N__43481\,
            I => \N__43478\
        );

    \I__10282\ : Span4Mux_h
    port map (
            O => \N__43478\,
            I => \N__43475\
        );

    \I__10281\ : Odrv4
    port map (
            O => \N__43475\,
            I => n14_adj_1208
        );

    \I__10280\ : CascadeMux
    port map (
            O => \N__43472\,
            I => \n26_adj_1192_cascade_\
        );

    \I__10279\ : CEMux
    port map (
            O => \N__43469\,
            I => \N__43466\
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__43466\,
            I => \N__43463\
        );

    \I__10277\ : Odrv4
    port map (
            O => \N__43463\,
            I => n18_adj_1191
        );

    \I__10276\ : InMux
    port map (
            O => \N__43460\,
            I => \N__43457\
        );

    \I__10275\ : LocalMux
    port map (
            O => \N__43457\,
            I => n15245
        );

    \I__10274\ : InMux
    port map (
            O => \N__43454\,
            I => \N__43451\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__43451\,
            I => \N__43442\
        );

    \I__10272\ : InMux
    port map (
            O => \N__43450\,
            I => \N__43433\
        );

    \I__10271\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43430\
        );

    \I__10270\ : InMux
    port map (
            O => \N__43448\,
            I => \N__43421\
        );

    \I__10269\ : InMux
    port map (
            O => \N__43447\,
            I => \N__43421\
        );

    \I__10268\ : InMux
    port map (
            O => \N__43446\,
            I => \N__43421\
        );

    \I__10267\ : InMux
    port map (
            O => \N__43445\,
            I => \N__43421\
        );

    \I__10266\ : Span4Mux_v
    port map (
            O => \N__43442\,
            I => \N__43418\
        );

    \I__10265\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43413\
        );

    \I__10264\ : InMux
    port map (
            O => \N__43440\,
            I => \N__43413\
        );

    \I__10263\ : CascadeMux
    port map (
            O => \N__43439\,
            I => \N__43410\
        );

    \I__10262\ : CascadeMux
    port map (
            O => \N__43438\,
            I => \N__43407\
        );

    \I__10261\ : CascadeMux
    port map (
            O => \N__43437\,
            I => \N__43403\
        );

    \I__10260\ : CascadeMux
    port map (
            O => \N__43436\,
            I => \N__43399\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__43433\,
            I => \N__43395\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__43430\,
            I => \N__43388\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__43421\,
            I => \N__43385\
        );

    \I__10256\ : Span4Mux_v
    port map (
            O => \N__43418\,
            I => \N__43380\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__43413\,
            I => \N__43380\
        );

    \I__10254\ : InMux
    port map (
            O => \N__43410\,
            I => \N__43376\
        );

    \I__10253\ : InMux
    port map (
            O => \N__43407\,
            I => \N__43371\
        );

    \I__10252\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43371\
        );

    \I__10251\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43362\
        );

    \I__10250\ : InMux
    port map (
            O => \N__43402\,
            I => \N__43362\
        );

    \I__10249\ : InMux
    port map (
            O => \N__43399\,
            I => \N__43362\
        );

    \I__10248\ : InMux
    port map (
            O => \N__43398\,
            I => \N__43362\
        );

    \I__10247\ : Sp12to4
    port map (
            O => \N__43395\,
            I => \N__43359\
        );

    \I__10246\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43350\
        );

    \I__10245\ : InMux
    port map (
            O => \N__43393\,
            I => \N__43350\
        );

    \I__10244\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43350\
        );

    \I__10243\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43350\
        );

    \I__10242\ : Span4Mux_v
    port map (
            O => \N__43388\,
            I => \N__43343\
        );

    \I__10241\ : Span4Mux_v
    port map (
            O => \N__43385\,
            I => \N__43343\
        );

    \I__10240\ : Span4Mux_h
    port map (
            O => \N__43380\,
            I => \N__43343\
        );

    \I__10239\ : InMux
    port map (
            O => \N__43379\,
            I => \N__43340\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__43376\,
            I => \N__43333\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__43371\,
            I => \N__43333\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__43362\,
            I => \N__43333\
        );

    \I__10235\ : Span12Mux_h
    port map (
            O => \N__43359\,
            I => \N__43330\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__43350\,
            I => \N__43323\
        );

    \I__10233\ : Sp12to4
    port map (
            O => \N__43343\,
            I => \N__43323\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__43340\,
            I => \N__43323\
        );

    \I__10231\ : Span12Mux_h
    port map (
            O => \N__43333\,
            I => \N__43320\
        );

    \I__10230\ : Span12Mux_v
    port map (
            O => \N__43330\,
            I => \N__43317\
        );

    \I__10229\ : Span12Mux_v
    port map (
            O => \N__43323\,
            I => \N__43314\
        );

    \I__10228\ : Span12Mux_v
    port map (
            O => \N__43320\,
            I => \N__43311\
        );

    \I__10227\ : Odrv12
    port map (
            O => \N__43317\,
            I => \ICE_SPI_CE0\
        );

    \I__10226\ : Odrv12
    port map (
            O => \N__43314\,
            I => \ICE_SPI_CE0\
        );

    \I__10225\ : Odrv12
    port map (
            O => \N__43311\,
            I => \ICE_SPI_CE0\
        );

    \I__10224\ : CascadeMux
    port map (
            O => \N__43304\,
            I => \n15245_cascade_\
        );

    \I__10223\ : InMux
    port map (
            O => \N__43301\,
            I => \N__43290\
        );

    \I__10222\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43290\
        );

    \I__10221\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43290\
        );

    \I__10220\ : InMux
    port map (
            O => \N__43298\,
            I => \N__43282\
        );

    \I__10219\ : InMux
    port map (
            O => \N__43297\,
            I => \N__43282\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__43290\,
            I => \N__43278\
        );

    \I__10217\ : InMux
    port map (
            O => \N__43289\,
            I => \N__43275\
        );

    \I__10216\ : InMux
    port map (
            O => \N__43288\,
            I => \N__43272\
        );

    \I__10215\ : InMux
    port map (
            O => \N__43287\,
            I => \N__43269\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__43282\,
            I => \N__43262\
        );

    \I__10213\ : InMux
    port map (
            O => \N__43281\,
            I => \N__43259\
        );

    \I__10212\ : Span4Mux_h
    port map (
            O => \N__43278\,
            I => \N__43256\
        );

    \I__10211\ : LocalMux
    port map (
            O => \N__43275\,
            I => \N__43248\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__43272\,
            I => \N__43248\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__43269\,
            I => \N__43248\
        );

    \I__10208\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43239\
        );

    \I__10207\ : InMux
    port map (
            O => \N__43267\,
            I => \N__43239\
        );

    \I__10206\ : InMux
    port map (
            O => \N__43266\,
            I => \N__43239\
        );

    \I__10205\ : InMux
    port map (
            O => \N__43265\,
            I => \N__43239\
        );

    \I__10204\ : Span4Mux_v
    port map (
            O => \N__43262\,
            I => \N__43235\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__43259\,
            I => \N__43232\
        );

    \I__10202\ : Span4Mux_h
    port map (
            O => \N__43256\,
            I => \N__43229\
        );

    \I__10201\ : InMux
    port map (
            O => \N__43255\,
            I => \N__43226\
        );

    \I__10200\ : Span4Mux_v
    port map (
            O => \N__43248\,
            I => \N__43221\
        );

    \I__10199\ : LocalMux
    port map (
            O => \N__43239\,
            I => \N__43221\
        );

    \I__10198\ : InMux
    port map (
            O => \N__43238\,
            I => \N__43218\
        );

    \I__10197\ : Odrv4
    port map (
            O => \N__43235\,
            I => comm_data_vld
        );

    \I__10196\ : Odrv4
    port map (
            O => \N__43232\,
            I => comm_data_vld
        );

    \I__10195\ : Odrv4
    port map (
            O => \N__43229\,
            I => comm_data_vld
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__43226\,
            I => comm_data_vld
        );

    \I__10193\ : Odrv4
    port map (
            O => \N__43221\,
            I => comm_data_vld
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__43218\,
            I => comm_data_vld
        );

    \I__10191\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43202\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__43202\,
            I => n8544
        );

    \I__10189\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43194\
        );

    \I__10188\ : InMux
    port map (
            O => \N__43198\,
            I => \N__43189\
        );

    \I__10187\ : InMux
    port map (
            O => \N__43197\,
            I => \N__43189\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__43194\,
            I => \N__43185\
        );

    \I__10185\ : LocalMux
    port map (
            O => \N__43189\,
            I => \N__43182\
        );

    \I__10184\ : InMux
    port map (
            O => \N__43188\,
            I => \N__43179\
        );

    \I__10183\ : Span4Mux_v
    port map (
            O => \N__43185\,
            I => \N__43174\
        );

    \I__10182\ : Span4Mux_v
    port map (
            O => \N__43182\,
            I => \N__43174\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__43179\,
            I => \N__43171\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__43174\,
            I => n9_adj_1028
        );

    \I__10179\ : Odrv12
    port map (
            O => \N__43171\,
            I => n9_adj_1028
        );

    \I__10178\ : CascadeMux
    port map (
            O => \N__43166\,
            I => \N__43162\
        );

    \I__10177\ : InMux
    port map (
            O => \N__43165\,
            I => \N__43159\
        );

    \I__10176\ : InMux
    port map (
            O => \N__43162\,
            I => \N__43156\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__43159\,
            I => \N__43153\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__43156\,
            I => \N__43150\
        );

    \I__10173\ : Span4Mux_h
    port map (
            O => \N__43153\,
            I => \N__43145\
        );

    \I__10172\ : Span4Mux_v
    port map (
            O => \N__43150\,
            I => \N__43145\
        );

    \I__10171\ : Odrv4
    port map (
            O => \N__43145\,
            I => n9011
        );

    \I__10170\ : CascadeMux
    port map (
            O => \N__43142\,
            I => \n9011_cascade_\
        );

    \I__10169\ : CEMux
    port map (
            O => \N__43139\,
            I => \N__43135\
        );

    \I__10168\ : CEMux
    port map (
            O => \N__43138\,
            I => \N__43131\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__43135\,
            I => \N__43128\
        );

    \I__10166\ : CEMux
    port map (
            O => \N__43134\,
            I => \N__43123\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__43131\,
            I => \N__43117\
        );

    \I__10164\ : Span4Mux_v
    port map (
            O => \N__43128\,
            I => \N__43117\
        );

    \I__10163\ : CEMux
    port map (
            O => \N__43127\,
            I => \N__43114\
        );

    \I__10162\ : CEMux
    port map (
            O => \N__43126\,
            I => \N__43111\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__43123\,
            I => \N__43106\
        );

    \I__10160\ : CEMux
    port map (
            O => \N__43122\,
            I => \N__43103\
        );

    \I__10159\ : Span4Mux_h
    port map (
            O => \N__43117\,
            I => \N__43096\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__43114\,
            I => \N__43096\
        );

    \I__10157\ : LocalMux
    port map (
            O => \N__43111\,
            I => \N__43096\
        );

    \I__10156\ : CEMux
    port map (
            O => \N__43110\,
            I => \N__43093\
        );

    \I__10155\ : CEMux
    port map (
            O => \N__43109\,
            I => \N__43090\
        );

    \I__10154\ : Span4Mux_v
    port map (
            O => \N__43106\,
            I => \N__43085\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__43103\,
            I => \N__43085\
        );

    \I__10152\ : Span4Mux_v
    port map (
            O => \N__43096\,
            I => \N__43082\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__43093\,
            I => \N__43079\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__43090\,
            I => \N__43075\
        );

    \I__10149\ : Span4Mux_v
    port map (
            O => \N__43085\,
            I => \N__43072\
        );

    \I__10148\ : Sp12to4
    port map (
            O => \N__43082\,
            I => \N__43069\
        );

    \I__10147\ : Sp12to4
    port map (
            O => \N__43079\,
            I => \N__43066\
        );

    \I__10146\ : InMux
    port map (
            O => \N__43078\,
            I => \N__43063\
        );

    \I__10145\ : Sp12to4
    port map (
            O => \N__43075\,
            I => \N__43058\
        );

    \I__10144\ : Sp12to4
    port map (
            O => \N__43072\,
            I => \N__43058\
        );

    \I__10143\ : Span12Mux_v
    port map (
            O => \N__43069\,
            I => \N__43051\
        );

    \I__10142\ : Span12Mux_v
    port map (
            O => \N__43066\,
            I => \N__43051\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__43063\,
            I => \N__43051\
        );

    \I__10140\ : Span12Mux_h
    port map (
            O => \N__43058\,
            I => \N__43048\
        );

    \I__10139\ : Span12Mux_h
    port map (
            O => \N__43051\,
            I => \N__43045\
        );

    \I__10138\ : Odrv12
    port map (
            O => \N__43048\,
            I => n9215
        );

    \I__10137\ : Odrv12
    port map (
            O => \N__43045\,
            I => n9215
        );

    \I__10136\ : InMux
    port map (
            O => \N__43040\,
            I => \N__43037\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__43037\,
            I => \N__43034\
        );

    \I__10134\ : Odrv4
    port map (
            O => \N__43034\,
            I => buf_data2_19
        );

    \I__10133\ : InMux
    port map (
            O => \N__43031\,
            I => \N__43028\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__43028\,
            I => \N__43025\
        );

    \I__10131\ : Span4Mux_h
    port map (
            O => \N__43025\,
            I => \N__43021\
        );

    \I__10130\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43018\
        );

    \I__10129\ : Sp12to4
    port map (
            O => \N__43021\,
            I => \N__43012\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__43018\,
            I => \N__43012\
        );

    \I__10127\ : InMux
    port map (
            O => \N__43017\,
            I => \N__43009\
        );

    \I__10126\ : Span12Mux_v
    port map (
            O => \N__43012\,
            I => \N__43006\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__43009\,
            I => buf_adcdata4_19
        );

    \I__10124\ : Odrv12
    port map (
            O => \N__43006\,
            I => buf_adcdata4_19
        );

    \I__10123\ : InMux
    port map (
            O => \N__43001\,
            I => \N__42998\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__42998\,
            I => \N__42995\
        );

    \I__10121\ : Sp12to4
    port map (
            O => \N__42995\,
            I => \N__42992\
        );

    \I__10120\ : Span12Mux_v
    port map (
            O => \N__42992\,
            I => \N__42989\
        );

    \I__10119\ : Odrv12
    port map (
            O => \N__42989\,
            I => \comm_buf_3_7_N_501_3\
        );

    \I__10118\ : CascadeMux
    port map (
            O => \N__42986\,
            I => \N__42982\
        );

    \I__10117\ : CascadeMux
    port map (
            O => \N__42985\,
            I => \N__42979\
        );

    \I__10116\ : InMux
    port map (
            O => \N__42982\,
            I => \N__42976\
        );

    \I__10115\ : InMux
    port map (
            O => \N__42979\,
            I => \N__42973\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__42976\,
            I => buf_control_6
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__42973\,
            I => buf_control_6
        );

    \I__10112\ : InMux
    port map (
            O => \N__42968\,
            I => \N__42965\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__42965\,
            I => \N__42962\
        );

    \I__10110\ : Span4Mux_h
    port map (
            O => \N__42962\,
            I => \N__42959\
        );

    \I__10109\ : Span4Mux_h
    port map (
            O => \N__42959\,
            I => \N__42956\
        );

    \I__10108\ : Odrv4
    port map (
            O => \N__42956\,
            I => n60
        );

    \I__10107\ : SRMux
    port map (
            O => \N__42953\,
            I => \N__42950\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__42950\,
            I => \N__42947\
        );

    \I__10105\ : Odrv12
    port map (
            O => \N__42947\,
            I => \comm_spi.imosi_N_791\
        );

    \I__10104\ : CascadeMux
    port map (
            O => \N__42944\,
            I => \N__42941\
        );

    \I__10103\ : InMux
    port map (
            O => \N__42941\,
            I => \N__42938\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__42938\,
            I => \N__42935\
        );

    \I__10101\ : Span4Mux_v
    port map (
            O => \N__42935\,
            I => \N__42932\
        );

    \I__10100\ : Sp12to4
    port map (
            O => \N__42932\,
            I => \N__42928\
        );

    \I__10099\ : CascadeMux
    port map (
            O => \N__42931\,
            I => \N__42924\
        );

    \I__10098\ : Span12Mux_h
    port map (
            O => \N__42928\,
            I => \N__42921\
        );

    \I__10097\ : InMux
    port map (
            O => \N__42927\,
            I => \N__42916\
        );

    \I__10096\ : InMux
    port map (
            O => \N__42924\,
            I => \N__42916\
        );

    \I__10095\ : Span12Mux_h
    port map (
            O => \N__42921\,
            I => \N__42913\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__42916\,
            I => cmd_rdadctmp_9_adj_1067
        );

    \I__10093\ : Odrv12
    port map (
            O => \N__42913\,
            I => cmd_rdadctmp_9_adj_1067
        );

    \I__10092\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42905\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__42905\,
            I => \N__42901\
        );

    \I__10090\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42898\
        );

    \I__10089\ : Span4Mux_v
    port map (
            O => \N__42901\,
            I => \N__42895\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__42898\,
            I => buf_adcdata2_1
        );

    \I__10087\ : Odrv4
    port map (
            O => \N__42895\,
            I => buf_adcdata2_1
        );

    \I__10086\ : InMux
    port map (
            O => \N__42890\,
            I => \N__42886\
        );

    \I__10085\ : InMux
    port map (
            O => \N__42889\,
            I => \N__42883\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__42886\,
            I => \comm_spi.imosi\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__42883\,
            I => \comm_spi.imosi\
        );

    \I__10082\ : SRMux
    port map (
            O => \N__42878\,
            I => \N__42875\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__42875\,
            I => \N__42872\
        );

    \I__10080\ : Span4Mux_h
    port map (
            O => \N__42872\,
            I => \N__42869\
        );

    \I__10079\ : Span4Mux_h
    port map (
            O => \N__42869\,
            I => \N__42866\
        );

    \I__10078\ : Odrv4
    port map (
            O => \N__42866\,
            I => \comm_spi.DOUT_7__N_786\
        );

    \I__10077\ : InMux
    port map (
            O => \N__42863\,
            I => \N__42857\
        );

    \I__10076\ : InMux
    port map (
            O => \N__42862\,
            I => \N__42857\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__42857\,
            I => \N__42853\
        );

    \I__10074\ : InMux
    port map (
            O => \N__42856\,
            I => \N__42850\
        );

    \I__10073\ : Span4Mux_v
    port map (
            O => \N__42853\,
            I => \N__42846\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__42850\,
            I => \N__42843\
        );

    \I__10071\ : InMux
    port map (
            O => \N__42849\,
            I => \N__42840\
        );

    \I__10070\ : Span4Mux_h
    port map (
            O => \N__42846\,
            I => \N__42833\
        );

    \I__10069\ : Span4Mux_v
    port map (
            O => \N__42843\,
            I => \N__42833\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__42840\,
            I => \N__42830\
        );

    \I__10067\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42825\
        );

    \I__10066\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42825\
        );

    \I__10065\ : Sp12to4
    port map (
            O => \N__42833\,
            I => \N__42820\
        );

    \I__10064\ : Span12Mux_h
    port map (
            O => \N__42830\,
            I => \N__42820\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__42825\,
            I => n15131
        );

    \I__10062\ : Odrv12
    port map (
            O => \N__42820\,
            I => n15131
        );

    \I__10061\ : CascadeMux
    port map (
            O => \N__42815\,
            I => \N__42812\
        );

    \I__10060\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42808\
        );

    \I__10059\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42805\
        );

    \I__10058\ : LocalMux
    port map (
            O => \N__42808\,
            I => n15241
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__42805\,
            I => n15241
        );

    \I__10056\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42788\
        );

    \I__10055\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42788\
        );

    \I__10054\ : InMux
    port map (
            O => \N__42798\,
            I => \N__42788\
        );

    \I__10053\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42785\
        );

    \I__10052\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42780\
        );

    \I__10051\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42780\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__42788\,
            I => \N__42775\
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__42785\,
            I => \N__42775\
        );

    \I__10048\ : LocalMux
    port map (
            O => \N__42780\,
            I => \N__42772\
        );

    \I__10047\ : Span4Mux_h
    port map (
            O => \N__42775\,
            I => \N__42769\
        );

    \I__10046\ : Span4Mux_h
    port map (
            O => \N__42772\,
            I => \N__42766\
        );

    \I__10045\ : Span4Mux_h
    port map (
            O => \N__42769\,
            I => \N__42763\
        );

    \I__10044\ : Span4Mux_h
    port map (
            O => \N__42766\,
            I => \N__42760\
        );

    \I__10043\ : Odrv4
    port map (
            O => \N__42763\,
            I => n15191
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__42760\,
            I => n15191
        );

    \I__10041\ : CascadeMux
    port map (
            O => \N__42755\,
            I => \N__42752\
        );

    \I__10040\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42749\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__42749\,
            I => \N__42745\
        );

    \I__10038\ : CascadeMux
    port map (
            O => \N__42748\,
            I => \N__42742\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__42745\,
            I => \N__42739\
        );

    \I__10036\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42736\
        );

    \I__10035\ : Odrv4
    port map (
            O => \N__42739\,
            I => n10148
        );

    \I__10034\ : LocalMux
    port map (
            O => \N__42736\,
            I => n10148
        );

    \I__10033\ : CascadeMux
    port map (
            O => \N__42731\,
            I => \N__42728\
        );

    \I__10032\ : InMux
    port map (
            O => \N__42728\,
            I => \N__42723\
        );

    \I__10031\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42718\
        );

    \I__10030\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42718\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__42723\,
            I => \N__42713\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__42718\,
            I => \N__42713\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__42713\,
            I => \N__42710\
        );

    \I__10026\ : Odrv4
    port map (
            O => \N__42710\,
            I => n7
        );

    \I__10025\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42703\
        );

    \I__10024\ : InMux
    port map (
            O => \N__42706\,
            I => \N__42700\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__42703\,
            I => \comm_state_3_N_418_1\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__42700\,
            I => \comm_state_3_N_418_1\
        );

    \I__10021\ : CascadeMux
    port map (
            O => \N__42695\,
            I => \n15711_cascade_\
        );

    \I__10020\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42689\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__42689\,
            I => n8_adj_1193
        );

    \I__10018\ : InMux
    port map (
            O => \N__42686\,
            I => \N__42683\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__42683\,
            I => \N__42680\
        );

    \I__10016\ : Span4Mux_h
    port map (
            O => \N__42680\,
            I => \N__42677\
        );

    \I__10015\ : Odrv4
    port map (
            O => \N__42677\,
            I => buf_data2_9
        );

    \I__10014\ : CascadeMux
    port map (
            O => \N__42674\,
            I => \N__42671\
        );

    \I__10013\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42667\
        );

    \I__10012\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42664\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__42667\,
            I => \N__42661\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__42664\,
            I => \N__42658\
        );

    \I__10009\ : Span4Mux_v
    port map (
            O => \N__42661\,
            I => \N__42653\
        );

    \I__10008\ : Span4Mux_h
    port map (
            O => \N__42658\,
            I => \N__42653\
        );

    \I__10007\ : Span4Mux_v
    port map (
            O => \N__42653\,
            I => \N__42649\
        );

    \I__10006\ : CascadeMux
    port map (
            O => \N__42652\,
            I => \N__42646\
        );

    \I__10005\ : Sp12to4
    port map (
            O => \N__42649\,
            I => \N__42643\
        );

    \I__10004\ : InMux
    port map (
            O => \N__42646\,
            I => \N__42640\
        );

    \I__10003\ : Span12Mux_h
    port map (
            O => \N__42643\,
            I => \N__42637\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__42640\,
            I => buf_adcdata4_9
        );

    \I__10001\ : Odrv12
    port map (
            O => \N__42637\,
            I => buf_adcdata4_9
        );

    \I__10000\ : InMux
    port map (
            O => \N__42632\,
            I => \N__42629\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42626\
        );

    \I__9998\ : Span12Mux_h
    port map (
            O => \N__42626\,
            I => \N__42623\
        );

    \I__9997\ : Odrv12
    port map (
            O => \N__42623\,
            I => n4063
        );

    \I__9996\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42617\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__42617\,
            I => \N__42613\
        );

    \I__9994\ : InMux
    port map (
            O => \N__42616\,
            I => \N__42610\
        );

    \I__9993\ : Span4Mux_h
    port map (
            O => \N__42613\,
            I => \N__42607\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__42610\,
            I => buf_adcdata2_11
        );

    \I__9991\ : Odrv4
    port map (
            O => \N__42607\,
            I => buf_adcdata2_11
        );

    \I__9990\ : InMux
    port map (
            O => \N__42602\,
            I => \N__42598\
        );

    \I__9989\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42595\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__42598\,
            I => \N__42592\
        );

    \I__9987\ : LocalMux
    port map (
            O => \N__42595\,
            I => \N__42589\
        );

    \I__9986\ : Span4Mux_v
    port map (
            O => \N__42592\,
            I => \N__42586\
        );

    \I__9985\ : Odrv4
    port map (
            O => \N__42589\,
            I => n8_adj_1219
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__42586\,
            I => n8_adj_1219
        );

    \I__9983\ : InMux
    port map (
            O => \N__42581\,
            I => \N__42577\
        );

    \I__9982\ : InMux
    port map (
            O => \N__42580\,
            I => \N__42574\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__42577\,
            I => \N__42571\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__42574\,
            I => \N__42566\
        );

    \I__9979\ : Span4Mux_h
    port map (
            O => \N__42571\,
            I => \N__42566\
        );

    \I__9978\ : Odrv4
    port map (
            O => \N__42566\,
            I => n7_adj_1218
        );

    \I__9977\ : CascadeMux
    port map (
            O => \N__42563\,
            I => \N__42560\
        );

    \I__9976\ : CascadeBuf
    port map (
            O => \N__42560\,
            I => \N__42557\
        );

    \I__9975\ : CascadeMux
    port map (
            O => \N__42557\,
            I => \N__42554\
        );

    \I__9974\ : CascadeBuf
    port map (
            O => \N__42554\,
            I => \N__42551\
        );

    \I__9973\ : CascadeMux
    port map (
            O => \N__42551\,
            I => \N__42548\
        );

    \I__9972\ : CascadeBuf
    port map (
            O => \N__42548\,
            I => \N__42545\
        );

    \I__9971\ : CascadeMux
    port map (
            O => \N__42545\,
            I => \N__42542\
        );

    \I__9970\ : CascadeBuf
    port map (
            O => \N__42542\,
            I => \N__42539\
        );

    \I__9969\ : CascadeMux
    port map (
            O => \N__42539\,
            I => \N__42536\
        );

    \I__9968\ : CascadeBuf
    port map (
            O => \N__42536\,
            I => \N__42533\
        );

    \I__9967\ : CascadeMux
    port map (
            O => \N__42533\,
            I => \N__42530\
        );

    \I__9966\ : CascadeBuf
    port map (
            O => \N__42530\,
            I => \N__42527\
        );

    \I__9965\ : CascadeMux
    port map (
            O => \N__42527\,
            I => \N__42524\
        );

    \I__9964\ : CascadeBuf
    port map (
            O => \N__42524\,
            I => \N__42520\
        );

    \I__9963\ : CascadeMux
    port map (
            O => \N__42523\,
            I => \N__42517\
        );

    \I__9962\ : CascadeMux
    port map (
            O => \N__42520\,
            I => \N__42514\
        );

    \I__9961\ : CascadeBuf
    port map (
            O => \N__42517\,
            I => \N__42511\
        );

    \I__9960\ : CascadeBuf
    port map (
            O => \N__42514\,
            I => \N__42508\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__42511\,
            I => \N__42505\
        );

    \I__9958\ : CascadeMux
    port map (
            O => \N__42508\,
            I => \N__42502\
        );

    \I__9957\ : InMux
    port map (
            O => \N__42505\,
            I => \N__42499\
        );

    \I__9956\ : CascadeBuf
    port map (
            O => \N__42502\,
            I => \N__42496\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__42499\,
            I => \N__42493\
        );

    \I__9954\ : CascadeMux
    port map (
            O => \N__42496\,
            I => \N__42490\
        );

    \I__9953\ : Span12Mux_h
    port map (
            O => \N__42493\,
            I => \N__42487\
        );

    \I__9952\ : InMux
    port map (
            O => \N__42490\,
            I => \N__42484\
        );

    \I__9951\ : Span12Mux_v
    port map (
            O => \N__42487\,
            I => \N__42481\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__42484\,
            I => \N__42478\
        );

    \I__9949\ : Odrv12
    port map (
            O => \N__42481\,
            I => \data_index_9_N_258_8\
        );

    \I__9948\ : Odrv4
    port map (
            O => \N__42478\,
            I => \data_index_9_N_258_8\
        );

    \I__9947\ : InMux
    port map (
            O => \N__42473\,
            I => \N__42470\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__42470\,
            I => \comm_spi.n10456\
        );

    \I__9945\ : ClkMux
    port map (
            O => \N__42467\,
            I => \N__42456\
        );

    \I__9944\ : ClkMux
    port map (
            O => \N__42466\,
            I => \N__42452\
        );

    \I__9943\ : ClkMux
    port map (
            O => \N__42465\,
            I => \N__42449\
        );

    \I__9942\ : ClkMux
    port map (
            O => \N__42464\,
            I => \N__42444\
        );

    \I__9941\ : ClkMux
    port map (
            O => \N__42463\,
            I => \N__42441\
        );

    \I__9940\ : ClkMux
    port map (
            O => \N__42462\,
            I => \N__42435\
        );

    \I__9939\ : ClkMux
    port map (
            O => \N__42461\,
            I => \N__42432\
        );

    \I__9938\ : ClkMux
    port map (
            O => \N__42460\,
            I => \N__42428\
        );

    \I__9937\ : ClkMux
    port map (
            O => \N__42459\,
            I => \N__42425\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__42456\,
            I => \N__42421\
        );

    \I__9935\ : ClkMux
    port map (
            O => \N__42455\,
            I => \N__42417\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__42452\,
            I => \N__42414\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__42449\,
            I => \N__42411\
        );

    \I__9932\ : ClkMux
    port map (
            O => \N__42448\,
            I => \N__42408\
        );

    \I__9931\ : ClkMux
    port map (
            O => \N__42447\,
            I => \N__42405\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__42444\,
            I => \N__42399\
        );

    \I__9929\ : LocalMux
    port map (
            O => \N__42441\,
            I => \N__42399\
        );

    \I__9928\ : ClkMux
    port map (
            O => \N__42440\,
            I => \N__42396\
        );

    \I__9927\ : ClkMux
    port map (
            O => \N__42439\,
            I => \N__42393\
        );

    \I__9926\ : ClkMux
    port map (
            O => \N__42438\,
            I => \N__42390\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__42435\,
            I => \N__42385\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__42432\,
            I => \N__42385\
        );

    \I__9923\ : ClkMux
    port map (
            O => \N__42431\,
            I => \N__42382\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__42428\,
            I => \N__42376\
        );

    \I__9921\ : LocalMux
    port map (
            O => \N__42425\,
            I => \N__42376\
        );

    \I__9920\ : ClkMux
    port map (
            O => \N__42424\,
            I => \N__42372\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__42421\,
            I => \N__42368\
        );

    \I__9918\ : ClkMux
    port map (
            O => \N__42420\,
            I => \N__42365\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__42417\,
            I => \N__42362\
        );

    \I__9916\ : Span4Mux_h
    port map (
            O => \N__42414\,
            I => \N__42353\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__42411\,
            I => \N__42353\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__42408\,
            I => \N__42353\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__42405\,
            I => \N__42353\
        );

    \I__9912\ : ClkMux
    port map (
            O => \N__42404\,
            I => \N__42350\
        );

    \I__9911\ : Span4Mux_v
    port map (
            O => \N__42399\,
            I => \N__42345\
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__42396\,
            I => \N__42345\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__42393\,
            I => \N__42342\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__42390\,
            I => \N__42339\
        );

    \I__9907\ : Span4Mux_v
    port map (
            O => \N__42385\,
            I => \N__42334\
        );

    \I__9906\ : LocalMux
    port map (
            O => \N__42382\,
            I => \N__42334\
        );

    \I__9905\ : ClkMux
    port map (
            O => \N__42381\,
            I => \N__42331\
        );

    \I__9904\ : Span4Mux_v
    port map (
            O => \N__42376\,
            I => \N__42328\
        );

    \I__9903\ : ClkMux
    port map (
            O => \N__42375\,
            I => \N__42325\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__42372\,
            I => \N__42322\
        );

    \I__9901\ : ClkMux
    port map (
            O => \N__42371\,
            I => \N__42319\
        );

    \I__9900\ : Span4Mux_h
    port map (
            O => \N__42368\,
            I => \N__42314\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__42365\,
            I => \N__42314\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__42362\,
            I => \N__42307\
        );

    \I__9897\ : Span4Mux_h
    port map (
            O => \N__42353\,
            I => \N__42307\
        );

    \I__9896\ : LocalMux
    port map (
            O => \N__42350\,
            I => \N__42307\
        );

    \I__9895\ : Span4Mux_v
    port map (
            O => \N__42345\,
            I => \N__42302\
        );

    \I__9894\ : Span4Mux_v
    port map (
            O => \N__42342\,
            I => \N__42302\
        );

    \I__9893\ : Span4Mux_h
    port map (
            O => \N__42339\,
            I => \N__42299\
        );

    \I__9892\ : Span4Mux_h
    port map (
            O => \N__42334\,
            I => \N__42294\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42294\
        );

    \I__9890\ : Span4Mux_h
    port map (
            O => \N__42328\,
            I => \N__42285\
        );

    \I__9889\ : LocalMux
    port map (
            O => \N__42325\,
            I => \N__42285\
        );

    \I__9888\ : Span4Mux_v
    port map (
            O => \N__42322\,
            I => \N__42285\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__42319\,
            I => \N__42285\
        );

    \I__9886\ : Span4Mux_h
    port map (
            O => \N__42314\,
            I => \N__42280\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__42307\,
            I => \N__42280\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__42302\,
            I => \N__42277\
        );

    \I__9883\ : Span4Mux_v
    port map (
            O => \N__42299\,
            I => \N__42272\
        );

    \I__9882\ : Span4Mux_h
    port map (
            O => \N__42294\,
            I => \N__42272\
        );

    \I__9881\ : Span4Mux_h
    port map (
            O => \N__42285\,
            I => \N__42269\
        );

    \I__9880\ : Odrv4
    port map (
            O => \N__42280\,
            I => \comm_spi.iclk\
        );

    \I__9879\ : Odrv4
    port map (
            O => \N__42277\,
            I => \comm_spi.iclk\
        );

    \I__9878\ : Odrv4
    port map (
            O => \N__42272\,
            I => \comm_spi.iclk\
        );

    \I__9877\ : Odrv4
    port map (
            O => \N__42269\,
            I => \comm_spi.iclk\
        );

    \I__9876\ : InMux
    port map (
            O => \N__42260\,
            I => \N__42257\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__42257\,
            I => \N__42254\
        );

    \I__9874\ : Span4Mux_v
    port map (
            O => \N__42254\,
            I => \N__42249\
        );

    \I__9873\ : InMux
    port map (
            O => \N__42253\,
            I => \N__42246\
        );

    \I__9872\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42243\
        );

    \I__9871\ : Odrv4
    port map (
            O => \N__42249\,
            I => \comm_spi.n16893\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__42246\,
            I => \comm_spi.n16893\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__42243\,
            I => \comm_spi.n16893\
        );

    \I__9868\ : InMux
    port map (
            O => \N__42236\,
            I => \N__42233\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__42233\,
            I => \N__42229\
        );

    \I__9866\ : InMux
    port map (
            O => \N__42232\,
            I => \N__42225\
        );

    \I__9865\ : Span4Mux_v
    port map (
            O => \N__42229\,
            I => \N__42222\
        );

    \I__9864\ : InMux
    port map (
            O => \N__42228\,
            I => \N__42219\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__42225\,
            I => \N__42216\
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__42222\,
            I => \comm_spi.n10441\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__42219\,
            I => \comm_spi.n10441\
        );

    \I__9860\ : Odrv4
    port map (
            O => \N__42216\,
            I => \comm_spi.n10441\
        );

    \I__9859\ : CascadeMux
    port map (
            O => \N__42209\,
            I => \comm_spi.n16893_cascade_\
        );

    \I__9858\ : CascadeMux
    port map (
            O => \N__42206\,
            I => \comm_spi.imosi_cascade_\
        );

    \I__9857\ : SRMux
    port map (
            O => \N__42203\,
            I => \N__42200\
        );

    \I__9856\ : LocalMux
    port map (
            O => \N__42200\,
            I => \N__42197\
        );

    \I__9855\ : Span4Mux_h
    port map (
            O => \N__42197\,
            I => \N__42194\
        );

    \I__9854\ : Odrv4
    port map (
            O => \N__42194\,
            I => \comm_spi.DOUT_7__N_785\
        );

    \I__9853\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42188\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__42188\,
            I => \N__42184\
        );

    \I__9851\ : CascadeMux
    port map (
            O => \N__42187\,
            I => \N__42181\
        );

    \I__9850\ : Span4Mux_v
    port map (
            O => \N__42184\,
            I => \N__42178\
        );

    \I__9849\ : InMux
    port map (
            O => \N__42181\,
            I => \N__42174\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__42178\,
            I => \N__42171\
        );

    \I__9847\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42168\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__42174\,
            I => \acadc_skipCount_1\
        );

    \I__9845\ : Odrv4
    port map (
            O => \N__42171\,
            I => \acadc_skipCount_1\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__42168\,
            I => \acadc_skipCount_1\
        );

    \I__9843\ : InMux
    port map (
            O => \N__42161\,
            I => \N__42156\
        );

    \I__9842\ : InMux
    port map (
            O => \N__42160\,
            I => \N__42153\
        );

    \I__9841\ : InMux
    port map (
            O => \N__42159\,
            I => \N__42150\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__42156\,
            I => req_data_cnt_1
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__42153\,
            I => req_data_cnt_1
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__42150\,
            I => req_data_cnt_1
        );

    \I__9837\ : CascadeMux
    port map (
            O => \N__42143\,
            I => \n4220_cascade_\
        );

    \I__9836\ : CascadeMux
    port map (
            O => \N__42140\,
            I => \n4253_cascade_\
        );

    \I__9835\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42134\
        );

    \I__9834\ : LocalMux
    port map (
            O => \N__42134\,
            I => \N__42131\
        );

    \I__9833\ : Span12Mux_v
    port map (
            O => \N__42131\,
            I => \N__42128\
        );

    \I__9832\ : Odrv12
    port map (
            O => \N__42128\,
            I => n4263
        );

    \I__9831\ : InMux
    port map (
            O => \N__42125\,
            I => \N__42121\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__42124\,
            I => \N__42117\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__42121\,
            I => \N__42114\
        );

    \I__9828\ : InMux
    port map (
            O => \N__42120\,
            I => \N__42111\
        );

    \I__9827\ : InMux
    port map (
            O => \N__42117\,
            I => \N__42108\
        );

    \I__9826\ : Span4Mux_v
    port map (
            O => \N__42114\,
            I => \N__42105\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__42111\,
            I => \N__42102\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__42108\,
            I => buf_dds_1
        );

    \I__9823\ : Odrv4
    port map (
            O => \N__42105\,
            I => buf_dds_1
        );

    \I__9822\ : Odrv12
    port map (
            O => \N__42102\,
            I => buf_dds_1
        );

    \I__9821\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42092\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__42092\,
            I => \N__42089\
        );

    \I__9819\ : Span4Mux_v
    port map (
            O => \N__42089\,
            I => \N__42084\
        );

    \I__9818\ : InMux
    port map (
            O => \N__42088\,
            I => \N__42081\
        );

    \I__9817\ : InMux
    port map (
            O => \N__42087\,
            I => \N__42078\
        );

    \I__9816\ : Sp12to4
    port map (
            O => \N__42084\,
            I => \N__42073\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__42081\,
            I => \N__42073\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__42078\,
            I => buf_adcdata3_9
        );

    \I__9813\ : Odrv12
    port map (
            O => \N__42073\,
            I => buf_adcdata3_9
        );

    \I__9812\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42065\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__42065\,
            I => n4208
        );

    \I__9810\ : CascadeMux
    port map (
            O => \N__42062\,
            I => \N__42059\
        );

    \I__9809\ : InMux
    port map (
            O => \N__42059\,
            I => \N__42056\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__42056\,
            I => \N__42053\
        );

    \I__9807\ : Span4Mux_h
    port map (
            O => \N__42053\,
            I => \N__42050\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__42050\,
            I => buf_data1_9
        );

    \I__9805\ : InMux
    port map (
            O => \N__42047\,
            I => \N__42044\
        );

    \I__9804\ : LocalMux
    port map (
            O => \N__42044\,
            I => n4196
        );

    \I__9803\ : InMux
    port map (
            O => \N__42041\,
            I => \N__42038\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__42038\,
            I => n4233
        );

    \I__9801\ : InMux
    port map (
            O => \N__42035\,
            I => \N__42032\
        );

    \I__9800\ : LocalMux
    port map (
            O => \N__42032\,
            I => \N__42028\
        );

    \I__9799\ : InMux
    port map (
            O => \N__42031\,
            I => \N__42025\
        );

    \I__9798\ : Span4Mux_v
    port map (
            O => \N__42028\,
            I => \N__42022\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__42025\,
            I => data_idxvec_3
        );

    \I__9796\ : Odrv4
    port map (
            O => \N__42022\,
            I => data_idxvec_3
        );

    \I__9795\ : InMux
    port map (
            O => \N__42017\,
            I => \N__42012\
        );

    \I__9794\ : InMux
    port map (
            O => \N__42016\,
            I => \N__42009\
        );

    \I__9793\ : InMux
    port map (
            O => \N__42015\,
            I => \N__42006\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__42012\,
            I => \N__42003\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__42009\,
            I => data_cntvec_3
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__42006\,
            I => data_cntvec_3
        );

    \I__9789\ : Odrv4
    port map (
            O => \N__42003\,
            I => data_cntvec_3
        );

    \I__9788\ : InMux
    port map (
            O => \N__41996\,
            I => \N__41993\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__41993\,
            I => \N__41990\
        );

    \I__9786\ : Span4Mux_v
    port map (
            O => \N__41990\,
            I => \N__41987\
        );

    \I__9785\ : Span4Mux_h
    port map (
            O => \N__41987\,
            I => \N__41984\
        );

    \I__9784\ : Odrv4
    port map (
            O => \N__41984\,
            I => buf_data1_11
        );

    \I__9783\ : CascadeMux
    port map (
            O => \N__41981\,
            I => \n4194_cascade_\
        );

    \I__9782\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41975\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__41975\,
            I => n4218
        );

    \I__9780\ : CascadeMux
    port map (
            O => \N__41972\,
            I => \n4231_cascade_\
        );

    \I__9779\ : InMux
    port map (
            O => \N__41969\,
            I => \N__41966\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__41966\,
            I => \N__41963\
        );

    \I__9777\ : Odrv4
    port map (
            O => \N__41963\,
            I => n4206
        );

    \I__9776\ : CascadeMux
    port map (
            O => \N__41960\,
            I => \n4251_cascade_\
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__41957\,
            I => \N__41953\
        );

    \I__9774\ : CascadeMux
    port map (
            O => \N__41956\,
            I => \N__41950\
        );

    \I__9773\ : InMux
    port map (
            O => \N__41953\,
            I => \N__41944\
        );

    \I__9772\ : InMux
    port map (
            O => \N__41950\,
            I => \N__41944\
        );

    \I__9771\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41941\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__41944\,
            I => cmd_rdadctmp_21_adj_1091
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__41941\,
            I => cmd_rdadctmp_21_adj_1091
        );

    \I__9768\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41932\
        );

    \I__9767\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41928\
        );

    \I__9766\ : LocalMux
    port map (
            O => \N__41932\,
            I => \N__41925\
        );

    \I__9765\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41922\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41919\
        );

    \I__9763\ : Span4Mux_v
    port map (
            O => \N__41925\,
            I => \N__41914\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__41922\,
            I => \N__41914\
        );

    \I__9761\ : Span4Mux_v
    port map (
            O => \N__41919\,
            I => \N__41910\
        );

    \I__9760\ : Span4Mux_h
    port map (
            O => \N__41914\,
            I => \N__41907\
        );

    \I__9759\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41904\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__41910\,
            I => n4_adj_1041
        );

    \I__9757\ : Odrv4
    port map (
            O => \N__41907\,
            I => n4_adj_1041
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__41904\,
            I => n4_adj_1041
        );

    \I__9755\ : CascadeMux
    port map (
            O => \N__41897\,
            I => \N__41891\
        );

    \I__9754\ : InMux
    port map (
            O => \N__41896\,
            I => \N__41888\
        );

    \I__9753\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41883\
        );

    \I__9752\ : InMux
    port map (
            O => \N__41894\,
            I => \N__41880\
        );

    \I__9751\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41877\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__41888\,
            I => \N__41874\
        );

    \I__9749\ : InMux
    port map (
            O => \N__41887\,
            I => \N__41869\
        );

    \I__9748\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41869\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41864\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__41880\,
            I => \N__41864\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__41877\,
            I => \N__41860\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__41874\,
            I => \N__41855\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__41869\,
            I => \N__41855\
        );

    \I__9742\ : Span4Mux_v
    port map (
            O => \N__41864\,
            I => \N__41852\
        );

    \I__9741\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41849\
        );

    \I__9740\ : Span4Mux_h
    port map (
            O => \N__41860\,
            I => \N__41846\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__41855\,
            I => \N__41843\
        );

    \I__9738\ : Sp12to4
    port map (
            O => \N__41852\,
            I => \N__41838\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__41849\,
            I => \N__41838\
        );

    \I__9736\ : Span4Mux_v
    port map (
            O => \N__41846\,
            I => \N__41835\
        );

    \I__9735\ : Odrv4
    port map (
            O => \N__41843\,
            I => comm_buf_0_6
        );

    \I__9734\ : Odrv12
    port map (
            O => \N__41838\,
            I => comm_buf_0_6
        );

    \I__9733\ : Odrv4
    port map (
            O => \N__41835\,
            I => comm_buf_0_6
        );

    \I__9732\ : CascadeMux
    port map (
            O => \N__41828\,
            I => \N__41815\
        );

    \I__9731\ : InMux
    port map (
            O => \N__41827\,
            I => \N__41812\
        );

    \I__9730\ : InMux
    port map (
            O => \N__41826\,
            I => \N__41807\
        );

    \I__9729\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41807\
        );

    \I__9728\ : InMux
    port map (
            O => \N__41824\,
            I => \N__41804\
        );

    \I__9727\ : InMux
    port map (
            O => \N__41823\,
            I => \N__41801\
        );

    \I__9726\ : InMux
    port map (
            O => \N__41822\,
            I => \N__41798\
        );

    \I__9725\ : InMux
    port map (
            O => \N__41821\,
            I => \N__41791\
        );

    \I__9724\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41791\
        );

    \I__9723\ : InMux
    port map (
            O => \N__41819\,
            I => \N__41791\
        );

    \I__9722\ : InMux
    port map (
            O => \N__41818\,
            I => \N__41786\
        );

    \I__9721\ : InMux
    port map (
            O => \N__41815\,
            I => \N__41782\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__41812\,
            I => \N__41779\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__41807\,
            I => \N__41776\
        );

    \I__9718\ : LocalMux
    port map (
            O => \N__41804\,
            I => \N__41773\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__41801\,
            I => \N__41766\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__41798\,
            I => \N__41766\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__41791\,
            I => \N__41766\
        );

    \I__9714\ : InMux
    port map (
            O => \N__41790\,
            I => \N__41761\
        );

    \I__9713\ : InMux
    port map (
            O => \N__41789\,
            I => \N__41761\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__41786\,
            I => \N__41758\
        );

    \I__9711\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41753\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__41782\,
            I => \N__41746\
        );

    \I__9709\ : Span4Mux_v
    port map (
            O => \N__41779\,
            I => \N__41746\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__41776\,
            I => \N__41746\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__41773\,
            I => \N__41739\
        );

    \I__9706\ : Span4Mux_v
    port map (
            O => \N__41766\,
            I => \N__41739\
        );

    \I__9705\ : LocalMux
    port map (
            O => \N__41761\,
            I => \N__41739\
        );

    \I__9704\ : Span4Mux_h
    port map (
            O => \N__41758\,
            I => \N__41736\
        );

    \I__9703\ : InMux
    port map (
            O => \N__41757\,
            I => \N__41733\
        );

    \I__9702\ : InMux
    port map (
            O => \N__41756\,
            I => \N__41730\
        );

    \I__9701\ : LocalMux
    port map (
            O => \N__41753\,
            I => \N__41727\
        );

    \I__9700\ : Span4Mux_h
    port map (
            O => \N__41746\,
            I => \N__41724\
        );

    \I__9699\ : Span4Mux_h
    port map (
            O => \N__41739\,
            I => \N__41719\
        );

    \I__9698\ : Span4Mux_h
    port map (
            O => \N__41736\,
            I => \N__41719\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__41733\,
            I => n8250
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__41730\,
            I => n8250
        );

    \I__9695\ : Odrv12
    port map (
            O => \N__41727\,
            I => n8250
        );

    \I__9694\ : Odrv4
    port map (
            O => \N__41724\,
            I => n8250
        );

    \I__9693\ : Odrv4
    port map (
            O => \N__41719\,
            I => n8250
        );

    \I__9692\ : InMux
    port map (
            O => \N__41708\,
            I => \N__41705\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__41705\,
            I => \N__41701\
        );

    \I__9690\ : InMux
    port map (
            O => \N__41704\,
            I => \N__41698\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__41701\,
            I => \N__41694\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__41698\,
            I => \N__41691\
        );

    \I__9687\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41688\
        );

    \I__9686\ : Span4Mux_h
    port map (
            O => \N__41694\,
            I => \N__41685\
        );

    \I__9685\ : Span4Mux_v
    port map (
            O => \N__41691\,
            I => \N__41682\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__41688\,
            I => \acadc_skipCount_14\
        );

    \I__9683\ : Odrv4
    port map (
            O => \N__41685\,
            I => \acadc_skipCount_14\
        );

    \I__9682\ : Odrv4
    port map (
            O => \N__41682\,
            I => \acadc_skipCount_14\
        );

    \I__9681\ : CascadeMux
    port map (
            O => \N__41675\,
            I => \N__41671\
        );

    \I__9680\ : CascadeMux
    port map (
            O => \N__41674\,
            I => \N__41668\
        );

    \I__9679\ : InMux
    port map (
            O => \N__41671\,
            I => \N__41665\
        );

    \I__9678\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41662\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__41665\,
            I => data_idxvec_15
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__41662\,
            I => data_idxvec_15
        );

    \I__9675\ : CascadeMux
    port map (
            O => \N__41657\,
            I => \N__41653\
        );

    \I__9674\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41649\
        );

    \I__9673\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41646\
        );

    \I__9672\ : InMux
    port map (
            O => \N__41652\,
            I => \N__41643\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__41649\,
            I => \N__41640\
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__41646\,
            I => \acadc_skipCount_15\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__41643\,
            I => \acadc_skipCount_15\
        );

    \I__9668\ : Odrv4
    port map (
            O => \N__41640\,
            I => \acadc_skipCount_15\
        );

    \I__9667\ : CascadeMux
    port map (
            O => \N__41633\,
            I => \N__41630\
        );

    \I__9666\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41627\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__41627\,
            I => \N__41624\
        );

    \I__9664\ : Span4Mux_v
    port map (
            O => \N__41624\,
            I => \N__41621\
        );

    \I__9663\ : Span4Mux_h
    port map (
            O => \N__41621\,
            I => \N__41618\
        );

    \I__9662\ : Odrv4
    port map (
            O => \N__41618\,
            I => n15468
        );

    \I__9661\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41612\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__41612\,
            I => \N__41609\
        );

    \I__9659\ : Odrv4
    port map (
            O => \N__41609\,
            I => n4217
        );

    \I__9658\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41603\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__41603\,
            I => n4230
        );

    \I__9656\ : InMux
    port map (
            O => \N__41600\,
            I => \N__41597\
        );

    \I__9655\ : LocalMux
    port map (
            O => \N__41597\,
            I => \N__41594\
        );

    \I__9654\ : Span4Mux_h
    port map (
            O => \N__41594\,
            I => \N__41591\
        );

    \I__9653\ : Span4Mux_v
    port map (
            O => \N__41591\,
            I => \N__41588\
        );

    \I__9652\ : Odrv4
    port map (
            O => \N__41588\,
            I => n4250
        );

    \I__9651\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41582\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__41582\,
            I => \N__41579\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__41579\,
            I => \N__41575\
        );

    \I__9648\ : InMux
    port map (
            O => \N__41578\,
            I => \N__41571\
        );

    \I__9647\ : Span4Mux_h
    port map (
            O => \N__41575\,
            I => \N__41568\
        );

    \I__9646\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41565\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__41571\,
            I => cmd_rdadctmp_22_adj_1090
        );

    \I__9644\ : Odrv4
    port map (
            O => \N__41568\,
            I => cmd_rdadctmp_22_adj_1090
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__41565\,
            I => cmd_rdadctmp_22_adj_1090
        );

    \I__9642\ : InMux
    port map (
            O => \N__41558\,
            I => \N__41554\
        );

    \I__9641\ : InMux
    port map (
            O => \N__41557\,
            I => \N__41551\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__41554\,
            I => \N__41547\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__41551\,
            I => \N__41544\
        );

    \I__9638\ : InMux
    port map (
            O => \N__41550\,
            I => \N__41541\
        );

    \I__9637\ : Span4Mux_v
    port map (
            O => \N__41547\,
            I => \N__41538\
        );

    \I__9636\ : Span4Mux_v
    port map (
            O => \N__41544\,
            I => \N__41535\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__41541\,
            I => buf_adcdata3_14
        );

    \I__9634\ : Odrv4
    port map (
            O => \N__41538\,
            I => buf_adcdata3_14
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__41535\,
            I => buf_adcdata3_14
        );

    \I__9632\ : CascadeMux
    port map (
            O => \N__41528\,
            I => \N__41521\
        );

    \I__9631\ : CascadeMux
    port map (
            O => \N__41527\,
            I => \N__41515\
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__41526\,
            I => \N__41512\
        );

    \I__9629\ : InMux
    port map (
            O => \N__41525\,
            I => \N__41507\
        );

    \I__9628\ : InMux
    port map (
            O => \N__41524\,
            I => \N__41502\
        );

    \I__9627\ : InMux
    port map (
            O => \N__41521\,
            I => \N__41499\
        );

    \I__9626\ : CascadeMux
    port map (
            O => \N__41520\,
            I => \N__41494\
        );

    \I__9625\ : CascadeMux
    port map (
            O => \N__41519\,
            I => \N__41491\
        );

    \I__9624\ : CascadeMux
    port map (
            O => \N__41518\,
            I => \N__41488\
        );

    \I__9623\ : InMux
    port map (
            O => \N__41515\,
            I => \N__41485\
        );

    \I__9622\ : InMux
    port map (
            O => \N__41512\,
            I => \N__41482\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__41511\,
            I => \N__41479\
        );

    \I__9620\ : InMux
    port map (
            O => \N__41510\,
            I => \N__41476\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__41507\,
            I => \N__41473\
        );

    \I__9618\ : CascadeMux
    port map (
            O => \N__41506\,
            I => \N__41470\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__41505\,
            I => \N__41467\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__41502\,
            I => \N__41464\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__41499\,
            I => \N__41461\
        );

    \I__9614\ : InMux
    port map (
            O => \N__41498\,
            I => \N__41454\
        );

    \I__9613\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41454\
        );

    \I__9612\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41454\
        );

    \I__9611\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41451\
        );

    \I__9610\ : InMux
    port map (
            O => \N__41488\,
            I => \N__41448\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__41485\,
            I => \N__41443\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__41482\,
            I => \N__41443\
        );

    \I__9607\ : InMux
    port map (
            O => \N__41479\,
            I => \N__41440\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__41476\,
            I => \N__41437\
        );

    \I__9605\ : Span4Mux_h
    port map (
            O => \N__41473\,
            I => \N__41434\
        );

    \I__9604\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41429\
        );

    \I__9603\ : InMux
    port map (
            O => \N__41467\,
            I => \N__41429\
        );

    \I__9602\ : Span4Mux_v
    port map (
            O => \N__41464\,
            I => \N__41426\
        );

    \I__9601\ : Span4Mux_v
    port map (
            O => \N__41461\,
            I => \N__41423\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__41454\,
            I => \N__41420\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__41451\,
            I => \N__41417\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41404\
        );

    \I__9597\ : Span4Mux_h
    port map (
            O => \N__41443\,
            I => \N__41404\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__41440\,
            I => \N__41404\
        );

    \I__9595\ : Span4Mux_v
    port map (
            O => \N__41437\,
            I => \N__41404\
        );

    \I__9594\ : Span4Mux_h
    port map (
            O => \N__41434\,
            I => \N__41404\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__41429\,
            I => \N__41404\
        );

    \I__9592\ : Span4Mux_h
    port map (
            O => \N__41426\,
            I => \N__41399\
        );

    \I__9591\ : Span4Mux_h
    port map (
            O => \N__41423\,
            I => \N__41399\
        );

    \I__9590\ : Span4Mux_v
    port map (
            O => \N__41420\,
            I => \N__41396\
        );

    \I__9589\ : Span4Mux_h
    port map (
            O => \N__41417\,
            I => \N__41391\
        );

    \I__9588\ : Span4Mux_v
    port map (
            O => \N__41404\,
            I => \N__41391\
        );

    \I__9587\ : Span4Mux_v
    port map (
            O => \N__41399\,
            I => \N__41388\
        );

    \I__9586\ : Odrv4
    port map (
            O => \N__41396\,
            I => n1
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__41391\,
            I => n1
        );

    \I__9584\ : Odrv4
    port map (
            O => \N__41388\,
            I => n1
        );

    \I__9583\ : CascadeMux
    port map (
            O => \N__41381\,
            I => \N__41375\
        );

    \I__9582\ : InMux
    port map (
            O => \N__41380\,
            I => \N__41370\
        );

    \I__9581\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41365\
        );

    \I__9580\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41362\
        );

    \I__9579\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41357\
        );

    \I__9578\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41353\
        );

    \I__9577\ : InMux
    port map (
            O => \N__41373\,
            I => \N__41350\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__41370\,
            I => \N__41347\
        );

    \I__9575\ : InMux
    port map (
            O => \N__41369\,
            I => \N__41343\
        );

    \I__9574\ : InMux
    port map (
            O => \N__41368\,
            I => \N__41340\
        );

    \I__9573\ : LocalMux
    port map (
            O => \N__41365\,
            I => \N__41337\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__41362\,
            I => \N__41334\
        );

    \I__9571\ : InMux
    port map (
            O => \N__41361\,
            I => \N__41329\
        );

    \I__9570\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41329\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__41357\,
            I => \N__41326\
        );

    \I__9568\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41323\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__41353\,
            I => \N__41320\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__41350\,
            I => \N__41315\
        );

    \I__9565\ : Span4Mux_h
    port map (
            O => \N__41347\,
            I => \N__41315\
        );

    \I__9564\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41309\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__41343\,
            I => \N__41306\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__41340\,
            I => \N__41301\
        );

    \I__9561\ : Span4Mux_v
    port map (
            O => \N__41337\,
            I => \N__41301\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__41334\,
            I => \N__41288\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__41329\,
            I => \N__41288\
        );

    \I__9558\ : Span4Mux_h
    port map (
            O => \N__41326\,
            I => \N__41288\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__41323\,
            I => \N__41288\
        );

    \I__9556\ : Span4Mux_v
    port map (
            O => \N__41320\,
            I => \N__41288\
        );

    \I__9555\ : Span4Mux_h
    port map (
            O => \N__41315\,
            I => \N__41288\
        );

    \I__9554\ : InMux
    port map (
            O => \N__41314\,
            I => \N__41285\
        );

    \I__9553\ : InMux
    port map (
            O => \N__41313\,
            I => \N__41280\
        );

    \I__9552\ : InMux
    port map (
            O => \N__41312\,
            I => \N__41280\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__41309\,
            I => \N__41277\
        );

    \I__9550\ : Span4Mux_v
    port map (
            O => \N__41306\,
            I => \N__41272\
        );

    \I__9549\ : Span4Mux_v
    port map (
            O => \N__41301\,
            I => \N__41272\
        );

    \I__9548\ : Span4Mux_v
    port map (
            O => \N__41288\,
            I => \N__41269\
        );

    \I__9547\ : LocalMux
    port map (
            O => \N__41285\,
            I => n8525
        );

    \I__9546\ : LocalMux
    port map (
            O => \N__41280\,
            I => n8525
        );

    \I__9545\ : Odrv4
    port map (
            O => \N__41277\,
            I => n8525
        );

    \I__9544\ : Odrv4
    port map (
            O => \N__41272\,
            I => n8525
        );

    \I__9543\ : Odrv4
    port map (
            O => \N__41269\,
            I => n8525
        );

    \I__9542\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41254\
        );

    \I__9541\ : InMux
    port map (
            O => \N__41257\,
            I => \N__41251\
        );

    \I__9540\ : LocalMux
    port map (
            O => \N__41254\,
            I => \N__41248\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__41251\,
            I => \N__41245\
        );

    \I__9538\ : Span4Mux_v
    port map (
            O => \N__41248\,
            I => \N__41242\
        );

    \I__9537\ : Span4Mux_h
    port map (
            O => \N__41245\,
            I => \N__41238\
        );

    \I__9536\ : Span4Mux_h
    port map (
            O => \N__41242\,
            I => \N__41235\
        );

    \I__9535\ : InMux
    port map (
            O => \N__41241\,
            I => \N__41232\
        );

    \I__9534\ : Span4Mux_v
    port map (
            O => \N__41238\,
            I => \N__41227\
        );

    \I__9533\ : Span4Mux_h
    port map (
            O => \N__41235\,
            I => \N__41227\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__41232\,
            I => buf_dds_11
        );

    \I__9531\ : Odrv4
    port map (
            O => \N__41227\,
            I => buf_dds_11
        );

    \I__9530\ : CascadeMux
    port map (
            O => \N__41222\,
            I => \N__41218\
        );

    \I__9529\ : InMux
    port map (
            O => \N__41221\,
            I => \N__41215\
        );

    \I__9528\ : InMux
    port map (
            O => \N__41218\,
            I => \N__41212\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__41215\,
            I => \N__41207\
        );

    \I__9526\ : LocalMux
    port map (
            O => \N__41212\,
            I => \N__41204\
        );

    \I__9525\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41201\
        );

    \I__9524\ : InMux
    port map (
            O => \N__41210\,
            I => \N__41197\
        );

    \I__9523\ : Span4Mux_h
    port map (
            O => \N__41207\,
            I => \N__41190\
        );

    \I__9522\ : Span4Mux_v
    port map (
            O => \N__41204\,
            I => \N__41190\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__41201\,
            I => \N__41190\
        );

    \I__9520\ : InMux
    port map (
            O => \N__41200\,
            I => \N__41187\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__41197\,
            I => n12
        );

    \I__9518\ : Odrv4
    port map (
            O => \N__41190\,
            I => n12
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__41187\,
            I => n12
        );

    \I__9516\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41177\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__41177\,
            I => \N__41174\
        );

    \I__9514\ : Odrv4
    port map (
            O => \N__41174\,
            I => n13_adj_1025
        );

    \I__9513\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41161\
        );

    \I__9512\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41161\
        );

    \I__9511\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41158\
        );

    \I__9510\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41155\
        );

    \I__9509\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41152\
        );

    \I__9508\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41148\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__41161\,
            I => \N__41139\
        );

    \I__9506\ : LocalMux
    port map (
            O => \N__41158\,
            I => \N__41139\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__41155\,
            I => \N__41139\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__41152\,
            I => \N__41139\
        );

    \I__9503\ : InMux
    port map (
            O => \N__41151\,
            I => \N__41136\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__41148\,
            I => \N__41133\
        );

    \I__9501\ : Span4Mux_v
    port map (
            O => \N__41139\,
            I => \N__41130\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__41136\,
            I => \N__41127\
        );

    \I__9499\ : Span12Mux_v
    port map (
            O => \N__41133\,
            I => \N__41123\
        );

    \I__9498\ : Span4Mux_h
    port map (
            O => \N__41130\,
            I => \N__41120\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__41127\,
            I => \N__41117\
        );

    \I__9496\ : InMux
    port map (
            O => \N__41126\,
            I => \N__41114\
        );

    \I__9495\ : Odrv12
    port map (
            O => \N__41123\,
            I => n7511
        );

    \I__9494\ : Odrv4
    port map (
            O => \N__41120\,
            I => n7511
        );

    \I__9493\ : Odrv4
    port map (
            O => \N__41117\,
            I => n7511
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__41114\,
            I => n7511
        );

    \I__9491\ : InMux
    port map (
            O => \N__41105\,
            I => \N__41102\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__41102\,
            I => \N__41098\
        );

    \I__9489\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41093\
        );

    \I__9488\ : Span4Mux_v
    port map (
            O => \N__41098\,
            I => \N__41089\
        );

    \I__9487\ : InMux
    port map (
            O => \N__41097\,
            I => \N__41086\
        );

    \I__9486\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41083\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__41093\,
            I => \N__41080\
        );

    \I__9484\ : InMux
    port map (
            O => \N__41092\,
            I => \N__41077\
        );

    \I__9483\ : Span4Mux_h
    port map (
            O => \N__41089\,
            I => \N__41074\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__41086\,
            I => \N__41071\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__41083\,
            I => \N__41068\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__41080\,
            I => \N__41063\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__41077\,
            I => \N__41063\
        );

    \I__9478\ : Span4Mux_h
    port map (
            O => \N__41074\,
            I => \N__41060\
        );

    \I__9477\ : Span4Mux_h
    port map (
            O => \N__41071\,
            I => \N__41055\
        );

    \I__9476\ : Span4Mux_h
    port map (
            O => \N__41068\,
            I => \N__41055\
        );

    \I__9475\ : Span4Mux_h
    port map (
            O => \N__41063\,
            I => \N__41052\
        );

    \I__9474\ : Odrv4
    port map (
            O => \N__41060\,
            I => comm_buf_1_1
        );

    \I__9473\ : Odrv4
    port map (
            O => \N__41055\,
            I => comm_buf_1_1
        );

    \I__9472\ : Odrv4
    port map (
            O => \N__41052\,
            I => comm_buf_1_1
        );

    \I__9471\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41041\
        );

    \I__9470\ : InMux
    port map (
            O => \N__41044\,
            I => \N__41034\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__41041\,
            I => \N__41031\
        );

    \I__9468\ : InMux
    port map (
            O => \N__41040\,
            I => \N__41028\
        );

    \I__9467\ : InMux
    port map (
            O => \N__41039\,
            I => \N__41021\
        );

    \I__9466\ : InMux
    port map (
            O => \N__41038\,
            I => \N__41021\
        );

    \I__9465\ : InMux
    port map (
            O => \N__41037\,
            I => \N__41021\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__41034\,
            I => \N__41016\
        );

    \I__9463\ : Span4Mux_v
    port map (
            O => \N__41031\,
            I => \N__41016\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41013\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__41021\,
            I => \N__41010\
        );

    \I__9460\ : Odrv4
    port map (
            O => \N__41016\,
            I => eis_start
        );

    \I__9459\ : Odrv12
    port map (
            O => \N__41013\,
            I => eis_start
        );

    \I__9458\ : Odrv4
    port map (
            O => \N__41010\,
            I => eis_start
        );

    \I__9457\ : CascadeMux
    port map (
            O => \N__41003\,
            I => \N__40999\
        );

    \I__9456\ : CascadeMux
    port map (
            O => \N__41002\,
            I => \N__40996\
        );

    \I__9455\ : InMux
    port map (
            O => \N__40999\,
            I => \N__40993\
        );

    \I__9454\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40990\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__40993\,
            I => \N__40985\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__40990\,
            I => \N__40985\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__40985\,
            I => data_idxvec_8
        );

    \I__9450\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40979\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40976\
        );

    \I__9448\ : Span4Mux_h
    port map (
            O => \N__40976\,
            I => \N__40973\
        );

    \I__9447\ : Odrv4
    port map (
            O => \N__40973\,
            I => n78_adj_1022
        );

    \I__9446\ : InMux
    port map (
            O => \N__40970\,
            I => \N__40966\
        );

    \I__9445\ : InMux
    port map (
            O => \N__40969\,
            I => \N__40962\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__40966\,
            I => \N__40959\
        );

    \I__9443\ : InMux
    port map (
            O => \N__40965\,
            I => \N__40956\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__40962\,
            I => \N__40951\
        );

    \I__9441\ : Span4Mux_v
    port map (
            O => \N__40959\,
            I => \N__40951\
        );

    \I__9440\ : LocalMux
    port map (
            O => \N__40956\,
            I => buf_dds_3
        );

    \I__9439\ : Odrv4
    port map (
            O => \N__40951\,
            I => buf_dds_3
        );

    \I__9438\ : InMux
    port map (
            O => \N__40946\,
            I => \N__40941\
        );

    \I__9437\ : InMux
    port map (
            O => \N__40945\,
            I => \N__40938\
        );

    \I__9436\ : InMux
    port map (
            O => \N__40944\,
            I => \N__40935\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__40941\,
            I => \N__40930\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__40938\,
            I => \N__40930\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__40935\,
            I => n8
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__40930\,
            I => n8
        );

    \I__9431\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40922\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__40922\,
            I => \N__40919\
        );

    \I__9429\ : Span4Mux_h
    port map (
            O => \N__40919\,
            I => \N__40916\
        );

    \I__9428\ : Span4Mux_v
    port map (
            O => \N__40916\,
            I => \N__40913\
        );

    \I__9427\ : Odrv4
    port map (
            O => \N__40913\,
            I => n15188
        );

    \I__9426\ : InMux
    port map (
            O => \N__40910\,
            I => \N__40907\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__40907\,
            I => \N__40903\
        );

    \I__9424\ : InMux
    port map (
            O => \N__40906\,
            I => \N__40900\
        );

    \I__9423\ : Span4Mux_h
    port map (
            O => \N__40903\,
            I => \N__40897\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__40900\,
            I => \N__40894\
        );

    \I__9421\ : Odrv4
    port map (
            O => \N__40897\,
            I => n12702
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__40894\,
            I => n12702
        );

    \I__9419\ : CascadeMux
    port map (
            O => \N__40889\,
            I => \n15188_cascade_\
        );

    \I__9418\ : InMux
    port map (
            O => \N__40886\,
            I => \N__40881\
        );

    \I__9417\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40876\
        );

    \I__9416\ : InMux
    port map (
            O => \N__40884\,
            I => \N__40872\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__40881\,
            I => \N__40869\
        );

    \I__9414\ : InMux
    port map (
            O => \N__40880\,
            I => \N__40864\
        );

    \I__9413\ : InMux
    port map (
            O => \N__40879\,
            I => \N__40864\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__40876\,
            I => \N__40856\
        );

    \I__9411\ : InMux
    port map (
            O => \N__40875\,
            I => \N__40853\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__40872\,
            I => \N__40850\
        );

    \I__9409\ : Span4Mux_h
    port map (
            O => \N__40869\,
            I => \N__40847\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__40864\,
            I => \N__40844\
        );

    \I__9407\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40837\
        );

    \I__9406\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40837\
        );

    \I__9405\ : InMux
    port map (
            O => \N__40861\,
            I => \N__40837\
        );

    \I__9404\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40834\
        );

    \I__9403\ : InMux
    port map (
            O => \N__40859\,
            I => \N__40831\
        );

    \I__9402\ : Span4Mux_v
    port map (
            O => \N__40856\,
            I => \N__40827\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__40853\,
            I => \N__40822\
        );

    \I__9400\ : Span12Mux_h
    port map (
            O => \N__40850\,
            I => \N__40822\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__40847\,
            I => \N__40813\
        );

    \I__9398\ : Span4Mux_h
    port map (
            O => \N__40844\,
            I => \N__40813\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__40837\,
            I => \N__40813\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__40834\,
            I => \N__40813\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__40831\,
            I => \N__40810\
        );

    \I__9394\ : InMux
    port map (
            O => \N__40830\,
            I => \N__40807\
        );

    \I__9393\ : Odrv4
    port map (
            O => \N__40827\,
            I => n8085
        );

    \I__9392\ : Odrv12
    port map (
            O => \N__40822\,
            I => n8085
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__40813\,
            I => n8085
        );

    \I__9390\ : Odrv4
    port map (
            O => \N__40810\,
            I => n8085
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__40807\,
            I => n8085
        );

    \I__9388\ : CascadeMux
    port map (
            O => \N__40796\,
            I => \n6_adj_1171_cascade_\
        );

    \I__9387\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40790\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__40790\,
            I => \N__40787\
        );

    \I__9385\ : Odrv12
    port map (
            O => \N__40787\,
            I => n15190
        );

    \I__9384\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40779\
        );

    \I__9383\ : InMux
    port map (
            O => \N__40783\,
            I => \N__40776\
        );

    \I__9382\ : CascadeMux
    port map (
            O => \N__40782\,
            I => \N__40773\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__40779\,
            I => \N__40770\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__40776\,
            I => \N__40767\
        );

    \I__9379\ : InMux
    port map (
            O => \N__40773\,
            I => \N__40764\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__40770\,
            I => \N__40759\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__40767\,
            I => \N__40759\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__40764\,
            I => buf_adcdata3_12
        );

    \I__9375\ : Odrv4
    port map (
            O => \N__40759\,
            I => buf_adcdata3_12
        );

    \I__9374\ : InMux
    port map (
            O => \N__40754\,
            I => \N__40750\
        );

    \I__9373\ : InMux
    port map (
            O => \N__40753\,
            I => \N__40747\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__40750\,
            I => \N__40744\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__40747\,
            I => n24
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__40744\,
            I => n24
        );

    \I__9369\ : InMux
    port map (
            O => \N__40739\,
            I => \N__40736\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__40736\,
            I => \N__40733\
        );

    \I__9367\ : Span4Mux_v
    port map (
            O => \N__40733\,
            I => \N__40727\
        );

    \I__9366\ : InMux
    port map (
            O => \N__40732\,
            I => \N__40724\
        );

    \I__9365\ : InMux
    port map (
            O => \N__40731\,
            I => \N__40719\
        );

    \I__9364\ : InMux
    port map (
            O => \N__40730\,
            I => \N__40716\
        );

    \I__9363\ : Span4Mux_h
    port map (
            O => \N__40727\,
            I => \N__40710\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__40724\,
            I => \N__40710\
        );

    \I__9361\ : InMux
    port map (
            O => \N__40723\,
            I => \N__40707\
        );

    \I__9360\ : CascadeMux
    port map (
            O => \N__40722\,
            I => \N__40703\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__40719\,
            I => \N__40700\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__40716\,
            I => \N__40697\
        );

    \I__9357\ : InMux
    port map (
            O => \N__40715\,
            I => \N__40694\
        );

    \I__9356\ : Span4Mux_v
    port map (
            O => \N__40710\,
            I => \N__40687\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__40707\,
            I => \N__40684\
        );

    \I__9354\ : InMux
    port map (
            O => \N__40706\,
            I => \N__40681\
        );

    \I__9353\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40678\
        );

    \I__9352\ : Span4Mux_v
    port map (
            O => \N__40700\,
            I => \N__40673\
        );

    \I__9351\ : Span4Mux_h
    port map (
            O => \N__40697\,
            I => \N__40673\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__40694\,
            I => \N__40670\
        );

    \I__9349\ : InMux
    port map (
            O => \N__40693\,
            I => \N__40667\
        );

    \I__9348\ : InMux
    port map (
            O => \N__40692\,
            I => \N__40664\
        );

    \I__9347\ : InMux
    port map (
            O => \N__40691\,
            I => \N__40661\
        );

    \I__9346\ : InMux
    port map (
            O => \N__40690\,
            I => \N__40658\
        );

    \I__9345\ : Span4Mux_h
    port map (
            O => \N__40687\,
            I => \N__40652\
        );

    \I__9344\ : Span4Mux_v
    port map (
            O => \N__40684\,
            I => \N__40652\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__40681\,
            I => \N__40647\
        );

    \I__9342\ : LocalMux
    port map (
            O => \N__40678\,
            I => \N__40647\
        );

    \I__9341\ : Span4Mux_h
    port map (
            O => \N__40673\,
            I => \N__40644\
        );

    \I__9340\ : Span4Mux_h
    port map (
            O => \N__40670\,
            I => \N__40641\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__40667\,
            I => \N__40632\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__40664\,
            I => \N__40632\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__40661\,
            I => \N__40632\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__40658\,
            I => \N__40632\
        );

    \I__9335\ : InMux
    port map (
            O => \N__40657\,
            I => \N__40629\
        );

    \I__9334\ : Span4Mux_h
    port map (
            O => \N__40652\,
            I => \N__40625\
        );

    \I__9333\ : Span12Mux_h
    port map (
            O => \N__40647\,
            I => \N__40622\
        );

    \I__9332\ : Span4Mux_h
    port map (
            O => \N__40644\,
            I => \N__40617\
        );

    \I__9331\ : Span4Mux_v
    port map (
            O => \N__40641\,
            I => \N__40617\
        );

    \I__9330\ : Span12Mux_h
    port map (
            O => \N__40632\,
            I => \N__40614\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__40629\,
            I => \N__40611\
        );

    \I__9328\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40608\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__40625\,
            I => comm_rx_buf_6
        );

    \I__9326\ : Odrv12
    port map (
            O => \N__40622\,
            I => comm_rx_buf_6
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__40617\,
            I => comm_rx_buf_6
        );

    \I__9324\ : Odrv12
    port map (
            O => \N__40614\,
            I => comm_rx_buf_6
        );

    \I__9323\ : Odrv12
    port map (
            O => \N__40611\,
            I => comm_rx_buf_6
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__40608\,
            I => comm_rx_buf_6
        );

    \I__9321\ : InMux
    port map (
            O => \N__40595\,
            I => \N__40592\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__40592\,
            I => \N__40589\
        );

    \I__9319\ : Span4Mux_h
    port map (
            O => \N__40589\,
            I => \N__40586\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__40586\,
            I => buf_data1_19
        );

    \I__9317\ : CascadeMux
    port map (
            O => \N__40583\,
            I => \N__40580\
        );

    \I__9316\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40576\
        );

    \I__9315\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40573\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__40576\,
            I => \N__40570\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__40573\,
            I => data_idxvec_11
        );

    \I__9312\ : Odrv4
    port map (
            O => \N__40570\,
            I => data_idxvec_11
        );

    \I__9311\ : InMux
    port map (
            O => \N__40565\,
            I => \N__40562\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__40562\,
            I => \N__40559\
        );

    \I__9309\ : Span4Mux_h
    port map (
            O => \N__40559\,
            I => \N__40556\
        );

    \I__9308\ : Span4Mux_h
    port map (
            O => \N__40556\,
            I => \N__40553\
        );

    \I__9307\ : Odrv4
    port map (
            O => \N__40553\,
            I => n75
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__40550\,
            I => \n12_cascade_\
        );

    \I__9305\ : InMux
    port map (
            O => \N__40547\,
            I => \N__40540\
        );

    \I__9304\ : InMux
    port map (
            O => \N__40546\,
            I => \N__40535\
        );

    \I__9303\ : InMux
    port map (
            O => \N__40545\,
            I => \N__40535\
        );

    \I__9302\ : InMux
    port map (
            O => \N__40544\,
            I => \N__40529\
        );

    \I__9301\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40525\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__40540\,
            I => \N__40520\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__40535\,
            I => \N__40520\
        );

    \I__9298\ : InMux
    port map (
            O => \N__40534\,
            I => \N__40517\
        );

    \I__9297\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40512\
        );

    \I__9296\ : InMux
    port map (
            O => \N__40532\,
            I => \N__40512\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__40529\,
            I => \N__40509\
        );

    \I__9294\ : InMux
    port map (
            O => \N__40528\,
            I => \N__40506\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__40525\,
            I => \N__40496\
        );

    \I__9292\ : Span4Mux_v
    port map (
            O => \N__40520\,
            I => \N__40496\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__40517\,
            I => \N__40496\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40496\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__40509\,
            I => \N__40493\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__40506\,
            I => \N__40490\
        );

    \I__9287\ : InMux
    port map (
            O => \N__40505\,
            I => \N__40487\
        );

    \I__9286\ : Span4Mux_v
    port map (
            O => \N__40496\,
            I => \N__40484\
        );

    \I__9285\ : Sp12to4
    port map (
            O => \N__40493\,
            I => \N__40477\
        );

    \I__9284\ : Span12Mux_v
    port map (
            O => \N__40490\,
            I => \N__40477\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__40487\,
            I => \N__40477\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__40484\,
            I => n6301
        );

    \I__9281\ : Odrv12
    port map (
            O => \N__40477\,
            I => n6301
        );

    \I__9280\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40465\
        );

    \I__9279\ : InMux
    port map (
            O => \N__40471\,
            I => \N__40465\
        );

    \I__9278\ : InMux
    port map (
            O => \N__40470\,
            I => \N__40451\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__40465\,
            I => \N__40448\
        );

    \I__9276\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40445\
        );

    \I__9275\ : InMux
    port map (
            O => \N__40463\,
            I => \N__40438\
        );

    \I__9274\ : InMux
    port map (
            O => \N__40462\,
            I => \N__40438\
        );

    \I__9273\ : InMux
    port map (
            O => \N__40461\,
            I => \N__40438\
        );

    \I__9272\ : CascadeMux
    port map (
            O => \N__40460\,
            I => \N__40435\
        );

    \I__9271\ : InMux
    port map (
            O => \N__40459\,
            I => \N__40428\
        );

    \I__9270\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40428\
        );

    \I__9269\ : InMux
    port map (
            O => \N__40457\,
            I => \N__40425\
        );

    \I__9268\ : InMux
    port map (
            O => \N__40456\,
            I => \N__40422\
        );

    \I__9267\ : InMux
    port map (
            O => \N__40455\,
            I => \N__40419\
        );

    \I__9266\ : InMux
    port map (
            O => \N__40454\,
            I => \N__40416\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__40451\,
            I => \N__40413\
        );

    \I__9264\ : Span4Mux_v
    port map (
            O => \N__40448\,
            I => \N__40408\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__40445\,
            I => \N__40408\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40405\
        );

    \I__9261\ : InMux
    port map (
            O => \N__40435\,
            I => \N__40400\
        );

    \I__9260\ : InMux
    port map (
            O => \N__40434\,
            I => \N__40400\
        );

    \I__9259\ : InMux
    port map (
            O => \N__40433\,
            I => \N__40397\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__40428\,
            I => \N__40394\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__40425\,
            I => \N__40391\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__40422\,
            I => \N__40388\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__40419\,
            I => \N__40381\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__40416\,
            I => \N__40381\
        );

    \I__9253\ : Span4Mux_v
    port map (
            O => \N__40413\,
            I => \N__40381\
        );

    \I__9252\ : Span4Mux_v
    port map (
            O => \N__40408\,
            I => \N__40378\
        );

    \I__9251\ : Span4Mux_v
    port map (
            O => \N__40405\,
            I => \N__40375\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__40400\,
            I => \N__40368\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__40397\,
            I => \N__40368\
        );

    \I__9248\ : Span4Mux_v
    port map (
            O => \N__40394\,
            I => \N__40368\
        );

    \I__9247\ : Span12Mux_v
    port map (
            O => \N__40391\,
            I => \N__40365\
        );

    \I__9246\ : Span4Mux_v
    port map (
            O => \N__40388\,
            I => \N__40358\
        );

    \I__9245\ : Span4Mux_v
    port map (
            O => \N__40381\,
            I => \N__40358\
        );

    \I__9244\ : Span4Mux_h
    port map (
            O => \N__40378\,
            I => \N__40358\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__40375\,
            I => n8253
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__40368\,
            I => n8253
        );

    \I__9241\ : Odrv12
    port map (
            O => \N__40365\,
            I => n8253
        );

    \I__9240\ : Odrv4
    port map (
            O => \N__40358\,
            I => n8253
        );

    \I__9239\ : InMux
    port map (
            O => \N__40349\,
            I => \N__40346\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__40346\,
            I => \N__40342\
        );

    \I__9237\ : InMux
    port map (
            O => \N__40345\,
            I => \N__40339\
        );

    \I__9236\ : Span4Mux_v
    port map (
            O => \N__40342\,
            I => \N__40336\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__40339\,
            I => \N__40333\
        );

    \I__9234\ : Sp12to4
    port map (
            O => \N__40336\,
            I => \N__40330\
        );

    \I__9233\ : Odrv4
    port map (
            O => \N__40333\,
            I => n14_adj_1197
        );

    \I__9232\ : Odrv12
    port map (
            O => \N__40330\,
            I => n14_adj_1197
        );

    \I__9231\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40320\
        );

    \I__9230\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40317\
        );

    \I__9229\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40314\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__40320\,
            I => \N__40309\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__40317\,
            I => \N__40309\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__40314\,
            I => req_data_cnt_2
        );

    \I__9225\ : Odrv12
    port map (
            O => \N__40309\,
            I => req_data_cnt_2
        );

    \I__9224\ : InMux
    port map (
            O => \N__40304\,
            I => \N__40299\
        );

    \I__9223\ : InMux
    port map (
            O => \N__40303\,
            I => \N__40294\
        );

    \I__9222\ : InMux
    port map (
            O => \N__40302\,
            I => \N__40294\
        );

    \I__9221\ : LocalMux
    port map (
            O => \N__40299\,
            I => comm_cmd_5
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__40294\,
            I => comm_cmd_5
        );

    \I__9219\ : InMux
    port map (
            O => \N__40289\,
            I => \N__40285\
        );

    \I__9218\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40281\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__40285\,
            I => \N__40278\
        );

    \I__9216\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40275\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__40281\,
            I => comm_cmd_4
        );

    \I__9214\ : Odrv4
    port map (
            O => \N__40278\,
            I => comm_cmd_4
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__40275\,
            I => comm_cmd_4
        );

    \I__9212\ : InMux
    port map (
            O => \N__40268\,
            I => \N__40263\
        );

    \I__9211\ : InMux
    port map (
            O => \N__40267\,
            I => \N__40258\
        );

    \I__9210\ : InMux
    port map (
            O => \N__40266\,
            I => \N__40258\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__40263\,
            I => comm_cmd_6
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__40258\,
            I => comm_cmd_6
        );

    \I__9207\ : InMux
    port map (
            O => \N__40253\,
            I => \N__40248\
        );

    \I__9206\ : InMux
    port map (
            O => \N__40252\,
            I => \N__40245\
        );

    \I__9205\ : InMux
    port map (
            O => \N__40251\,
            I => \N__40242\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__40248\,
            I => \N__40234\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__40245\,
            I => \N__40229\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__40242\,
            I => \N__40229\
        );

    \I__9201\ : InMux
    port map (
            O => \N__40241\,
            I => \N__40226\
        );

    \I__9200\ : InMux
    port map (
            O => \N__40240\,
            I => \N__40221\
        );

    \I__9199\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40218\
        );

    \I__9198\ : InMux
    port map (
            O => \N__40238\,
            I => \N__40213\
        );

    \I__9197\ : InMux
    port map (
            O => \N__40237\,
            I => \N__40213\
        );

    \I__9196\ : Span4Mux_v
    port map (
            O => \N__40234\,
            I => \N__40203\
        );

    \I__9195\ : Span4Mux_h
    port map (
            O => \N__40229\,
            I => \N__40203\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__40226\,
            I => \N__40203\
        );

    \I__9193\ : CascadeMux
    port map (
            O => \N__40225\,
            I => \N__40200\
        );

    \I__9192\ : CascadeMux
    port map (
            O => \N__40224\,
            I => \N__40197\
        );

    \I__9191\ : LocalMux
    port map (
            O => \N__40221\,
            I => \N__40190\
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__40218\,
            I => \N__40190\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__40213\,
            I => \N__40187\
        );

    \I__9188\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40184\
        );

    \I__9187\ : InMux
    port map (
            O => \N__40211\,
            I => \N__40181\
        );

    \I__9186\ : InMux
    port map (
            O => \N__40210\,
            I => \N__40178\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__40203\,
            I => \N__40175\
        );

    \I__9184\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40172\
        );

    \I__9183\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40165\
        );

    \I__9182\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40165\
        );

    \I__9181\ : InMux
    port map (
            O => \N__40195\,
            I => \N__40165\
        );

    \I__9180\ : Span4Mux_v
    port map (
            O => \N__40190\,
            I => \N__40161\
        );

    \I__9179\ : Span4Mux_v
    port map (
            O => \N__40187\,
            I => \N__40156\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__40184\,
            I => \N__40156\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__40181\,
            I => \N__40151\
        );

    \I__9176\ : LocalMux
    port map (
            O => \N__40178\,
            I => \N__40151\
        );

    \I__9175\ : Span4Mux_h
    port map (
            O => \N__40175\,
            I => \N__40148\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__40172\,
            I => \N__40143\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__40165\,
            I => \N__40143\
        );

    \I__9172\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40140\
        );

    \I__9171\ : Span4Mux_h
    port map (
            O => \N__40161\,
            I => \N__40135\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__40156\,
            I => \N__40135\
        );

    \I__9169\ : Odrv12
    port map (
            O => \N__40151\,
            I => n8043
        );

    \I__9168\ : Odrv4
    port map (
            O => \N__40148\,
            I => n8043
        );

    \I__9167\ : Odrv4
    port map (
            O => \N__40143\,
            I => n8043
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__40140\,
            I => n8043
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__40135\,
            I => n8043
        );

    \I__9164\ : InMux
    port map (
            O => \N__40124\,
            I => \N__40113\
        );

    \I__9163\ : InMux
    port map (
            O => \N__40123\,
            I => \N__40110\
        );

    \I__9162\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40107\
        );

    \I__9161\ : InMux
    port map (
            O => \N__40121\,
            I => \N__40104\
        );

    \I__9160\ : InMux
    port map (
            O => \N__40120\,
            I => \N__40101\
        );

    \I__9159\ : InMux
    port map (
            O => \N__40119\,
            I => \N__40098\
        );

    \I__9158\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40095\
        );

    \I__9157\ : InMux
    port map (
            O => \N__40117\,
            I => \N__40092\
        );

    \I__9156\ : InMux
    port map (
            O => \N__40116\,
            I => \N__40089\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__40113\,
            I => \N__40082\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__40110\,
            I => \N__40082\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__40107\,
            I => \N__40082\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__40104\,
            I => \N__40077\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__40077\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__40098\,
            I => \N__40068\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__40095\,
            I => \N__40068\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__40092\,
            I => \N__40068\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__40089\,
            I => \N__40065\
        );

    \I__9146\ : Span4Mux_v
    port map (
            O => \N__40082\,
            I => \N__40060\
        );

    \I__9145\ : Span4Mux_v
    port map (
            O => \N__40077\,
            I => \N__40060\
        );

    \I__9144\ : InMux
    port map (
            O => \N__40076\,
            I => \N__40057\
        );

    \I__9143\ : InMux
    port map (
            O => \N__40075\,
            I => \N__40054\
        );

    \I__9142\ : Span4Mux_v
    port map (
            O => \N__40068\,
            I => \N__40050\
        );

    \I__9141\ : Span4Mux_h
    port map (
            O => \N__40065\,
            I => \N__40047\
        );

    \I__9140\ : Span4Mux_h
    port map (
            O => \N__40060\,
            I => \N__40040\
        );

    \I__9139\ : LocalMux
    port map (
            O => \N__40057\,
            I => \N__40040\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__40054\,
            I => \N__40040\
        );

    \I__9137\ : InMux
    port map (
            O => \N__40053\,
            I => \N__40037\
        );

    \I__9136\ : Span4Mux_h
    port map (
            O => \N__40050\,
            I => \N__40033\
        );

    \I__9135\ : Span4Mux_v
    port map (
            O => \N__40047\,
            I => \N__40028\
        );

    \I__9134\ : Span4Mux_h
    port map (
            O => \N__40040\,
            I => \N__40028\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__40037\,
            I => \N__40025\
        );

    \I__9132\ : InMux
    port map (
            O => \N__40036\,
            I => \N__40022\
        );

    \I__9131\ : Span4Mux_h
    port map (
            O => \N__40033\,
            I => \N__40018\
        );

    \I__9130\ : Span4Mux_h
    port map (
            O => \N__40028\,
            I => \N__40015\
        );

    \I__9129\ : Span12Mux_h
    port map (
            O => \N__40025\,
            I => \N__40010\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__40022\,
            I => \N__40010\
        );

    \I__9127\ : InMux
    port map (
            O => \N__40021\,
            I => \N__40007\
        );

    \I__9126\ : Odrv4
    port map (
            O => \N__40018\,
            I => comm_rx_buf_2
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__40015\,
            I => comm_rx_buf_2
        );

    \I__9124\ : Odrv12
    port map (
            O => \N__40010\,
            I => comm_rx_buf_2
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__40007\,
            I => comm_rx_buf_2
        );

    \I__9122\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39992\
        );

    \I__9121\ : InMux
    port map (
            O => \N__39997\,
            I => \N__39989\
        );

    \I__9120\ : InMux
    port map (
            O => \N__39996\,
            I => \N__39986\
        );

    \I__9119\ : InMux
    port map (
            O => \N__39995\,
            I => \N__39983\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__39992\,
            I => \N__39980\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__39989\,
            I => \N__39977\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__39986\,
            I => \N__39974\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__39983\,
            I => \N__39971\
        );

    \I__9114\ : Span4Mux_h
    port map (
            O => \N__39980\,
            I => \N__39965\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__39977\,
            I => \N__39965\
        );

    \I__9112\ : Span4Mux_v
    port map (
            O => \N__39974\,
            I => \N__39960\
        );

    \I__9111\ : Span4Mux_h
    port map (
            O => \N__39971\,
            I => \N__39960\
        );

    \I__9110\ : InMux
    port map (
            O => \N__39970\,
            I => \N__39957\
        );

    \I__9109\ : Sp12to4
    port map (
            O => \N__39965\,
            I => \N__39952\
        );

    \I__9108\ : Sp12to4
    port map (
            O => \N__39960\,
            I => \N__39952\
        );

    \I__9107\ : LocalMux
    port map (
            O => \N__39957\,
            I => comm_buf_1_2
        );

    \I__9106\ : Odrv12
    port map (
            O => \N__39952\,
            I => comm_buf_1_2
        );

    \I__9105\ : InMux
    port map (
            O => \N__39947\,
            I => \N__39944\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__39944\,
            I => \N__39941\
        );

    \I__9103\ : Span4Mux_v
    port map (
            O => \N__39941\,
            I => \N__39936\
        );

    \I__9102\ : InMux
    port map (
            O => \N__39940\,
            I => \N__39933\
        );

    \I__9101\ : InMux
    port map (
            O => \N__39939\,
            I => \N__39929\
        );

    \I__9100\ : Span4Mux_h
    port map (
            O => \N__39936\,
            I => \N__39923\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__39933\,
            I => \N__39923\
        );

    \I__9098\ : InMux
    port map (
            O => \N__39932\,
            I => \N__39919\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__39929\,
            I => \N__39916\
        );

    \I__9096\ : InMux
    port map (
            O => \N__39928\,
            I => \N__39911\
        );

    \I__9095\ : Span4Mux_v
    port map (
            O => \N__39923\,
            I => \N__39908\
        );

    \I__9094\ : InMux
    port map (
            O => \N__39922\,
            I => \N__39905\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__39919\,
            I => \N__39900\
        );

    \I__9092\ : Span4Mux_h
    port map (
            O => \N__39916\,
            I => \N__39897\
        );

    \I__9091\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39894\
        );

    \I__9090\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39891\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__39911\,
            I => \N__39888\
        );

    \I__9088\ : Span4Mux_v
    port map (
            O => \N__39908\,
            I => \N__39882\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__39905\,
            I => \N__39882\
        );

    \I__9086\ : InMux
    port map (
            O => \N__39904\,
            I => \N__39879\
        );

    \I__9085\ : InMux
    port map (
            O => \N__39903\,
            I => \N__39875\
        );

    \I__9084\ : Span4Mux_h
    port map (
            O => \N__39900\,
            I => \N__39872\
        );

    \I__9083\ : Span4Mux_v
    port map (
            O => \N__39897\,
            I => \N__39863\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39863\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__39891\,
            I => \N__39863\
        );

    \I__9080\ : Span4Mux_v
    port map (
            O => \N__39888\,
            I => \N__39863\
        );

    \I__9079\ : InMux
    port map (
            O => \N__39887\,
            I => \N__39860\
        );

    \I__9078\ : Span4Mux_h
    port map (
            O => \N__39882\,
            I => \N__39854\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__39879\,
            I => \N__39854\
        );

    \I__9076\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39851\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__39875\,
            I => \N__39848\
        );

    \I__9074\ : Sp12to4
    port map (
            O => \N__39872\,
            I => \N__39841\
        );

    \I__9073\ : Sp12to4
    port map (
            O => \N__39863\,
            I => \N__39841\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__39860\,
            I => \N__39841\
        );

    \I__9071\ : InMux
    port map (
            O => \N__39859\,
            I => \N__39838\
        );

    \I__9070\ : Span4Mux_h
    port map (
            O => \N__39854\,
            I => \N__39833\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__39851\,
            I => \N__39833\
        );

    \I__9068\ : Span12Mux_h
    port map (
            O => \N__39848\,
            I => \N__39825\
        );

    \I__9067\ : Span12Mux_v
    port map (
            O => \N__39841\,
            I => \N__39825\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__39838\,
            I => \N__39825\
        );

    \I__9065\ : Span4Mux_v
    port map (
            O => \N__39833\,
            I => \N__39822\
        );

    \I__9064\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39819\
        );

    \I__9063\ : Odrv12
    port map (
            O => \N__39825\,
            I => comm_rx_buf_4
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__39822\,
            I => comm_rx_buf_4
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__39819\,
            I => comm_rx_buf_4
        );

    \I__9060\ : CascadeMux
    port map (
            O => \N__39812\,
            I => \n10363_cascade_\
        );

    \I__9059\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39805\
        );

    \I__9058\ : InMux
    port map (
            O => \N__39808\,
            I => \N__39799\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__39805\,
            I => \N__39792\
        );

    \I__9056\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39789\
        );

    \I__9055\ : InMux
    port map (
            O => \N__39803\,
            I => \N__39786\
        );

    \I__9054\ : CascadeMux
    port map (
            O => \N__39802\,
            I => \N__39782\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__39799\,
            I => \N__39779\
        );

    \I__9052\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39776\
        );

    \I__9051\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39773\
        );

    \I__9050\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39770\
        );

    \I__9049\ : CascadeMux
    port map (
            O => \N__39795\,
            I => \N__39767\
        );

    \I__9048\ : Span4Mux_v
    port map (
            O => \N__39792\,
            I => \N__39760\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__39789\,
            I => \N__39760\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__39786\,
            I => \N__39757\
        );

    \I__9045\ : InMux
    port map (
            O => \N__39785\,
            I => \N__39754\
        );

    \I__9044\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39751\
        );

    \I__9043\ : Span4Mux_v
    port map (
            O => \N__39779\,
            I => \N__39746\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__39776\,
            I => \N__39746\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__39773\,
            I => \N__39741\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__39770\,
            I => \N__39741\
        );

    \I__9039\ : InMux
    port map (
            O => \N__39767\,
            I => \N__39738\
        );

    \I__9038\ : InMux
    port map (
            O => \N__39766\,
            I => \N__39735\
        );

    \I__9037\ : InMux
    port map (
            O => \N__39765\,
            I => \N__39732\
        );

    \I__9036\ : Span4Mux_h
    port map (
            O => \N__39760\,
            I => \N__39728\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__39757\,
            I => \N__39723\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__39754\,
            I => \N__39723\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__39751\,
            I => \N__39720\
        );

    \I__9032\ : Span4Mux_v
    port map (
            O => \N__39746\,
            I => \N__39711\
        );

    \I__9031\ : Span4Mux_h
    port map (
            O => \N__39741\,
            I => \N__39711\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__39738\,
            I => \N__39711\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__39735\,
            I => \N__39711\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__39732\,
            I => \N__39708\
        );

    \I__9027\ : CascadeMux
    port map (
            O => \N__39731\,
            I => \N__39705\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__39728\,
            I => \N__39700\
        );

    \I__9025\ : Span4Mux_h
    port map (
            O => \N__39723\,
            I => \N__39700\
        );

    \I__9024\ : Span4Mux_v
    port map (
            O => \N__39720\,
            I => \N__39695\
        );

    \I__9023\ : Span4Mux_h
    port map (
            O => \N__39711\,
            I => \N__39695\
        );

    \I__9022\ : Span4Mux_v
    port map (
            O => \N__39708\,
            I => \N__39692\
        );

    \I__9021\ : InMux
    port map (
            O => \N__39705\,
            I => \N__39689\
        );

    \I__9020\ : Span4Mux_h
    port map (
            O => \N__39700\,
            I => \N__39685\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__39695\,
            I => \N__39682\
        );

    \I__9018\ : Sp12to4
    port map (
            O => \N__39692\,
            I => \N__39677\
        );

    \I__9017\ : LocalMux
    port map (
            O => \N__39689\,
            I => \N__39677\
        );

    \I__9016\ : InMux
    port map (
            O => \N__39688\,
            I => \N__39674\
        );

    \I__9015\ : Odrv4
    port map (
            O => \N__39685\,
            I => comm_rx_buf_5
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__39682\,
            I => comm_rx_buf_5
        );

    \I__9013\ : Odrv12
    port map (
            O => \N__39677\,
            I => comm_rx_buf_5
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__39674\,
            I => comm_rx_buf_5
        );

    \I__9011\ : InMux
    port map (
            O => \N__39665\,
            I => \N__39659\
        );

    \I__9010\ : CascadeMux
    port map (
            O => \N__39664\,
            I => \N__39656\
        );

    \I__9009\ : CascadeMux
    port map (
            O => \N__39663\,
            I => \N__39651\
        );

    \I__9008\ : InMux
    port map (
            O => \N__39662\,
            I => \N__39647\
        );

    \I__9007\ : LocalMux
    port map (
            O => \N__39659\,
            I => \N__39644\
        );

    \I__9006\ : InMux
    port map (
            O => \N__39656\,
            I => \N__39641\
        );

    \I__9005\ : InMux
    port map (
            O => \N__39655\,
            I => \N__39635\
        );

    \I__9004\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39635\
        );

    \I__9003\ : InMux
    port map (
            O => \N__39651\,
            I => \N__39632\
        );

    \I__9002\ : InMux
    port map (
            O => \N__39650\,
            I => \N__39629\
        );

    \I__9001\ : LocalMux
    port map (
            O => \N__39647\,
            I => \N__39622\
        );

    \I__9000\ : Span4Mux_v
    port map (
            O => \N__39644\,
            I => \N__39622\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__39641\,
            I => \N__39622\
        );

    \I__8998\ : InMux
    port map (
            O => \N__39640\,
            I => \N__39619\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__39635\,
            I => \N__39614\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__39632\,
            I => \N__39614\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__39629\,
            I => \N__39609\
        );

    \I__8994\ : Span4Mux_h
    port map (
            O => \N__39622\,
            I => \N__39609\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__39619\,
            I => \N__39606\
        );

    \I__8992\ : Span4Mux_h
    port map (
            O => \N__39614\,
            I => \N__39603\
        );

    \I__8991\ : Span4Mux_h
    port map (
            O => \N__39609\,
            I => \N__39600\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__39606\,
            I => n8062
        );

    \I__8989\ : Odrv4
    port map (
            O => \N__39603\,
            I => n8062
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__39600\,
            I => n8062
        );

    \I__8987\ : CascadeMux
    port map (
            O => \N__39593\,
            I => \n8085_cascade_\
        );

    \I__8986\ : InMux
    port map (
            O => \N__39590\,
            I => \N__39587\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__8984\ : Odrv4
    port map (
            O => \N__39584\,
            I => n14_adj_1152
        );

    \I__8983\ : CascadeMux
    port map (
            O => \N__39581\,
            I => \N__39577\
        );

    \I__8982\ : CascadeMux
    port map (
            O => \N__39580\,
            I => \N__39574\
        );

    \I__8981\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39571\
        );

    \I__8980\ : InMux
    port map (
            O => \N__39574\,
            I => \N__39565\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__39571\,
            I => \N__39562\
        );

    \I__8978\ : InMux
    port map (
            O => \N__39570\,
            I => \N__39557\
        );

    \I__8977\ : InMux
    port map (
            O => \N__39569\,
            I => \N__39557\
        );

    \I__8976\ : InMux
    port map (
            O => \N__39568\,
            I => \N__39553\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__39565\,
            I => \N__39549\
        );

    \I__8974\ : Span4Mux_v
    port map (
            O => \N__39562\,
            I => \N__39544\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__39557\,
            I => \N__39544\
        );

    \I__8972\ : CascadeMux
    port map (
            O => \N__39556\,
            I => \N__39538\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__39553\,
            I => \N__39535\
        );

    \I__8970\ : InMux
    port map (
            O => \N__39552\,
            I => \N__39532\
        );

    \I__8969\ : Span4Mux_h
    port map (
            O => \N__39549\,
            I => \N__39527\
        );

    \I__8968\ : Span4Mux_h
    port map (
            O => \N__39544\,
            I => \N__39527\
        );

    \I__8967\ : InMux
    port map (
            O => \N__39543\,
            I => \N__39524\
        );

    \I__8966\ : InMux
    port map (
            O => \N__39542\,
            I => \N__39521\
        );

    \I__8965\ : InMux
    port map (
            O => \N__39541\,
            I => \N__39518\
        );

    \I__8964\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39515\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__39535\,
            I => \N__39512\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__39532\,
            I => \N__39509\
        );

    \I__8961\ : Span4Mux_h
    port map (
            O => \N__39527\,
            I => \N__39506\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__39524\,
            I => \N__39497\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__39521\,
            I => \N__39497\
        );

    \I__8958\ : LocalMux
    port map (
            O => \N__39518\,
            I => \N__39497\
        );

    \I__8957\ : LocalMux
    port map (
            O => \N__39515\,
            I => \N__39497\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__39512\,
            I => \N__39494\
        );

    \I__8955\ : Span4Mux_h
    port map (
            O => \N__39509\,
            I => \N__39491\
        );

    \I__8954\ : Span4Mux_h
    port map (
            O => \N__39506\,
            I => \N__39488\
        );

    \I__8953\ : Span12Mux_h
    port map (
            O => \N__39497\,
            I => \N__39485\
        );

    \I__8952\ : Odrv4
    port map (
            O => \N__39494\,
            I => n93
        );

    \I__8951\ : Odrv4
    port map (
            O => \N__39491\,
            I => n93
        );

    \I__8950\ : Odrv4
    port map (
            O => \N__39488\,
            I => n93
        );

    \I__8949\ : Odrv12
    port map (
            O => \N__39485\,
            I => n93
        );

    \I__8948\ : CascadeMux
    port map (
            O => \N__39476\,
            I => \N__39472\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__39475\,
            I => \N__39469\
        );

    \I__8946\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39466\
        );

    \I__8945\ : InMux
    port map (
            O => \N__39469\,
            I => \N__39463\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__39466\,
            I => \N__39458\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__39463\,
            I => \N__39458\
        );

    \I__8942\ : Span4Mux_h
    port map (
            O => \N__39458\,
            I => \N__39455\
        );

    \I__8941\ : Odrv4
    port map (
            O => \N__39455\,
            I => n27
        );

    \I__8940\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__39449\,
            I => n4
        );

    \I__8938\ : CascadeMux
    port map (
            O => \N__39446\,
            I => \n15309_cascade_\
        );

    \I__8937\ : CascadeMux
    port map (
            O => \N__39443\,
            I => \N__39440\
        );

    \I__8936\ : InMux
    port map (
            O => \N__39440\,
            I => \N__39437\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__39437\,
            I => \N__39433\
        );

    \I__8934\ : InMux
    port map (
            O => \N__39436\,
            I => \N__39430\
        );

    \I__8933\ : Odrv4
    port map (
            O => \N__39433\,
            I => \comm_state_3_N_402_3\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__39430\,
            I => \comm_state_3_N_402_3\
        );

    \I__8931\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39422\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__39422\,
            I => \N__39419\
        );

    \I__8929\ : Odrv4
    port map (
            O => \N__39419\,
            I => n15637
        );

    \I__8928\ : InMux
    port map (
            O => \N__39416\,
            I => \N__39413\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__39413\,
            I => n13_adj_1040
        );

    \I__8926\ : InMux
    port map (
            O => \N__39410\,
            I => \N__39407\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__39407\,
            I => \N__39404\
        );

    \I__8924\ : Odrv4
    port map (
            O => \N__39404\,
            I => n22_adj_1078
        );

    \I__8923\ : CascadeMux
    port map (
            O => \N__39401\,
            I => \N__39398\
        );

    \I__8922\ : InMux
    port map (
            O => \N__39398\,
            I => \N__39391\
        );

    \I__8921\ : InMux
    port map (
            O => \N__39397\,
            I => \N__39387\
        );

    \I__8920\ : InMux
    port map (
            O => \N__39396\,
            I => \N__39384\
        );

    \I__8919\ : InMux
    port map (
            O => \N__39395\,
            I => \N__39380\
        );

    \I__8918\ : InMux
    port map (
            O => \N__39394\,
            I => \N__39377\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__39391\,
            I => \N__39374\
        );

    \I__8916\ : InMux
    port map (
            O => \N__39390\,
            I => \N__39371\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__39387\,
            I => \N__39368\
        );

    \I__8914\ : LocalMux
    port map (
            O => \N__39384\,
            I => \N__39365\
        );

    \I__8913\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39362\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__39380\,
            I => \N__39355\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__39377\,
            I => \N__39355\
        );

    \I__8910\ : Span4Mux_v
    port map (
            O => \N__39374\,
            I => \N__39350\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__39371\,
            I => \N__39350\
        );

    \I__8908\ : Span4Mux_v
    port map (
            O => \N__39368\,
            I => \N__39347\
        );

    \I__8907\ : Span4Mux_v
    port map (
            O => \N__39365\,
            I => \N__39342\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__39362\,
            I => \N__39342\
        );

    \I__8905\ : InMux
    port map (
            O => \N__39361\,
            I => \N__39339\
        );

    \I__8904\ : InMux
    port map (
            O => \N__39360\,
            I => \N__39335\
        );

    \I__8903\ : Span4Mux_v
    port map (
            O => \N__39355\,
            I => \N__39328\
        );

    \I__8902\ : Span4Mux_v
    port map (
            O => \N__39350\,
            I => \N__39328\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__39347\,
            I => \N__39323\
        );

    \I__8900\ : Span4Mux_v
    port map (
            O => \N__39342\,
            I => \N__39323\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__39339\,
            I => \N__39320\
        );

    \I__8898\ : InMux
    port map (
            O => \N__39338\,
            I => \N__39317\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__39335\,
            I => \N__39314\
        );

    \I__8896\ : InMux
    port map (
            O => \N__39334\,
            I => \N__39311\
        );

    \I__8895\ : InMux
    port map (
            O => \N__39333\,
            I => \N__39308\
        );

    \I__8894\ : Span4Mux_h
    port map (
            O => \N__39328\,
            I => \N__39304\
        );

    \I__8893\ : Span4Mux_h
    port map (
            O => \N__39323\,
            I => \N__39301\
        );

    \I__8892\ : Span4Mux_v
    port map (
            O => \N__39320\,
            I => \N__39298\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__39317\,
            I => \N__39289\
        );

    \I__8890\ : Sp12to4
    port map (
            O => \N__39314\,
            I => \N__39289\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__39311\,
            I => \N__39289\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__39308\,
            I => \N__39289\
        );

    \I__8887\ : InMux
    port map (
            O => \N__39307\,
            I => \N__39286\
        );

    \I__8886\ : Span4Mux_h
    port map (
            O => \N__39304\,
            I => \N__39283\
        );

    \I__8885\ : Span4Mux_h
    port map (
            O => \N__39301\,
            I => \N__39278\
        );

    \I__8884\ : Span4Mux_v
    port map (
            O => \N__39298\,
            I => \N__39278\
        );

    \I__8883\ : Span12Mux_h
    port map (
            O => \N__39289\,
            I => \N__39275\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__39286\,
            I => \N__39272\
        );

    \I__8881\ : Odrv4
    port map (
            O => \N__39283\,
            I => comm_rx_buf_7
        );

    \I__8880\ : Odrv4
    port map (
            O => \N__39278\,
            I => comm_rx_buf_7
        );

    \I__8879\ : Odrv12
    port map (
            O => \N__39275\,
            I => comm_rx_buf_7
        );

    \I__8878\ : Odrv12
    port map (
            O => \N__39272\,
            I => comm_rx_buf_7
        );

    \I__8877\ : InMux
    port map (
            O => \N__39263\,
            I => \N__39260\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__39260\,
            I => \N__39257\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__39257\,
            I => \N__39251\
        );

    \I__8874\ : InMux
    port map (
            O => \N__39256\,
            I => \N__39248\
        );

    \I__8873\ : CascadeMux
    port map (
            O => \N__39255\,
            I => \N__39245\
        );

    \I__8872\ : InMux
    port map (
            O => \N__39254\,
            I => \N__39242\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__39251\,
            I => \N__39239\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__39248\,
            I => \N__39236\
        );

    \I__8869\ : InMux
    port map (
            O => \N__39245\,
            I => \N__39233\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__39242\,
            I => \N__39230\
        );

    \I__8867\ : Span4Mux_h
    port map (
            O => \N__39239\,
            I => \N__39227\
        );

    \I__8866\ : Span12Mux_v
    port map (
            O => \N__39236\,
            I => \N__39224\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__39233\,
            I => comm_cmd_7
        );

    \I__8864\ : Odrv4
    port map (
            O => \N__39230\,
            I => comm_cmd_7
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__39227\,
            I => comm_cmd_7
        );

    \I__8862\ : Odrv12
    port map (
            O => \N__39224\,
            I => comm_cmd_7
        );

    \I__8861\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39210\
        );

    \I__8860\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39206\
        );

    \I__8859\ : InMux
    port map (
            O => \N__39213\,
            I => \N__39202\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__39210\,
            I => \N__39198\
        );

    \I__8857\ : InMux
    port map (
            O => \N__39209\,
            I => \N__39195\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__39206\,
            I => \N__39192\
        );

    \I__8855\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39189\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__39202\,
            I => \N__39184\
        );

    \I__8853\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39181\
        );

    \I__8852\ : Span4Mux_v
    port map (
            O => \N__39198\,
            I => \N__39170\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39170\
        );

    \I__8850\ : Span4Mux_v
    port map (
            O => \N__39192\,
            I => \N__39170\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__39189\,
            I => \N__39167\
        );

    \I__8848\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39164\
        );

    \I__8847\ : InMux
    port map (
            O => \N__39187\,
            I => \N__39161\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__39184\,
            I => \N__39158\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__39181\,
            I => \N__39155\
        );

    \I__8844\ : InMux
    port map (
            O => \N__39180\,
            I => \N__39152\
        );

    \I__8843\ : InMux
    port map (
            O => \N__39179\,
            I => \N__39149\
        );

    \I__8842\ : InMux
    port map (
            O => \N__39178\,
            I => \N__39146\
        );

    \I__8841\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39143\
        );

    \I__8840\ : Span4Mux_h
    port map (
            O => \N__39170\,
            I => \N__39135\
        );

    \I__8839\ : Span4Mux_v
    port map (
            O => \N__39167\,
            I => \N__39135\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__39164\,
            I => \N__39135\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__39161\,
            I => \N__39132\
        );

    \I__8836\ : Span4Mux_h
    port map (
            O => \N__39158\,
            I => \N__39119\
        );

    \I__8835\ : Span4Mux_v
    port map (
            O => \N__39155\,
            I => \N__39119\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__39152\,
            I => \N__39119\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__39149\,
            I => \N__39119\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__39146\,
            I => \N__39119\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__39143\,
            I => \N__39119\
        );

    \I__8830\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39115\
        );

    \I__8829\ : Span4Mux_h
    port map (
            O => \N__39135\,
            I => \N__39112\
        );

    \I__8828\ : Span4Mux_v
    port map (
            O => \N__39132\,
            I => \N__39109\
        );

    \I__8827\ : Span4Mux_v
    port map (
            O => \N__39119\,
            I => \N__39106\
        );

    \I__8826\ : InMux
    port map (
            O => \N__39118\,
            I => \N__39103\
        );

    \I__8825\ : LocalMux
    port map (
            O => \N__39115\,
            I => \N__39100\
        );

    \I__8824\ : Span4Mux_h
    port map (
            O => \N__39112\,
            I => \N__39097\
        );

    \I__8823\ : Span4Mux_v
    port map (
            O => \N__39109\,
            I => \N__39092\
        );

    \I__8822\ : Span4Mux_h
    port map (
            O => \N__39106\,
            I => \N__39092\
        );

    \I__8821\ : LocalMux
    port map (
            O => \N__39103\,
            I => comm_rx_buf_0
        );

    \I__8820\ : Odrv12
    port map (
            O => \N__39100\,
            I => comm_rx_buf_0
        );

    \I__8819\ : Odrv4
    port map (
            O => \N__39097\,
            I => comm_rx_buf_0
        );

    \I__8818\ : Odrv4
    port map (
            O => \N__39092\,
            I => comm_rx_buf_0
        );

    \I__8817\ : InMux
    port map (
            O => \N__39083\,
            I => \N__39077\
        );

    \I__8816\ : InMux
    port map (
            O => \N__39082\,
            I => \N__39077\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__39077\,
            I => n8530
        );

    \I__8814\ : InMux
    port map (
            O => \N__39074\,
            I => \N__39068\
        );

    \I__8813\ : InMux
    port map (
            O => \N__39073\,
            I => \N__39068\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__39068\,
            I => n15198
        );

    \I__8811\ : InMux
    port map (
            O => \N__39065\,
            I => \N__39062\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__39062\,
            I => n15266
        );

    \I__8809\ : CascadeMux
    port map (
            O => \N__39059\,
            I => \n15410_cascade_\
        );

    \I__8808\ : CEMux
    port map (
            O => \N__39056\,
            I => \N__39053\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__39053\,
            I => n15130
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__39050\,
            I => \N__39047\
        );

    \I__8805\ : InMux
    port map (
            O => \N__39047\,
            I => \N__39044\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__39044\,
            I => n15408
        );

    \I__8803\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39037\
        );

    \I__8802\ : InMux
    port map (
            O => \N__39040\,
            I => \N__39034\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__39037\,
            I => n10394
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__39034\,
            I => n10394
        );

    \I__8799\ : InMux
    port map (
            O => \N__39029\,
            I => \N__39026\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__39026\,
            I => n16190
        );

    \I__8797\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39020\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__39020\,
            I => n15635
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__39017\,
            I => \N__39014\
        );

    \I__8794\ : InMux
    port map (
            O => \N__39014\,
            I => \N__39010\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__39013\,
            I => \N__39007\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__39010\,
            I => \N__39004\
        );

    \I__8791\ : InMux
    port map (
            O => \N__39007\,
            I => \N__39001\
        );

    \I__8790\ : Odrv4
    port map (
            O => \N__39004\,
            I => n12_adj_1027
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__39001\,
            I => n12_adj_1027
        );

    \I__8788\ : InMux
    port map (
            O => \N__38996\,
            I => \N__38992\
        );

    \I__8787\ : InMux
    port map (
            O => \N__38995\,
            I => \N__38989\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__38992\,
            I => \N__38984\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__38989\,
            I => \N__38984\
        );

    \I__8784\ : Span4Mux_v
    port map (
            O => \N__38984\,
            I => \N__38981\
        );

    \I__8783\ : Odrv4
    port map (
            O => \N__38981\,
            I => n12622
        );

    \I__8782\ : InMux
    port map (
            O => \N__38978\,
            I => \N__38973\
        );

    \I__8781\ : InMux
    port map (
            O => \N__38977\,
            I => \N__38968\
        );

    \I__8780\ : InMux
    port map (
            O => \N__38976\,
            I => \N__38965\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__38973\,
            I => \N__38962\
        );

    \I__8778\ : InMux
    port map (
            O => \N__38972\,
            I => \N__38959\
        );

    \I__8777\ : CascadeMux
    port map (
            O => \N__38971\,
            I => \N__38956\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__38968\,
            I => \N__38953\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__38965\,
            I => \N__38948\
        );

    \I__8774\ : Span4Mux_h
    port map (
            O => \N__38962\,
            I => \N__38948\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__38959\,
            I => \N__38945\
        );

    \I__8772\ : InMux
    port map (
            O => \N__38956\,
            I => \N__38942\
        );

    \I__8771\ : Span4Mux_h
    port map (
            O => \N__38953\,
            I => \N__38939\
        );

    \I__8770\ : Sp12to4
    port map (
            O => \N__38948\,
            I => \N__38936\
        );

    \I__8769\ : Odrv4
    port map (
            O => \N__38945\,
            I => comm_buf_1_7
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__38942\,
            I => comm_buf_1_7
        );

    \I__8767\ : Odrv4
    port map (
            O => \N__38939\,
            I => comm_buf_1_7
        );

    \I__8766\ : Odrv12
    port map (
            O => \N__38936\,
            I => comm_buf_1_7
        );

    \I__8765\ : InMux
    port map (
            O => \N__38927\,
            I => \N__38920\
        );

    \I__8764\ : InMux
    port map (
            O => \N__38926\,
            I => \N__38917\
        );

    \I__8763\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38914\
        );

    \I__8762\ : InMux
    port map (
            O => \N__38924\,
            I => \N__38911\
        );

    \I__8761\ : InMux
    port map (
            O => \N__38923\,
            I => \N__38908\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__38920\,
            I => \N__38905\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__38917\,
            I => \N__38899\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38899\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__38911\,
            I => \N__38896\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__38908\,
            I => \N__38893\
        );

    \I__8755\ : Span4Mux_h
    port map (
            O => \N__38905\,
            I => \N__38890\
        );

    \I__8754\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38887\
        );

    \I__8753\ : Span4Mux_v
    port map (
            O => \N__38899\,
            I => \N__38884\
        );

    \I__8752\ : Span4Mux_v
    port map (
            O => \N__38896\,
            I => \N__38881\
        );

    \I__8751\ : Span4Mux_h
    port map (
            O => \N__38893\,
            I => \N__38878\
        );

    \I__8750\ : Span4Mux_h
    port map (
            O => \N__38890\,
            I => \N__38875\
        );

    \I__8749\ : LocalMux
    port map (
            O => \N__38887\,
            I => \N__38868\
        );

    \I__8748\ : Span4Mux_h
    port map (
            O => \N__38884\,
            I => \N__38868\
        );

    \I__8747\ : Span4Mux_h
    port map (
            O => \N__38881\,
            I => \N__38868\
        );

    \I__8746\ : Span4Mux_h
    port map (
            O => \N__38878\,
            I => \N__38865\
        );

    \I__8745\ : Span4Mux_v
    port map (
            O => \N__38875\,
            I => \N__38862\
        );

    \I__8744\ : Sp12to4
    port map (
            O => \N__38868\,
            I => \N__38859\
        );

    \I__8743\ : Span4Mux_h
    port map (
            O => \N__38865\,
            I => \N__38854\
        );

    \I__8742\ : Span4Mux_h
    port map (
            O => \N__38862\,
            I => \N__38854\
        );

    \I__8741\ : Odrv12
    port map (
            O => \N__38859\,
            I => comm_buf_0_7
        );

    \I__8740\ : Odrv4
    port map (
            O => \N__38854\,
            I => comm_buf_0_7
        );

    \I__8739\ : InMux
    port map (
            O => \N__38849\,
            I => \N__38816\
        );

    \I__8738\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38816\
        );

    \I__8737\ : InMux
    port map (
            O => \N__38847\,
            I => \N__38811\
        );

    \I__8736\ : InMux
    port map (
            O => \N__38846\,
            I => \N__38811\
        );

    \I__8735\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38802\
        );

    \I__8734\ : InMux
    port map (
            O => \N__38844\,
            I => \N__38802\
        );

    \I__8733\ : InMux
    port map (
            O => \N__38843\,
            I => \N__38802\
        );

    \I__8732\ : InMux
    port map (
            O => \N__38842\,
            I => \N__38795\
        );

    \I__8731\ : InMux
    port map (
            O => \N__38841\,
            I => \N__38795\
        );

    \I__8730\ : InMux
    port map (
            O => \N__38840\,
            I => \N__38795\
        );

    \I__8729\ : InMux
    port map (
            O => \N__38839\,
            I => \N__38790\
        );

    \I__8728\ : InMux
    port map (
            O => \N__38838\,
            I => \N__38790\
        );

    \I__8727\ : InMux
    port map (
            O => \N__38837\,
            I => \N__38776\
        );

    \I__8726\ : InMux
    port map (
            O => \N__38836\,
            I => \N__38767\
        );

    \I__8725\ : InMux
    port map (
            O => \N__38835\,
            I => \N__38767\
        );

    \I__8724\ : InMux
    port map (
            O => \N__38834\,
            I => \N__38767\
        );

    \I__8723\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38767\
        );

    \I__8722\ : InMux
    port map (
            O => \N__38832\,
            I => \N__38760\
        );

    \I__8721\ : InMux
    port map (
            O => \N__38831\,
            I => \N__38753\
        );

    \I__8720\ : InMux
    port map (
            O => \N__38830\,
            I => \N__38753\
        );

    \I__8719\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38753\
        );

    \I__8718\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38746\
        );

    \I__8717\ : InMux
    port map (
            O => \N__38827\,
            I => \N__38746\
        );

    \I__8716\ : InMux
    port map (
            O => \N__38826\,
            I => \N__38746\
        );

    \I__8715\ : InMux
    port map (
            O => \N__38825\,
            I => \N__38735\
        );

    \I__8714\ : InMux
    port map (
            O => \N__38824\,
            I => \N__38735\
        );

    \I__8713\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38735\
        );

    \I__8712\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38735\
        );

    \I__8711\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38735\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__38816\,
            I => \N__38730\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__38811\,
            I => \N__38730\
        );

    \I__8708\ : InMux
    port map (
            O => \N__38810\,
            I => \N__38725\
        );

    \I__8707\ : InMux
    port map (
            O => \N__38809\,
            I => \N__38725\
        );

    \I__8706\ : LocalMux
    port map (
            O => \N__38802\,
            I => \N__38718\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__38795\,
            I => \N__38718\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__38790\,
            I => \N__38718\
        );

    \I__8703\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38711\
        );

    \I__8702\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38711\
        );

    \I__8701\ : InMux
    port map (
            O => \N__38787\,
            I => \N__38711\
        );

    \I__8700\ : InMux
    port map (
            O => \N__38786\,
            I => \N__38704\
        );

    \I__8699\ : InMux
    port map (
            O => \N__38785\,
            I => \N__38704\
        );

    \I__8698\ : InMux
    port map (
            O => \N__38784\,
            I => \N__38704\
        );

    \I__8697\ : InMux
    port map (
            O => \N__38783\,
            I => \N__38699\
        );

    \I__8696\ : InMux
    port map (
            O => \N__38782\,
            I => \N__38699\
        );

    \I__8695\ : InMux
    port map (
            O => \N__38781\,
            I => \N__38694\
        );

    \I__8694\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38694\
        );

    \I__8693\ : InMux
    port map (
            O => \N__38779\,
            I => \N__38690\
        );

    \I__8692\ : LocalMux
    port map (
            O => \N__38776\,
            I => \N__38686\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__38767\,
            I => \N__38683\
        );

    \I__8690\ : InMux
    port map (
            O => \N__38766\,
            I => \N__38680\
        );

    \I__8689\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38675\
        );

    \I__8688\ : InMux
    port map (
            O => \N__38764\,
            I => \N__38675\
        );

    \I__8687\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38672\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__38760\,
            I => \N__38669\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__38753\,
            I => \N__38666\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__38746\,
            I => \N__38655\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__38735\,
            I => \N__38655\
        );

    \I__8682\ : Span4Mux_v
    port map (
            O => \N__38730\,
            I => \N__38655\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__38725\,
            I => \N__38655\
        );

    \I__8680\ : Span4Mux_v
    port map (
            O => \N__38718\,
            I => \N__38655\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__38711\,
            I => \N__38646\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__38704\,
            I => \N__38646\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__38699\,
            I => \N__38646\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__38694\,
            I => \N__38646\
        );

    \I__8675\ : CascadeMux
    port map (
            O => \N__38693\,
            I => \N__38643\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__38690\,
            I => \N__38639\
        );

    \I__8673\ : InMux
    port map (
            O => \N__38689\,
            I => \N__38636\
        );

    \I__8672\ : Span4Mux_v
    port map (
            O => \N__38686\,
            I => \N__38631\
        );

    \I__8671\ : Span4Mux_v
    port map (
            O => \N__38683\,
            I => \N__38631\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__38680\,
            I => \N__38619\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__38675\,
            I => \N__38619\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__38672\,
            I => \N__38619\
        );

    \I__8667\ : Span4Mux_v
    port map (
            O => \N__38669\,
            I => \N__38619\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__38666\,
            I => \N__38619\
        );

    \I__8665\ : Span4Mux_h
    port map (
            O => \N__38655\,
            I => \N__38614\
        );

    \I__8664\ : Span4Mux_v
    port map (
            O => \N__38646\,
            I => \N__38614\
        );

    \I__8663\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38609\
        );

    \I__8662\ : InMux
    port map (
            O => \N__38642\,
            I => \N__38609\
        );

    \I__8661\ : Span4Mux_v
    port map (
            O => \N__38639\,
            I => \N__38602\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__38636\,
            I => \N__38602\
        );

    \I__8659\ : Span4Mux_h
    port map (
            O => \N__38631\,
            I => \N__38602\
        );

    \I__8658\ : InMux
    port map (
            O => \N__38630\,
            I => \N__38599\
        );

    \I__8657\ : Span4Mux_h
    port map (
            O => \N__38619\,
            I => \N__38596\
        );

    \I__8656\ : Span4Mux_h
    port map (
            O => \N__38614\,
            I => \N__38593\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__38609\,
            I => comm_index_0
        );

    \I__8654\ : Odrv4
    port map (
            O => \N__38602\,
            I => comm_index_0
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__38599\,
            I => comm_index_0
        );

    \I__8652\ : Odrv4
    port map (
            O => \N__38596\,
            I => comm_index_0
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__38593\,
            I => comm_index_0
        );

    \I__8650\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38579\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__38579\,
            I => \N__38576\
        );

    \I__8648\ : Span12Mux_h
    port map (
            O => \N__38576\,
            I => \N__38573\
        );

    \I__8647\ : Odrv12
    port map (
            O => \N__38573\,
            I => n15381
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__38570\,
            I => \n12846_cascade_\
        );

    \I__8645\ : InMux
    port map (
            O => \N__38567\,
            I => \N__38564\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__38564\,
            I => n4_adj_1179
        );

    \I__8643\ : CascadeMux
    port map (
            O => \N__38561\,
            I => \N__38555\
        );

    \I__8642\ : CascadeMux
    port map (
            O => \N__38560\,
            I => \N__38552\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__38559\,
            I => \N__38549\
        );

    \I__8640\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38545\
        );

    \I__8639\ : InMux
    port map (
            O => \N__38555\,
            I => \N__38538\
        );

    \I__8638\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38538\
        );

    \I__8637\ : InMux
    port map (
            O => \N__38549\,
            I => \N__38538\
        );

    \I__8636\ : CascadeMux
    port map (
            O => \N__38548\,
            I => \N__38535\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__38545\,
            I => \N__38530\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__38538\,
            I => \N__38527\
        );

    \I__8633\ : InMux
    port map (
            O => \N__38535\,
            I => \N__38522\
        );

    \I__8632\ : InMux
    port map (
            O => \N__38534\,
            I => \N__38522\
        );

    \I__8631\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38519\
        );

    \I__8630\ : Span4Mux_h
    port map (
            O => \N__38530\,
            I => \N__38516\
        );

    \I__8629\ : Span4Mux_v
    port map (
            O => \N__38527\,
            I => \N__38511\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__38522\,
            I => \N__38511\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__38519\,
            I => \N__38508\
        );

    \I__8626\ : Odrv4
    port map (
            O => \N__38516\,
            I => n15204
        );

    \I__8625\ : Odrv4
    port map (
            O => \N__38511\,
            I => n15204
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__38508\,
            I => n15204
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__38501\,
            I => \n4_adj_1184_cascade_\
        );

    \I__8622\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38495\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__38495\,
            I => \N__38492\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__38492\,
            I => n15290
        );

    \I__8619\ : CascadeMux
    port map (
            O => \N__38489\,
            I => \n15241_cascade_\
        );

    \I__8618\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38480\
        );

    \I__8617\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38480\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__38480\,
            I => n15108
        );

    \I__8615\ : CEMux
    port map (
            O => \N__38477\,
            I => \N__38474\
        );

    \I__8614\ : LocalMux
    port map (
            O => \N__38474\,
            I => \N__38471\
        );

    \I__8613\ : Span4Mux_v
    port map (
            O => \N__38471\,
            I => \N__38468\
        );

    \I__8612\ : Odrv4
    port map (
            O => \N__38468\,
            I => n15128
        );

    \I__8611\ : InMux
    port map (
            O => \N__38465\,
            I => \N__38462\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__38462\,
            I => \N__38459\
        );

    \I__8609\ : Span4Mux_v
    port map (
            O => \N__38459\,
            I => \N__38456\
        );

    \I__8608\ : Odrv4
    port map (
            O => \N__38456\,
            I => \comm_spi.n10438\
        );

    \I__8607\ : SRMux
    port map (
            O => \N__38453\,
            I => \N__38450\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__38450\,
            I => \N__38447\
        );

    \I__8605\ : Span4Mux_h
    port map (
            O => \N__38447\,
            I => \N__38444\
        );

    \I__8604\ : Span4Mux_h
    port map (
            O => \N__38444\,
            I => \N__38441\
        );

    \I__8603\ : Odrv4
    port map (
            O => \N__38441\,
            I => \comm_spi.iclk_N_802\
        );

    \I__8602\ : InMux
    port map (
            O => \N__38438\,
            I => \N__38435\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__38435\,
            I => \comm_spi.n16890\
        );

    \I__8600\ : InMux
    port map (
            O => \N__38432\,
            I => \N__38429\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__38429\,
            I => \comm_spi.n10455\
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__38426\,
            I => \comm_spi.n16890_cascade_\
        );

    \I__8597\ : InMux
    port map (
            O => \N__38423\,
            I => \N__38420\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__38420\,
            I => \N__38409\
        );

    \I__8595\ : InMux
    port map (
            O => \N__38419\,
            I => \N__38406\
        );

    \I__8594\ : InMux
    port map (
            O => \N__38418\,
            I => \N__38391\
        );

    \I__8593\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38391\
        );

    \I__8592\ : InMux
    port map (
            O => \N__38416\,
            I => \N__38391\
        );

    \I__8591\ : InMux
    port map (
            O => \N__38415\,
            I => \N__38391\
        );

    \I__8590\ : InMux
    port map (
            O => \N__38414\,
            I => \N__38391\
        );

    \I__8589\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38391\
        );

    \I__8588\ : InMux
    port map (
            O => \N__38412\,
            I => \N__38391\
        );

    \I__8587\ : Odrv12
    port map (
            O => \N__38409\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__38406\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__38391\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__8584\ : InMux
    port map (
            O => \N__38384\,
            I => \N__38381\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__38381\,
            I => \N__38378\
        );

    \I__8582\ : Span4Mux_v
    port map (
            O => \N__38378\,
            I => \N__38368\
        );

    \I__8581\ : InMux
    port map (
            O => \N__38377\,
            I => \N__38353\
        );

    \I__8580\ : InMux
    port map (
            O => \N__38376\,
            I => \N__38353\
        );

    \I__8579\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38353\
        );

    \I__8578\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38353\
        );

    \I__8577\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38353\
        );

    \I__8576\ : InMux
    port map (
            O => \N__38372\,
            I => \N__38353\
        );

    \I__8575\ : InMux
    port map (
            O => \N__38371\,
            I => \N__38353\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__38368\,
            I => \comm_spi.n12175\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__38353\,
            I => \comm_spi.n12175\
        );

    \I__8572\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38344\
        );

    \I__8571\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38341\
        );

    \I__8570\ : LocalMux
    port map (
            O => \N__38344\,
            I => \N__38338\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__38341\,
            I => data_idxvec_5
        );

    \I__8568\ : Odrv4
    port map (
            O => \N__38338\,
            I => data_idxvec_5
        );

    \I__8567\ : InMux
    port map (
            O => \N__38333\,
            I => \N__38328\
        );

    \I__8566\ : InMux
    port map (
            O => \N__38332\,
            I => \N__38325\
        );

    \I__8565\ : InMux
    port map (
            O => \N__38331\,
            I => \N__38322\
        );

    \I__8564\ : LocalMux
    port map (
            O => \N__38328\,
            I => data_cntvec_5
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__38325\,
            I => data_cntvec_5
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__38322\,
            I => data_cntvec_5
        );

    \I__8561\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38312\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__38312\,
            I => \N__38309\
        );

    \I__8559\ : Span4Mux_h
    port map (
            O => \N__38309\,
            I => \N__38306\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__38306\,
            I => buf_data1_13
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__38303\,
            I => \n4192_cascade_\
        );

    \I__8556\ : InMux
    port map (
            O => \N__38300\,
            I => \N__38297\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__38297\,
            I => n4229
        );

    \I__8554\ : CascadeMux
    port map (
            O => \N__38294\,
            I => \N__38291\
        );

    \I__8553\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38288\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__38288\,
            I => \N__38285\
        );

    \I__8551\ : Sp12to4
    port map (
            O => \N__38285\,
            I => \N__38280\
        );

    \I__8550\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38277\
        );

    \I__8549\ : CascadeMux
    port map (
            O => \N__38283\,
            I => \N__38274\
        );

    \I__8548\ : Span12Mux_s9_v
    port map (
            O => \N__38280\,
            I => \N__38269\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__38277\,
            I => \N__38269\
        );

    \I__8546\ : InMux
    port map (
            O => \N__38274\,
            I => \N__38266\
        );

    \I__8545\ : Odrv12
    port map (
            O => \N__38269\,
            I => cmd_rdadctmp_18_adj_1058
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__38266\,
            I => cmd_rdadctmp_18_adj_1058
        );

    \I__8543\ : InMux
    port map (
            O => \N__38261\,
            I => \N__38258\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__38258\,
            I => \N__38254\
        );

    \I__8541\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38251\
        );

    \I__8540\ : Span4Mux_v
    port map (
            O => \N__38254\,
            I => \N__38248\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__38251\,
            I => buf_adcdata2_10
        );

    \I__8538\ : Odrv4
    port map (
            O => \N__38248\,
            I => buf_adcdata2_10
        );

    \I__8537\ : InMux
    port map (
            O => \N__38243\,
            I => \N__38239\
        );

    \I__8536\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38236\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38233\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__38236\,
            I => data_idxvec_1
        );

    \I__8533\ : Odrv12
    port map (
            O => \N__38233\,
            I => data_idxvec_1
        );

    \I__8532\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38224\
        );

    \I__8531\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38220\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__38224\,
            I => \N__38217\
        );

    \I__8529\ : InMux
    port map (
            O => \N__38223\,
            I => \N__38214\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__38220\,
            I => data_cntvec_1
        );

    \I__8527\ : Odrv4
    port map (
            O => \N__38217\,
            I => data_cntvec_1
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__38214\,
            I => data_cntvec_1
        );

    \I__8525\ : CascadeMux
    port map (
            O => \N__38207\,
            I => \N__38204\
        );

    \I__8524\ : InMux
    port map (
            O => \N__38204\,
            I => \N__38201\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__38201\,
            I => \N__38197\
        );

    \I__8522\ : InMux
    port map (
            O => \N__38200\,
            I => \N__38194\
        );

    \I__8521\ : Sp12to4
    port map (
            O => \N__38197\,
            I => \N__38188\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__38194\,
            I => \N__38188\
        );

    \I__8519\ : CascadeMux
    port map (
            O => \N__38193\,
            I => \N__38185\
        );

    \I__8518\ : Span12Mux_h
    port map (
            O => \N__38188\,
            I => \N__38182\
        );

    \I__8517\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38179\
        );

    \I__8516\ : Odrv12
    port map (
            O => \N__38182\,
            I => cmd_rdadctmp_16_adj_1096
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__38179\,
            I => cmd_rdadctmp_16_adj_1096
        );

    \I__8514\ : InMux
    port map (
            O => \N__38174\,
            I => \N__38171\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__38171\,
            I => \N__38167\
        );

    \I__8512\ : InMux
    port map (
            O => \N__38170\,
            I => \N__38163\
        );

    \I__8511\ : Span4Mux_v
    port map (
            O => \N__38167\,
            I => \N__38160\
        );

    \I__8510\ : InMux
    port map (
            O => \N__38166\,
            I => \N__38157\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__38163\,
            I => req_data_cnt_3
        );

    \I__8508\ : Odrv4
    port map (
            O => \N__38160\,
            I => req_data_cnt_3
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__38157\,
            I => req_data_cnt_3
        );

    \I__8506\ : InMux
    port map (
            O => \N__38150\,
            I => \N__38147\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__38147\,
            I => \N__38142\
        );

    \I__8504\ : InMux
    port map (
            O => \N__38146\,
            I => \N__38137\
        );

    \I__8503\ : InMux
    port map (
            O => \N__38145\,
            I => \N__38137\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__38142\,
            I => \acadc_skipCount_3\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__38137\,
            I => \acadc_skipCount_3\
        );

    \I__8500\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38128\
        );

    \I__8499\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38124\
        );

    \I__8498\ : LocalMux
    port map (
            O => \N__38128\,
            I => \N__38119\
        );

    \I__8497\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38116\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__38124\,
            I => \N__38113\
        );

    \I__8495\ : InMux
    port map (
            O => \N__38123\,
            I => \N__38108\
        );

    \I__8494\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38108\
        );

    \I__8493\ : Span4Mux_v
    port map (
            O => \N__38119\,
            I => \N__38103\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__38116\,
            I => \N__38103\
        );

    \I__8491\ : Span4Mux_h
    port map (
            O => \N__38113\,
            I => \N__38098\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__38108\,
            I => \N__38098\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__38103\,
            I => \N__38087\
        );

    \I__8488\ : Span4Mux_v
    port map (
            O => \N__38098\,
            I => \N__38084\
        );

    \I__8487\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38081\
        );

    \I__8486\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38074\
        );

    \I__8485\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38074\
        );

    \I__8484\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38074\
        );

    \I__8483\ : InMux
    port map (
            O => \N__38093\,
            I => \N__38071\
        );

    \I__8482\ : InMux
    port map (
            O => \N__38092\,
            I => \N__38064\
        );

    \I__8481\ : InMux
    port map (
            O => \N__38091\,
            I => \N__38064\
        );

    \I__8480\ : InMux
    port map (
            O => \N__38090\,
            I => \N__38064\
        );

    \I__8479\ : Span4Mux_h
    port map (
            O => \N__38087\,
            I => \N__38061\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__38084\,
            I => eis_state_1
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__38081\,
            I => eis_state_1
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__38074\,
            I => eis_state_1
        );

    \I__8475\ : LocalMux
    port map (
            O => \N__38071\,
            I => eis_state_1
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__38064\,
            I => eis_state_1
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__38061\,
            I => eis_state_1
        );

    \I__8472\ : CEMux
    port map (
            O => \N__38048\,
            I => \N__38044\
        );

    \I__8471\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38038\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__38044\,
            I => \N__38035\
        );

    \I__8469\ : CEMux
    port map (
            O => \N__38043\,
            I => \N__38032\
        );

    \I__8468\ : CEMux
    port map (
            O => \N__38042\,
            I => \N__38029\
        );

    \I__8467\ : CEMux
    port map (
            O => \N__38041\,
            I => \N__38026\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__38038\,
            I => \N__38023\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__38035\,
            I => \N__38016\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__38032\,
            I => \N__38016\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__38029\,
            I => \N__38016\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38011\
        );

    \I__8461\ : Span4Mux_v
    port map (
            O => \N__38023\,
            I => \N__38011\
        );

    \I__8460\ : Odrv4
    port map (
            O => \N__38016\,
            I => n9790
        );

    \I__8459\ : Odrv4
    port map (
            O => \N__38011\,
            I => n9790
        );

    \I__8458\ : SRMux
    port map (
            O => \N__38006\,
            I => \N__38002\
        );

    \I__8457\ : SRMux
    port map (
            O => \N__38005\,
            I => \N__37999\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__38002\,
            I => \N__37996\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__37999\,
            I => \N__37991\
        );

    \I__8454\ : Span4Mux_v
    port map (
            O => \N__37996\,
            I => \N__37988\
        );

    \I__8453\ : SRMux
    port map (
            O => \N__37995\,
            I => \N__37985\
        );

    \I__8452\ : SRMux
    port map (
            O => \N__37994\,
            I => \N__37982\
        );

    \I__8451\ : Span12Mux_v
    port map (
            O => \N__37991\,
            I => \N__37979\
        );

    \I__8450\ : Span4Mux_h
    port map (
            O => \N__37988\,
            I => \N__37976\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__37985\,
            I => n10483
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__37982\,
            I => n10483
        );

    \I__8447\ : Odrv12
    port map (
            O => \N__37979\,
            I => n10483
        );

    \I__8446\ : Odrv4
    port map (
            O => \N__37976\,
            I => n10483
        );

    \I__8445\ : InMux
    port map (
            O => \N__37967\,
            I => \N__37964\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__37964\,
            I => \N__37961\
        );

    \I__8443\ : Span4Mux_v
    port map (
            O => \N__37961\,
            I => \N__37957\
        );

    \I__8442\ : InMux
    port map (
            O => \N__37960\,
            I => \N__37954\
        );

    \I__8441\ : Odrv4
    port map (
            O => \N__37957\,
            I => \comm_spi.n16887\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__37954\,
            I => \comm_spi.n16887\
        );

    \I__8439\ : InMux
    port map (
            O => \N__37949\,
            I => \N__37946\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__37946\,
            I => \N__37942\
        );

    \I__8437\ : InMux
    port map (
            O => \N__37945\,
            I => \N__37939\
        );

    \I__8436\ : Span4Mux_v
    port map (
            O => \N__37942\,
            I => \N__37934\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__37939\,
            I => \N__37934\
        );

    \I__8434\ : Span4Mux_v
    port map (
            O => \N__37934\,
            I => \N__37931\
        );

    \I__8433\ : Span4Mux_h
    port map (
            O => \N__37931\,
            I => \N__37928\
        );

    \I__8432\ : Span4Mux_h
    port map (
            O => \N__37928\,
            I => \N__37925\
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__37925\,
            I => n14_adj_1169
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__37922\,
            I => \N__37918\
        );

    \I__8429\ : InMux
    port map (
            O => \N__37921\,
            I => \N__37912\
        );

    \I__8428\ : InMux
    port map (
            O => \N__37918\,
            I => \N__37912\
        );

    \I__8427\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37909\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__37912\,
            I => \N__37906\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__37909\,
            I => req_data_cnt_6
        );

    \I__8424\ : Odrv4
    port map (
            O => \N__37906\,
            I => req_data_cnt_6
        );

    \I__8423\ : InMux
    port map (
            O => \N__37901\,
            I => \N__37898\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__37898\,
            I => \N__37895\
        );

    \I__8421\ : Span4Mux_v
    port map (
            O => \N__37895\,
            I => \N__37892\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__37892\,
            I => n4204
        );

    \I__8419\ : CascadeMux
    port map (
            O => \N__37889\,
            I => \n4249_cascade_\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__37886\,
            I => \n4259_cascade_\
        );

    \I__8417\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37879\
        );

    \I__8416\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37875\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__37879\,
            I => \N__37871\
        );

    \I__8414\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37867\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__37875\,
            I => \N__37864\
        );

    \I__8412\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37861\
        );

    \I__8411\ : Span4Mux_h
    port map (
            O => \N__37871\,
            I => \N__37858\
        );

    \I__8410\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37855\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__37867\,
            I => \N__37852\
        );

    \I__8408\ : Span4Mux_v
    port map (
            O => \N__37864\,
            I => \N__37847\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__37861\,
            I => \N__37847\
        );

    \I__8406\ : Span4Mux_v
    port map (
            O => \N__37858\,
            I => \N__37844\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__37855\,
            I => \N__37841\
        );

    \I__8404\ : Span12Mux_h
    port map (
            O => \N__37852\,
            I => \N__37838\
        );

    \I__8403\ : Odrv4
    port map (
            O => \N__37847\,
            I => comm_buf_1_5
        );

    \I__8402\ : Odrv4
    port map (
            O => \N__37844\,
            I => comm_buf_1_5
        );

    \I__8401\ : Odrv4
    port map (
            O => \N__37841\,
            I => comm_buf_1_5
        );

    \I__8400\ : Odrv12
    port map (
            O => \N__37838\,
            I => comm_buf_1_5
        );

    \I__8399\ : CascadeMux
    port map (
            O => \N__37829\,
            I => \N__37825\
        );

    \I__8398\ : InMux
    port map (
            O => \N__37828\,
            I => \N__37822\
        );

    \I__8397\ : InMux
    port map (
            O => \N__37825\,
            I => \N__37819\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__37822\,
            I => \N__37816\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__37819\,
            I => data_idxvec_4
        );

    \I__8394\ : Odrv4
    port map (
            O => \N__37816\,
            I => data_idxvec_4
        );

    \I__8393\ : InMux
    port map (
            O => \N__37811\,
            I => \N__37807\
        );

    \I__8392\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37803\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__37807\,
            I => \N__37800\
        );

    \I__8390\ : InMux
    port map (
            O => \N__37806\,
            I => \N__37797\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__37803\,
            I => data_cntvec_4
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__37800\,
            I => data_cntvec_4
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__37797\,
            I => data_cntvec_4
        );

    \I__8386\ : InMux
    port map (
            O => \N__37790\,
            I => \N__37787\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__37787\,
            I => \N__37784\
        );

    \I__8384\ : Span4Mux_v
    port map (
            O => \N__37784\,
            I => \N__37781\
        );

    \I__8383\ : Span4Mux_h
    port map (
            O => \N__37781\,
            I => \N__37778\
        );

    \I__8382\ : Odrv4
    port map (
            O => \N__37778\,
            I => buf_data1_12
        );

    \I__8381\ : CascadeMux
    port map (
            O => \N__37775\,
            I => \n4193_cascade_\
        );

    \I__8380\ : CascadeMux
    port map (
            O => \N__37772\,
            I => \N__37768\
        );

    \I__8379\ : CascadeMux
    port map (
            O => \N__37771\,
            I => \N__37764\
        );

    \I__8378\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37761\
        );

    \I__8377\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37758\
        );

    \I__8376\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37755\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__37761\,
            I => req_data_cnt_5
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__37758\,
            I => req_data_cnt_5
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__37755\,
            I => req_data_cnt_5
        );

    \I__8372\ : InMux
    port map (
            O => \N__37748\,
            I => \N__37745\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37742\
        );

    \I__8370\ : Span4Mux_h
    port map (
            O => \N__37742\,
            I => \N__37737\
        );

    \I__8369\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37732\
        );

    \I__8368\ : InMux
    port map (
            O => \N__37740\,
            I => \N__37732\
        );

    \I__8367\ : Odrv4
    port map (
            O => \N__37737\,
            I => \acadc_skipCount_5\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__37732\,
            I => \acadc_skipCount_5\
        );

    \I__8365\ : InMux
    port map (
            O => \N__37727\,
            I => \N__37724\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__37724\,
            I => n4216
        );

    \I__8363\ : InMux
    port map (
            O => \N__37721\,
            I => n14050
        );

    \I__8362\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37715\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__37715\,
            I => \N__37712\
        );

    \I__8360\ : Span4Mux_v
    port map (
            O => \N__37712\,
            I => \N__37708\
        );

    \I__8359\ : InMux
    port map (
            O => \N__37711\,
            I => \N__37705\
        );

    \I__8358\ : Sp12to4
    port map (
            O => \N__37708\,
            I => \N__37702\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37699\
        );

    \I__8356\ : Span12Mux_s11_h
    port map (
            O => \N__37702\,
            I => \N__37696\
        );

    \I__8355\ : Span4Mux_h
    port map (
            O => \N__37699\,
            I => \N__37693\
        );

    \I__8354\ : Odrv12
    port map (
            O => \N__37696\,
            I => n14_adj_1207
        );

    \I__8353\ : Odrv4
    port map (
            O => \N__37693\,
            I => n14_adj_1207
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__37688\,
            I => \N__37684\
        );

    \I__8351\ : InMux
    port map (
            O => \N__37687\,
            I => \N__37681\
        );

    \I__8350\ : InMux
    port map (
            O => \N__37684\,
            I => \N__37678\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__37681\,
            I => \N__37675\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__37678\,
            I => data_idxvec_12
        );

    \I__8347\ : Odrv4
    port map (
            O => \N__37675\,
            I => data_idxvec_12
        );

    \I__8346\ : InMux
    port map (
            O => \N__37670\,
            I => n14051
        );

    \I__8345\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37664\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37660\
        );

    \I__8343\ : InMux
    port map (
            O => \N__37663\,
            I => \N__37657\
        );

    \I__8342\ : Span4Mux_h
    port map (
            O => \N__37660\,
            I => \N__37654\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__37657\,
            I => n14_adj_1202
        );

    \I__8340\ : Odrv4
    port map (
            O => \N__37654\,
            I => n14_adj_1202
        );

    \I__8339\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37645\
        );

    \I__8338\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37642\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__37645\,
            I => \N__37639\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__37642\,
            I => data_idxvec_13
        );

    \I__8335\ : Odrv4
    port map (
            O => \N__37639\,
            I => data_idxvec_13
        );

    \I__8334\ : InMux
    port map (
            O => \N__37634\,
            I => n14052
        );

    \I__8333\ : InMux
    port map (
            O => \N__37631\,
            I => \N__37627\
        );

    \I__8332\ : InMux
    port map (
            O => \N__37630\,
            I => \N__37624\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__37627\,
            I => \N__37621\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__37624\,
            I => \N__37618\
        );

    \I__8329\ : Span4Mux_h
    port map (
            O => \N__37621\,
            I => \N__37615\
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__37618\,
            I => n14_adj_1206
        );

    \I__8327\ : Odrv4
    port map (
            O => \N__37615\,
            I => n14_adj_1206
        );

    \I__8326\ : CascadeMux
    port map (
            O => \N__37610\,
            I => \N__37607\
        );

    \I__8325\ : InMux
    port map (
            O => \N__37607\,
            I => \N__37603\
        );

    \I__8324\ : CascadeMux
    port map (
            O => \N__37606\,
            I => \N__37600\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__37603\,
            I => \N__37597\
        );

    \I__8322\ : InMux
    port map (
            O => \N__37600\,
            I => \N__37594\
        );

    \I__8321\ : Span12Mux_v
    port map (
            O => \N__37597\,
            I => \N__37591\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__37594\,
            I => data_idxvec_14
        );

    \I__8319\ : Odrv12
    port map (
            O => \N__37591\,
            I => data_idxvec_14
        );

    \I__8318\ : InMux
    port map (
            O => \N__37586\,
            I => n14053
        );

    \I__8317\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37579\
        );

    \I__8316\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37576\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__37579\,
            I => \N__37573\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__37576\,
            I => \N__37570\
        );

    \I__8313\ : Span4Mux_h
    port map (
            O => \N__37573\,
            I => \N__37567\
        );

    \I__8312\ : Span12Mux_h
    port map (
            O => \N__37570\,
            I => \N__37564\
        );

    \I__8311\ : Odrv4
    port map (
            O => \N__37567\,
            I => n14_adj_1205
        );

    \I__8310\ : Odrv12
    port map (
            O => \N__37564\,
            I => n14_adj_1205
        );

    \I__8309\ : InMux
    port map (
            O => \N__37559\,
            I => n14054
        );

    \I__8308\ : CEMux
    port map (
            O => \N__37556\,
            I => \N__37553\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__37553\,
            I => \N__37549\
        );

    \I__8306\ : CEMux
    port map (
            O => \N__37552\,
            I => \N__37546\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__37549\,
            I => \N__37542\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__37546\,
            I => \N__37539\
        );

    \I__8303\ : CEMux
    port map (
            O => \N__37545\,
            I => \N__37536\
        );

    \I__8302\ : Sp12to4
    port map (
            O => \N__37542\,
            I => \N__37533\
        );

    \I__8301\ : Span4Mux_h
    port map (
            O => \N__37539\,
            I => \N__37530\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__37536\,
            I => \N__37527\
        );

    \I__8299\ : Odrv12
    port map (
            O => \N__37533\,
            I => n9187
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__37530\,
            I => n9187
        );

    \I__8297\ : Odrv12
    port map (
            O => \N__37527\,
            I => n9187
        );

    \I__8296\ : InMux
    port map (
            O => \N__37520\,
            I => \N__37517\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__37517\,
            I => \N__37513\
        );

    \I__8294\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37509\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__37513\,
            I => \N__37506\
        );

    \I__8292\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37503\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__37509\,
            I => buf_adcdata3_13
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__37506\,
            I => buf_adcdata3_13
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__37503\,
            I => buf_adcdata3_13
        );

    \I__8288\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37493\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__37493\,
            I => \N__37489\
        );

    \I__8286\ : InMux
    port map (
            O => \N__37492\,
            I => \N__37486\
        );

    \I__8285\ : Span4Mux_v
    port map (
            O => \N__37489\,
            I => \N__37481\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__37486\,
            I => \N__37481\
        );

    \I__8283\ : Span4Mux_v
    port map (
            O => \N__37481\,
            I => \N__37478\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__37478\,
            I => n14_adj_1198
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__37475\,
            I => \N__37472\
        );

    \I__8280\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37469\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37466\
        );

    \I__8278\ : Span4Mux_v
    port map (
            O => \N__37466\,
            I => \N__37463\
        );

    \I__8277\ : Sp12to4
    port map (
            O => \N__37463\,
            I => \N__37458\
        );

    \I__8276\ : InMux
    port map (
            O => \N__37462\,
            I => \N__37453\
        );

    \I__8275\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37453\
        );

    \I__8274\ : Span12Mux_h
    port map (
            O => \N__37458\,
            I => \N__37450\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__37453\,
            I => cmd_rdadctmp_22
        );

    \I__8272\ : Odrv12
    port map (
            O => \N__37450\,
            I => cmd_rdadctmp_22
        );

    \I__8271\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37442\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__37442\,
            I => \N__37438\
        );

    \I__8269\ : InMux
    port map (
            O => \N__37441\,
            I => \N__37435\
        );

    \I__8268\ : Span4Mux_h
    port map (
            O => \N__37438\,
            I => \N__37432\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__37435\,
            I => buf_adcdata1_14
        );

    \I__8266\ : Odrv4
    port map (
            O => \N__37432\,
            I => buf_adcdata1_14
        );

    \I__8265\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37424\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37419\
        );

    \I__8263\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37416\
        );

    \I__8262\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37413\
        );

    \I__8261\ : Span4Mux_v
    port map (
            O => \N__37419\,
            I => \N__37408\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__37416\,
            I => \N__37408\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__37413\,
            I => req_data_cnt_11
        );

    \I__8258\ : Odrv4
    port map (
            O => \N__37408\,
            I => req_data_cnt_11
        );

    \I__8257\ : InMux
    port map (
            O => \N__37403\,
            I => n14042
        );

    \I__8256\ : InMux
    port map (
            O => \N__37400\,
            I => \N__37396\
        );

    \I__8255\ : InMux
    port map (
            O => \N__37399\,
            I => \N__37393\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__37396\,
            I => \N__37390\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__37393\,
            I => \N__37387\
        );

    \I__8252\ : Span4Mux_h
    port map (
            O => \N__37390\,
            I => \N__37384\
        );

    \I__8251\ : Span4Mux_v
    port map (
            O => \N__37387\,
            I => \N__37381\
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__37384\,
            I => n14_adj_1196
        );

    \I__8249\ : Odrv4
    port map (
            O => \N__37381\,
            I => n14_adj_1196
        );

    \I__8248\ : InMux
    port map (
            O => \N__37376\,
            I => n14043
        );

    \I__8247\ : InMux
    port map (
            O => \N__37373\,
            I => \N__37370\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__37370\,
            I => \N__37366\
        );

    \I__8245\ : InMux
    port map (
            O => \N__37369\,
            I => \N__37363\
        );

    \I__8244\ : Span4Mux_h
    port map (
            O => \N__37366\,
            I => \N__37360\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__37363\,
            I => \N__37357\
        );

    \I__8242\ : Span4Mux_v
    port map (
            O => \N__37360\,
            I => \N__37354\
        );

    \I__8241\ : Odrv4
    port map (
            O => \N__37357\,
            I => n14_adj_1213
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__37354\,
            I => n14_adj_1213
        );

    \I__8239\ : InMux
    port map (
            O => \N__37349\,
            I => n14044
        );

    \I__8238\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37342\
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__37345\,
            I => \N__37339\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__37342\,
            I => \N__37336\
        );

    \I__8235\ : InMux
    port map (
            O => \N__37339\,
            I => \N__37333\
        );

    \I__8234\ : Span4Mux_h
    port map (
            O => \N__37336\,
            I => \N__37330\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__37333\,
            I => data_idxvec_6
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__37330\,
            I => data_idxvec_6
        );

    \I__8231\ : InMux
    port map (
            O => \N__37325\,
            I => n14045
        );

    \I__8230\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37319\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37315\
        );

    \I__8228\ : InMux
    port map (
            O => \N__37318\,
            I => \N__37312\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__37315\,
            I => \N__37309\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__37312\,
            I => \N__37304\
        );

    \I__8225\ : Span4Mux_h
    port map (
            O => \N__37309\,
            I => \N__37304\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__37304\,
            I => \N__37301\
        );

    \I__8223\ : Odrv4
    port map (
            O => \N__37301\,
            I => n14_adj_1168
        );

    \I__8222\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37295\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__37295\,
            I => \N__37291\
        );

    \I__8220\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37288\
        );

    \I__8219\ : Span4Mux_h
    port map (
            O => \N__37291\,
            I => \N__37285\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__37288\,
            I => data_idxvec_7
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__37285\,
            I => data_idxvec_7
        );

    \I__8216\ : InMux
    port map (
            O => \N__37280\,
            I => n14046
        );

    \I__8215\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37274\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__37274\,
            I => \N__37269\
        );

    \I__8213\ : InMux
    port map (
            O => \N__37273\,
            I => \N__37266\
        );

    \I__8212\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37263\
        );

    \I__8211\ : Span4Mux_v
    port map (
            O => \N__37269\,
            I => \N__37260\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__37266\,
            I => \N__37255\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__37263\,
            I => \N__37255\
        );

    \I__8208\ : Span4Mux_h
    port map (
            O => \N__37260\,
            I => \N__37252\
        );

    \I__8207\ : Span4Mux_v
    port map (
            O => \N__37255\,
            I => \N__37249\
        );

    \I__8206\ : Sp12to4
    port map (
            O => \N__37252\,
            I => \N__37246\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__37249\,
            I => n14_adj_1211
        );

    \I__8204\ : Odrv12
    port map (
            O => \N__37246\,
            I => n14_adj_1211
        );

    \I__8203\ : InMux
    port map (
            O => \N__37241\,
            I => \bfn_17_13_0_\
        );

    \I__8202\ : InMux
    port map (
            O => \N__37238\,
            I => \N__37234\
        );

    \I__8201\ : InMux
    port map (
            O => \N__37237\,
            I => \N__37231\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__37234\,
            I => \N__37228\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__37231\,
            I => \N__37225\
        );

    \I__8198\ : Span12Mux_v
    port map (
            O => \N__37228\,
            I => \N__37222\
        );

    \I__8197\ : Span4Mux_v
    port map (
            O => \N__37225\,
            I => \N__37219\
        );

    \I__8196\ : Odrv12
    port map (
            O => \N__37222\,
            I => n14_adj_1210
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__37219\,
            I => n14_adj_1210
        );

    \I__8194\ : CascadeMux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__8193\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37208\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__37208\,
            I => \N__37204\
        );

    \I__8191\ : InMux
    port map (
            O => \N__37207\,
            I => \N__37201\
        );

    \I__8190\ : Span4Mux_h
    port map (
            O => \N__37204\,
            I => \N__37198\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__37201\,
            I => data_idxvec_9
        );

    \I__8188\ : Odrv4
    port map (
            O => \N__37198\,
            I => data_idxvec_9
        );

    \I__8187\ : InMux
    port map (
            O => \N__37193\,
            I => n14048
        );

    \I__8186\ : InMux
    port map (
            O => \N__37190\,
            I => \N__37186\
        );

    \I__8185\ : InMux
    port map (
            O => \N__37189\,
            I => \N__37183\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__37186\,
            I => \N__37180\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__37183\,
            I => \N__37177\
        );

    \I__8182\ : Span4Mux_h
    port map (
            O => \N__37180\,
            I => \N__37172\
        );

    \I__8181\ : Span4Mux_h
    port map (
            O => \N__37177\,
            I => \N__37172\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__37172\,
            I => n14_adj_1209
        );

    \I__8179\ : CascadeMux
    port map (
            O => \N__37169\,
            I => \N__37165\
        );

    \I__8178\ : CascadeMux
    port map (
            O => \N__37168\,
            I => \N__37162\
        );

    \I__8177\ : InMux
    port map (
            O => \N__37165\,
            I => \N__37159\
        );

    \I__8176\ : InMux
    port map (
            O => \N__37162\,
            I => \N__37156\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__37159\,
            I => \N__37153\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__37156\,
            I => data_idxvec_10
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__37153\,
            I => data_idxvec_10
        );

    \I__8172\ : InMux
    port map (
            O => \N__37148\,
            I => n14049
        );

    \I__8171\ : InMux
    port map (
            O => \N__37145\,
            I => \N__37142\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37139\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__37139\,
            I => \N__37136\
        );

    \I__8168\ : Span4Mux_v
    port map (
            O => \N__37136\,
            I => \N__37133\
        );

    \I__8167\ : Span4Mux_h
    port map (
            O => \N__37133\,
            I => \N__37130\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__37130\,
            I => buf_data1_8
        );

    \I__8165\ : CascadeMux
    port map (
            O => \N__37127\,
            I => \n4197_cascade_\
        );

    \I__8164\ : InMux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__8162\ : Span4Mux_h
    port map (
            O => \N__37118\,
            I => \N__37115\
        );

    \I__8161\ : Odrv4
    port map (
            O => \N__37115\,
            I => n4221
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__37112\,
            I => \n4234_cascade_\
        );

    \I__8159\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37106\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__37106\,
            I => \N__37103\
        );

    \I__8157\ : Span4Mux_v
    port map (
            O => \N__37103\,
            I => \N__37100\
        );

    \I__8156\ : Span4Mux_h
    port map (
            O => \N__37100\,
            I => \N__37097\
        );

    \I__8155\ : Span4Mux_h
    port map (
            O => \N__37097\,
            I => \N__37094\
        );

    \I__8154\ : Odrv4
    port map (
            O => \N__37094\,
            I => n4209
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__37091\,
            I => \n4254_cascade_\
        );

    \I__8152\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37085\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__37085\,
            I => n4264
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__37082\,
            I => \n32_cascade_\
        );

    \I__8149\ : InMux
    port map (
            O => \N__37079\,
            I => \N__37076\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__37076\,
            I => \N__37073\
        );

    \I__8147\ : Span4Mux_h
    port map (
            O => \N__37073\,
            I => \N__37070\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__37070\,
            I => \N__37067\
        );

    \I__8145\ : Odrv4
    port map (
            O => \N__37067\,
            I => n15557
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__37064\,
            I => \N__37061\
        );

    \I__8143\ : InMux
    port map (
            O => \N__37061\,
            I => \N__37057\
        );

    \I__8142\ : InMux
    port map (
            O => \N__37060\,
            I => \N__37054\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__37057\,
            I => data_idxvec_0
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__37054\,
            I => data_idxvec_0
        );

    \I__8139\ : InMux
    port map (
            O => \N__37049\,
            I => \N__37046\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__37046\,
            I => \data_idxvec_15_N_673_0\
        );

    \I__8137\ : InMux
    port map (
            O => \N__37043\,
            I => n14040
        );

    \I__8136\ : CascadeMux
    port map (
            O => \N__37040\,
            I => \N__37036\
        );

    \I__8135\ : InMux
    port map (
            O => \N__37039\,
            I => \N__37033\
        );

    \I__8134\ : InMux
    port map (
            O => \N__37036\,
            I => \N__37030\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__37027\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__37030\,
            I => \N__37022\
        );

    \I__8131\ : Span4Mux_v
    port map (
            O => \N__37027\,
            I => \N__37022\
        );

    \I__8130\ : Odrv4
    port map (
            O => \N__37022\,
            I => data_idxvec_2
        );

    \I__8129\ : InMux
    port map (
            O => \N__37019\,
            I => n14041
        );

    \I__8128\ : CascadeMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__8127\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__8125\ : Span4Mux_h
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__8124\ : Span4Mux_v
    port map (
            O => \N__37004\,
            I => \N__37001\
        );

    \I__8123\ : Odrv4
    port map (
            O => \N__37001\,
            I => buf_data1_20
        );

    \I__8122\ : CascadeMux
    port map (
            O => \N__36998\,
            I => \n8058_cascade_\
        );

    \I__8121\ : InMux
    port map (
            O => \N__36995\,
            I => \N__36991\
        );

    \I__8120\ : InMux
    port map (
            O => \N__36994\,
            I => \N__36986\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__36991\,
            I => \N__36983\
        );

    \I__8118\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36980\
        );

    \I__8117\ : CascadeMux
    port map (
            O => \N__36989\,
            I => \N__36977\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__36986\,
            I => \N__36974\
        );

    \I__8115\ : Span4Mux_v
    port map (
            O => \N__36983\,
            I => \N__36969\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__36980\,
            I => \N__36964\
        );

    \I__8113\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36961\
        );

    \I__8112\ : Span4Mux_v
    port map (
            O => \N__36974\,
            I => \N__36957\
        );

    \I__8111\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36954\
        );

    \I__8110\ : CascadeMux
    port map (
            O => \N__36972\,
            I => \N__36951\
        );

    \I__8109\ : Span4Mux_h
    port map (
            O => \N__36969\,
            I => \N__36948\
        );

    \I__8108\ : InMux
    port map (
            O => \N__36968\,
            I => \N__36943\
        );

    \I__8107\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36943\
        );

    \I__8106\ : Span4Mux_v
    port map (
            O => \N__36964\,
            I => \N__36940\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__36961\,
            I => \N__36937\
        );

    \I__8104\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36934\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__36957\,
            I => \N__36929\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__36954\,
            I => \N__36929\
        );

    \I__8101\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36926\
        );

    \I__8100\ : Span4Mux_h
    port map (
            O => \N__36948\,
            I => \N__36923\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__36943\,
            I => \N__36920\
        );

    \I__8098\ : Span4Mux_h
    port map (
            O => \N__36940\,
            I => \N__36915\
        );

    \I__8097\ : Span4Mux_v
    port map (
            O => \N__36937\,
            I => \N__36915\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__36934\,
            I => \N__36908\
        );

    \I__8095\ : Sp12to4
    port map (
            O => \N__36929\,
            I => \N__36908\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__36926\,
            I => \N__36908\
        );

    \I__8093\ : Span4Mux_v
    port map (
            O => \N__36923\,
            I => \N__36903\
        );

    \I__8092\ : Span4Mux_h
    port map (
            O => \N__36920\,
            I => \N__36903\
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__36915\,
            I => comm_buf_0_4
        );

    \I__8090\ : Odrv12
    port map (
            O => \N__36908\,
            I => comm_buf_0_4
        );

    \I__8089\ : Odrv4
    port map (
            O => \N__36903\,
            I => comm_buf_0_4
        );

    \I__8088\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36893\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__36893\,
            I => n15584
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__36890\,
            I => \n83_cascade_\
        );

    \I__8085\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36884\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36881\
        );

    \I__8083\ : Odrv12
    port map (
            O => \N__36881\,
            I => n15581
        );

    \I__8082\ : InMux
    port map (
            O => \N__36878\,
            I => \N__36874\
        );

    \I__8081\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36871\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__36874\,
            I => \N__36868\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36865\
        );

    \I__8078\ : Span4Mux_h
    port map (
            O => \N__36868\,
            I => \N__36862\
        );

    \I__8077\ : Span12Mux_v
    port map (
            O => \N__36865\,
            I => \N__36858\
        );

    \I__8076\ : Span4Mux_h
    port map (
            O => \N__36862\,
            I => \N__36855\
        );

    \I__8075\ : InMux
    port map (
            O => \N__36861\,
            I => \N__36852\
        );

    \I__8074\ : Odrv12
    port map (
            O => \N__36858\,
            I => cmd_rdadctmp_29_adj_1083
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__36855\,
            I => cmd_rdadctmp_29_adj_1083
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__36852\,
            I => cmd_rdadctmp_29_adj_1083
        );

    \I__8071\ : InMux
    port map (
            O => \N__36845\,
            I => \N__36840\
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__36844\,
            I => \N__36837\
        );

    \I__8069\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36834\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N__36831\
        );

    \I__8067\ : InMux
    port map (
            O => \N__36837\,
            I => \N__36828\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__36834\,
            I => \N__36825\
        );

    \I__8065\ : Span4Mux_v
    port map (
            O => \N__36831\,
            I => \N__36822\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36817\
        );

    \I__8063\ : Span4Mux_v
    port map (
            O => \N__36825\,
            I => \N__36817\
        );

    \I__8062\ : Span4Mux_h
    port map (
            O => \N__36822\,
            I => \N__36814\
        );

    \I__8061\ : Sp12to4
    port map (
            O => \N__36817\,
            I => \N__36811\
        );

    \I__8060\ : Odrv4
    port map (
            O => \N__36814\,
            I => buf_adcdata3_21
        );

    \I__8059\ : Odrv12
    port map (
            O => \N__36811\,
            I => buf_adcdata3_21
        );

    \I__8058\ : CascadeMux
    port map (
            O => \N__36806\,
            I => \N__36803\
        );

    \I__8057\ : InMux
    port map (
            O => \N__36803\,
            I => \N__36800\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36797\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__36797\,
            I => \N__36794\
        );

    \I__8054\ : Span4Mux_h
    port map (
            O => \N__36794\,
            I => \N__36790\
        );

    \I__8053\ : CascadeMux
    port map (
            O => \N__36793\,
            I => \N__36786\
        );

    \I__8052\ : Span4Mux_v
    port map (
            O => \N__36790\,
            I => \N__36783\
        );

    \I__8051\ : InMux
    port map (
            O => \N__36789\,
            I => \N__36780\
        );

    \I__8050\ : InMux
    port map (
            O => \N__36786\,
            I => \N__36777\
        );

    \I__8049\ : Odrv4
    port map (
            O => \N__36783\,
            I => cmd_rdadctmp_23_adj_1089
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__36780\,
            I => cmd_rdadctmp_23_adj_1089
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__36777\,
            I => cmd_rdadctmp_23_adj_1089
        );

    \I__8046\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36767\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36764\
        );

    \I__8044\ : Span4Mux_v
    port map (
            O => \N__36764\,
            I => \N__36759\
        );

    \I__8043\ : InMux
    port map (
            O => \N__36763\,
            I => \N__36756\
        );

    \I__8042\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36753\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__36759\,
            I => \N__36748\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__36756\,
            I => \N__36748\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__36753\,
            I => buf_adcdata3_15
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__36748\,
            I => buf_adcdata3_15
        );

    \I__8037\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36740\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__36740\,
            I => \N__36737\
        );

    \I__8035\ : Odrv12
    port map (
            O => \N__36737\,
            I => buf_data1_18
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__36734\,
            I => \N__36731\
        );

    \I__8033\ : InMux
    port map (
            O => \N__36731\,
            I => \N__36728\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__36728\,
            I => \N__36725\
        );

    \I__8031\ : Span4Mux_h
    port map (
            O => \N__36725\,
            I => \N__36722\
        );

    \I__8030\ : Span4Mux_h
    port map (
            O => \N__36722\,
            I => \N__36719\
        );

    \I__8029\ : Odrv4
    port map (
            O => \N__36719\,
            I => n75_adj_1164
        );

    \I__8028\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36709\
        );

    \I__8027\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36706\
        );

    \I__8026\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36702\
        );

    \I__8025\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36699\
        );

    \I__8024\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36696\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__36709\,
            I => \N__36693\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__36706\,
            I => \N__36690\
        );

    \I__8021\ : CascadeMux
    port map (
            O => \N__36705\,
            I => \N__36687\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__36702\,
            I => \N__36684\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__36699\,
            I => \N__36681\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__36696\,
            I => \N__36678\
        );

    \I__8017\ : Span4Mux_h
    port map (
            O => \N__36693\,
            I => \N__36673\
        );

    \I__8016\ : Span4Mux_h
    port map (
            O => \N__36690\,
            I => \N__36673\
        );

    \I__8015\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36670\
        );

    \I__8014\ : Span4Mux_v
    port map (
            O => \N__36684\,
            I => \N__36667\
        );

    \I__8013\ : Span4Mux_v
    port map (
            O => \N__36681\,
            I => \N__36662\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__36678\,
            I => \N__36662\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__36673\,
            I => comm_buf_1_0
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__36670\,
            I => comm_buf_1_0
        );

    \I__8009\ : Odrv4
    port map (
            O => \N__36667\,
            I => comm_buf_1_0
        );

    \I__8008\ : Odrv4
    port map (
            O => \N__36662\,
            I => comm_buf_1_0
        );

    \I__8007\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36650\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__36650\,
            I => \N__36645\
        );

    \I__8005\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36642\
        );

    \I__8004\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36639\
        );

    \I__8003\ : Span4Mux_v
    port map (
            O => \N__36645\,
            I => \N__36636\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__36642\,
            I => data_cntvec_0
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__36639\,
            I => data_cntvec_0
        );

    \I__8000\ : Odrv4
    port map (
            O => \N__36636\,
            I => data_cntvec_0
        );

    \I__7999\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36626\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__36626\,
            I => \N__36623\
        );

    \I__7997\ : Odrv4
    port map (
            O => \N__36623\,
            I => n15527
        );

    \I__7996\ : CEMux
    port map (
            O => \N__36620\,
            I => \N__36617\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__36617\,
            I => \N__36614\
        );

    \I__7994\ : Span4Mux_h
    port map (
            O => \N__36614\,
            I => \N__36611\
        );

    \I__7993\ : Span4Mux_h
    port map (
            O => \N__36611\,
            I => \N__36608\
        );

    \I__7992\ : Odrv4
    port map (
            O => \N__36608\,
            I => n14_adj_1189
        );

    \I__7991\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36602\
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__36602\,
            I => n13_adj_1032
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__36599\,
            I => \n13_adj_1032_cascade_\
        );

    \I__7988\ : InMux
    port map (
            O => \N__36596\,
            I => \N__36590\
        );

    \I__7987\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36590\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__36590\,
            I => n8519
        );

    \I__7985\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36583\
        );

    \I__7984\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36580\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__36583\,
            I => \N__36577\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__36580\,
            I => \N__36574\
        );

    \I__7981\ : Span12Mux_h
    port map (
            O => \N__36577\,
            I => \N__36571\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__36574\,
            I => n22_adj_1115
        );

    \I__7979\ : Odrv12
    port map (
            O => \N__36571\,
            I => n22_adj_1115
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__36566\,
            I => \N__36563\
        );

    \I__7977\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36560\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__36560\,
            I => n15651
        );

    \I__7975\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36554\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__36554\,
            I => n15526
        );

    \I__7973\ : CascadeMux
    port map (
            O => \N__36551\,
            I => \n15668_cascade_\
        );

    \I__7972\ : InMux
    port map (
            O => \N__36548\,
            I => \N__36545\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__36545\,
            I => n1523
        );

    \I__7970\ : CascadeMux
    port map (
            O => \N__36542\,
            I => \n1523_cascade_\
        );

    \I__7969\ : CascadeMux
    port map (
            O => \N__36539\,
            I => \n2_adj_1200_cascade_\
        );

    \I__7968\ : InMux
    port map (
            O => \N__36536\,
            I => \N__36533\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__36533\,
            I => n16464
        );

    \I__7966\ : CascadeMux
    port map (
            O => \N__36530\,
            I => \n16467_cascade_\
        );

    \I__7965\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36524\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__36524\,
            I => n8_adj_1201
        );

    \I__7963\ : SRMux
    port map (
            O => \N__36521\,
            I => \N__36518\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36515\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__36515\,
            I => \N__36512\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__36512\,
            I => \ADC_VAC2.n14926\
        );

    \I__7959\ : InMux
    port map (
            O => \N__36509\,
            I => \N__36506\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36502\
        );

    \I__7957\ : CEMux
    port map (
            O => \N__36505\,
            I => \N__36499\
        );

    \I__7956\ : Sp12to4
    port map (
            O => \N__36502\,
            I => \N__36496\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__36499\,
            I => \N__36493\
        );

    \I__7954\ : Span12Mux_v
    port map (
            O => \N__36496\,
            I => \N__36490\
        );

    \I__7953\ : Odrv4
    port map (
            O => \N__36493\,
            I => \ADC_VAC2.n9413\
        );

    \I__7952\ : Odrv12
    port map (
            O => \N__36490\,
            I => \ADC_VAC2.n9413\
        );

    \I__7951\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36479\
        );

    \I__7950\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36479\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36476\
        );

    \I__7948\ : Span4Mux_h
    port map (
            O => \N__36476\,
            I => \N__36471\
        );

    \I__7947\ : InMux
    port map (
            O => \N__36475\,
            I => \N__36467\
        );

    \I__7946\ : InMux
    port map (
            O => \N__36474\,
            I => \N__36463\
        );

    \I__7945\ : Span4Mux_h
    port map (
            O => \N__36471\,
            I => \N__36460\
        );

    \I__7944\ : CascadeMux
    port map (
            O => \N__36470\,
            I => \N__36457\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__36467\,
            I => \N__36453\
        );

    \I__7942\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36450\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__36463\,
            I => \N__36446\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__36460\,
            I => \N__36443\
        );

    \I__7939\ : InMux
    port map (
            O => \N__36457\,
            I => \N__36438\
        );

    \I__7938\ : InMux
    port map (
            O => \N__36456\,
            I => \N__36438\
        );

    \I__7937\ : Span4Mux_v
    port map (
            O => \N__36453\,
            I => \N__36435\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__36450\,
            I => \N__36430\
        );

    \I__7935\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36425\
        );

    \I__7934\ : Span4Mux_v
    port map (
            O => \N__36446\,
            I => \N__36416\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__36443\,
            I => \N__36416\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__36438\,
            I => \N__36416\
        );

    \I__7931\ : Span4Mux_h
    port map (
            O => \N__36435\,
            I => \N__36416\
        );

    \I__7930\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36411\
        );

    \I__7929\ : InMux
    port map (
            O => \N__36433\,
            I => \N__36411\
        );

    \I__7928\ : Span4Mux_h
    port map (
            O => \N__36430\,
            I => \N__36407\
        );

    \I__7927\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36404\
        );

    \I__7926\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36401\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__36425\,
            I => \N__36398\
        );

    \I__7924\ : Sp12to4
    port map (
            O => \N__36416\,
            I => \N__36393\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__36411\,
            I => \N__36393\
        );

    \I__7922\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36390\
        );

    \I__7921\ : Odrv4
    port map (
            O => \N__36407\,
            I => \DTRIG_N_957_adj_1077\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__36404\,
            I => \DTRIG_N_957_adj_1077\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__36401\,
            I => \DTRIG_N_957_adj_1077\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__36398\,
            I => \DTRIG_N_957_adj_1077\
        );

    \I__7917\ : Odrv12
    port map (
            O => \N__36393\,
            I => \DTRIG_N_957_adj_1077\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__36390\,
            I => \DTRIG_N_957_adj_1077\
        );

    \I__7915\ : SRMux
    port map (
            O => \N__36377\,
            I => \N__36374\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__36374\,
            I => \N__36371\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__36371\,
            I => \N__36368\
        );

    \I__7912\ : Span4Mux_h
    port map (
            O => \N__36368\,
            I => \N__36365\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__36365\,
            I => \N__36362\
        );

    \I__7910\ : Odrv4
    port map (
            O => \N__36362\,
            I => \ADC_VAC2.n10706\
        );

    \I__7909\ : InMux
    port map (
            O => \N__36359\,
            I => \N__36352\
        );

    \I__7908\ : InMux
    port map (
            O => \N__36358\,
            I => \N__36352\
        );

    \I__7907\ : InMux
    port map (
            O => \N__36357\,
            I => \N__36349\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__36352\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__36349\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__7904\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36334\
        );

    \I__7903\ : InMux
    port map (
            O => \N__36343\,
            I => \N__36334\
        );

    \I__7902\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36334\
        );

    \I__7901\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36331\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__36334\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__36331\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__36326\,
            I => \N__36323\
        );

    \I__7897\ : InMux
    port map (
            O => \N__36323\,
            I => \N__36310\
        );

    \I__7896\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36310\
        );

    \I__7895\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36310\
        );

    \I__7894\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36310\
        );

    \I__7893\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36307\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__36310\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__36307\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__7890\ : CascadeMux
    port map (
            O => \N__36302\,
            I => \N__36299\
        );

    \I__7889\ : CascadeBuf
    port map (
            O => \N__36299\,
            I => \N__36296\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__36296\,
            I => \N__36293\
        );

    \I__7887\ : CascadeBuf
    port map (
            O => \N__36293\,
            I => \N__36290\
        );

    \I__7886\ : CascadeMux
    port map (
            O => \N__36290\,
            I => \N__36287\
        );

    \I__7885\ : CascadeBuf
    port map (
            O => \N__36287\,
            I => \N__36284\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__36284\,
            I => \N__36281\
        );

    \I__7883\ : CascadeBuf
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__36278\,
            I => \N__36275\
        );

    \I__7881\ : CascadeBuf
    port map (
            O => \N__36275\,
            I => \N__36272\
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__36272\,
            I => \N__36269\
        );

    \I__7879\ : CascadeBuf
    port map (
            O => \N__36269\,
            I => \N__36266\
        );

    \I__7878\ : CascadeMux
    port map (
            O => \N__36266\,
            I => \N__36263\
        );

    \I__7877\ : CascadeBuf
    port map (
            O => \N__36263\,
            I => \N__36259\
        );

    \I__7876\ : CascadeMux
    port map (
            O => \N__36262\,
            I => \N__36256\
        );

    \I__7875\ : CascadeMux
    port map (
            O => \N__36259\,
            I => \N__36253\
        );

    \I__7874\ : CascadeBuf
    port map (
            O => \N__36256\,
            I => \N__36250\
        );

    \I__7873\ : CascadeBuf
    port map (
            O => \N__36253\,
            I => \N__36247\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__36250\,
            I => \N__36244\
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__36247\,
            I => \N__36241\
        );

    \I__7870\ : InMux
    port map (
            O => \N__36244\,
            I => \N__36238\
        );

    \I__7869\ : CascadeBuf
    port map (
            O => \N__36241\,
            I => \N__36235\
        );

    \I__7868\ : LocalMux
    port map (
            O => \N__36238\,
            I => \N__36232\
        );

    \I__7867\ : CascadeMux
    port map (
            O => \N__36235\,
            I => \N__36229\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__36232\,
            I => \N__36226\
        );

    \I__7865\ : InMux
    port map (
            O => \N__36229\,
            I => \N__36223\
        );

    \I__7864\ : Span4Mux_v
    port map (
            O => \N__36226\,
            I => \N__36220\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__36223\,
            I => \N__36217\
        );

    \I__7862\ : Sp12to4
    port map (
            O => \N__36220\,
            I => \N__36213\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__36217\,
            I => \N__36210\
        );

    \I__7860\ : InMux
    port map (
            O => \N__36216\,
            I => \N__36207\
        );

    \I__7859\ : Span12Mux_v
    port map (
            O => \N__36213\,
            I => \N__36204\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__36210\,
            I => \N__36201\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__36207\,
            I => data_count_4
        );

    \I__7856\ : Odrv12
    port map (
            O => \N__36204\,
            I => data_count_4
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__36201\,
            I => data_count_4
        );

    \I__7854\ : InMux
    port map (
            O => \N__36194\,
            I => n13945
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__36191\,
            I => \N__36188\
        );

    \I__7852\ : CascadeBuf
    port map (
            O => \N__36188\,
            I => \N__36185\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__36185\,
            I => \N__36182\
        );

    \I__7850\ : CascadeBuf
    port map (
            O => \N__36182\,
            I => \N__36179\
        );

    \I__7849\ : CascadeMux
    port map (
            O => \N__36179\,
            I => \N__36176\
        );

    \I__7848\ : CascadeBuf
    port map (
            O => \N__36176\,
            I => \N__36173\
        );

    \I__7847\ : CascadeMux
    port map (
            O => \N__36173\,
            I => \N__36170\
        );

    \I__7846\ : CascadeBuf
    port map (
            O => \N__36170\,
            I => \N__36167\
        );

    \I__7845\ : CascadeMux
    port map (
            O => \N__36167\,
            I => \N__36164\
        );

    \I__7844\ : CascadeBuf
    port map (
            O => \N__36164\,
            I => \N__36161\
        );

    \I__7843\ : CascadeMux
    port map (
            O => \N__36161\,
            I => \N__36158\
        );

    \I__7842\ : CascadeBuf
    port map (
            O => \N__36158\,
            I => \N__36155\
        );

    \I__7841\ : CascadeMux
    port map (
            O => \N__36155\,
            I => \N__36152\
        );

    \I__7840\ : CascadeBuf
    port map (
            O => \N__36152\,
            I => \N__36149\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__36149\,
            I => \N__36145\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__36148\,
            I => \N__36142\
        );

    \I__7837\ : CascadeBuf
    port map (
            O => \N__36145\,
            I => \N__36139\
        );

    \I__7836\ : CascadeBuf
    port map (
            O => \N__36142\,
            I => \N__36136\
        );

    \I__7835\ : CascadeMux
    port map (
            O => \N__36139\,
            I => \N__36133\
        );

    \I__7834\ : CascadeMux
    port map (
            O => \N__36136\,
            I => \N__36130\
        );

    \I__7833\ : CascadeBuf
    port map (
            O => \N__36133\,
            I => \N__36127\
        );

    \I__7832\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36124\
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__36127\,
            I => \N__36121\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__36124\,
            I => \N__36118\
        );

    \I__7829\ : InMux
    port map (
            O => \N__36121\,
            I => \N__36115\
        );

    \I__7828\ : Span4Mux_v
    port map (
            O => \N__36118\,
            I => \N__36112\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36109\
        );

    \I__7826\ : Sp12to4
    port map (
            O => \N__36112\,
            I => \N__36105\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__36109\,
            I => \N__36102\
        );

    \I__7824\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36099\
        );

    \I__7823\ : Span12Mux_h
    port map (
            O => \N__36105\,
            I => \N__36096\
        );

    \I__7822\ : Span4Mux_h
    port map (
            O => \N__36102\,
            I => \N__36093\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__36099\,
            I => data_count_5
        );

    \I__7820\ : Odrv12
    port map (
            O => \N__36096\,
            I => data_count_5
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__36093\,
            I => data_count_5
        );

    \I__7818\ : InMux
    port map (
            O => \N__36086\,
            I => n13946
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__36083\,
            I => \N__36080\
        );

    \I__7816\ : CascadeBuf
    port map (
            O => \N__36080\,
            I => \N__36077\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__36077\,
            I => \N__36074\
        );

    \I__7814\ : CascadeBuf
    port map (
            O => \N__36074\,
            I => \N__36071\
        );

    \I__7813\ : CascadeMux
    port map (
            O => \N__36071\,
            I => \N__36068\
        );

    \I__7812\ : CascadeBuf
    port map (
            O => \N__36068\,
            I => \N__36065\
        );

    \I__7811\ : CascadeMux
    port map (
            O => \N__36065\,
            I => \N__36062\
        );

    \I__7810\ : CascadeBuf
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__7808\ : CascadeBuf
    port map (
            O => \N__36056\,
            I => \N__36053\
        );

    \I__7807\ : CascadeMux
    port map (
            O => \N__36053\,
            I => \N__36050\
        );

    \I__7806\ : CascadeBuf
    port map (
            O => \N__36050\,
            I => \N__36047\
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__36047\,
            I => \N__36044\
        );

    \I__7804\ : CascadeBuf
    port map (
            O => \N__36044\,
            I => \N__36041\
        );

    \I__7803\ : CascadeMux
    port map (
            O => \N__36041\,
            I => \N__36037\
        );

    \I__7802\ : CascadeMux
    port map (
            O => \N__36040\,
            I => \N__36034\
        );

    \I__7801\ : CascadeBuf
    port map (
            O => \N__36037\,
            I => \N__36031\
        );

    \I__7800\ : CascadeBuf
    port map (
            O => \N__36034\,
            I => \N__36028\
        );

    \I__7799\ : CascadeMux
    port map (
            O => \N__36031\,
            I => \N__36025\
        );

    \I__7798\ : CascadeMux
    port map (
            O => \N__36028\,
            I => \N__36022\
        );

    \I__7797\ : CascadeBuf
    port map (
            O => \N__36025\,
            I => \N__36019\
        );

    \I__7796\ : InMux
    port map (
            O => \N__36022\,
            I => \N__36016\
        );

    \I__7795\ : CascadeMux
    port map (
            O => \N__36019\,
            I => \N__36013\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__36016\,
            I => \N__36010\
        );

    \I__7793\ : InMux
    port map (
            O => \N__36013\,
            I => \N__36007\
        );

    \I__7792\ : Sp12to4
    port map (
            O => \N__36010\,
            I => \N__36004\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__36007\,
            I => \N__36001\
        );

    \I__7790\ : Span12Mux_v
    port map (
            O => \N__36004\,
            I => \N__35997\
        );

    \I__7789\ : Span4Mux_h
    port map (
            O => \N__36001\,
            I => \N__35994\
        );

    \I__7788\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35991\
        );

    \I__7787\ : Span12Mux_h
    port map (
            O => \N__35997\,
            I => \N__35988\
        );

    \I__7786\ : Span4Mux_h
    port map (
            O => \N__35994\,
            I => \N__35985\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__35991\,
            I => data_count_6
        );

    \I__7784\ : Odrv12
    port map (
            O => \N__35988\,
            I => data_count_6
        );

    \I__7783\ : Odrv4
    port map (
            O => \N__35985\,
            I => data_count_6
        );

    \I__7782\ : InMux
    port map (
            O => \N__35978\,
            I => n13947
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__35975\,
            I => \N__35972\
        );

    \I__7780\ : CascadeBuf
    port map (
            O => \N__35972\,
            I => \N__35969\
        );

    \I__7779\ : CascadeMux
    port map (
            O => \N__35969\,
            I => \N__35966\
        );

    \I__7778\ : CascadeBuf
    port map (
            O => \N__35966\,
            I => \N__35963\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__35963\,
            I => \N__35960\
        );

    \I__7776\ : CascadeBuf
    port map (
            O => \N__35960\,
            I => \N__35957\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__35957\,
            I => \N__35954\
        );

    \I__7774\ : CascadeBuf
    port map (
            O => \N__35954\,
            I => \N__35951\
        );

    \I__7773\ : CascadeMux
    port map (
            O => \N__35951\,
            I => \N__35948\
        );

    \I__7772\ : CascadeBuf
    port map (
            O => \N__35948\,
            I => \N__35945\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__35945\,
            I => \N__35942\
        );

    \I__7770\ : CascadeBuf
    port map (
            O => \N__35942\,
            I => \N__35939\
        );

    \I__7769\ : CascadeMux
    port map (
            O => \N__35939\,
            I => \N__35936\
        );

    \I__7768\ : CascadeBuf
    port map (
            O => \N__35936\,
            I => \N__35933\
        );

    \I__7767\ : CascadeMux
    port map (
            O => \N__35933\,
            I => \N__35930\
        );

    \I__7766\ : CascadeBuf
    port map (
            O => \N__35930\,
            I => \N__35926\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__35929\,
            I => \N__35923\
        );

    \I__7764\ : CascadeMux
    port map (
            O => \N__35926\,
            I => \N__35920\
        );

    \I__7763\ : CascadeBuf
    port map (
            O => \N__35923\,
            I => \N__35917\
        );

    \I__7762\ : CascadeBuf
    port map (
            O => \N__35920\,
            I => \N__35914\
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__35917\,
            I => \N__35911\
        );

    \I__7760\ : CascadeMux
    port map (
            O => \N__35914\,
            I => \N__35908\
        );

    \I__7759\ : InMux
    port map (
            O => \N__35911\,
            I => \N__35905\
        );

    \I__7758\ : InMux
    port map (
            O => \N__35908\,
            I => \N__35902\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__35905\,
            I => \N__35899\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__35902\,
            I => \N__35896\
        );

    \I__7755\ : Span12Mux_v
    port map (
            O => \N__35899\,
            I => \N__35892\
        );

    \I__7754\ : Span4Mux_h
    port map (
            O => \N__35896\,
            I => \N__35889\
        );

    \I__7753\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35886\
        );

    \I__7752\ : Span12Mux_h
    port map (
            O => \N__35892\,
            I => \N__35883\
        );

    \I__7751\ : Span4Mux_h
    port map (
            O => \N__35889\,
            I => \N__35880\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__35886\,
            I => data_count_7
        );

    \I__7749\ : Odrv12
    port map (
            O => \N__35883\,
            I => data_count_7
        );

    \I__7748\ : Odrv4
    port map (
            O => \N__35880\,
            I => data_count_7
        );

    \I__7747\ : InMux
    port map (
            O => \N__35873\,
            I => n13948
        );

    \I__7746\ : InMux
    port map (
            O => \N__35870\,
            I => \bfn_16_19_0_\
        );

    \I__7745\ : CascadeMux
    port map (
            O => \N__35867\,
            I => \N__35864\
        );

    \I__7744\ : CascadeBuf
    port map (
            O => \N__35864\,
            I => \N__35861\
        );

    \I__7743\ : CascadeMux
    port map (
            O => \N__35861\,
            I => \N__35858\
        );

    \I__7742\ : CascadeBuf
    port map (
            O => \N__35858\,
            I => \N__35855\
        );

    \I__7741\ : CascadeMux
    port map (
            O => \N__35855\,
            I => \N__35852\
        );

    \I__7740\ : CascadeBuf
    port map (
            O => \N__35852\,
            I => \N__35849\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__35849\,
            I => \N__35846\
        );

    \I__7738\ : CascadeBuf
    port map (
            O => \N__35846\,
            I => \N__35843\
        );

    \I__7737\ : CascadeMux
    port map (
            O => \N__35843\,
            I => \N__35840\
        );

    \I__7736\ : CascadeBuf
    port map (
            O => \N__35840\,
            I => \N__35837\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__35837\,
            I => \N__35834\
        );

    \I__7734\ : CascadeBuf
    port map (
            O => \N__35834\,
            I => \N__35831\
        );

    \I__7733\ : CascadeMux
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__7732\ : CascadeBuf
    port map (
            O => \N__35828\,
            I => \N__35825\
        );

    \I__7731\ : CascadeMux
    port map (
            O => \N__35825\,
            I => \N__35822\
        );

    \I__7730\ : CascadeBuf
    port map (
            O => \N__35822\,
            I => \N__35818\
        );

    \I__7729\ : CascadeMux
    port map (
            O => \N__35821\,
            I => \N__35815\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__35818\,
            I => \N__35812\
        );

    \I__7727\ : CascadeBuf
    port map (
            O => \N__35815\,
            I => \N__35809\
        );

    \I__7726\ : CascadeBuf
    port map (
            O => \N__35812\,
            I => \N__35806\
        );

    \I__7725\ : CascadeMux
    port map (
            O => \N__35809\,
            I => \N__35803\
        );

    \I__7724\ : CascadeMux
    port map (
            O => \N__35806\,
            I => \N__35800\
        );

    \I__7723\ : InMux
    port map (
            O => \N__35803\,
            I => \N__35797\
        );

    \I__7722\ : InMux
    port map (
            O => \N__35800\,
            I => \N__35794\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__35797\,
            I => \N__35791\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__35794\,
            I => \N__35788\
        );

    \I__7719\ : Span12Mux_v
    port map (
            O => \N__35791\,
            I => \N__35784\
        );

    \I__7718\ : Span4Mux_h
    port map (
            O => \N__35788\,
            I => \N__35781\
        );

    \I__7717\ : InMux
    port map (
            O => \N__35787\,
            I => \N__35778\
        );

    \I__7716\ : Span12Mux_h
    port map (
            O => \N__35784\,
            I => \N__35775\
        );

    \I__7715\ : Span4Mux_h
    port map (
            O => \N__35781\,
            I => \N__35772\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__35778\,
            I => data_count_8
        );

    \I__7713\ : Odrv12
    port map (
            O => \N__35775\,
            I => data_count_8
        );

    \I__7712\ : Odrv4
    port map (
            O => \N__35772\,
            I => data_count_8
        );

    \I__7711\ : InMux
    port map (
            O => \N__35765\,
            I => \N__35760\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__35764\,
            I => \N__35756\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__35763\,
            I => \N__35749\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__35760\,
            I => \N__35743\
        );

    \I__7707\ : CascadeMux
    port map (
            O => \N__35759\,
            I => \N__35738\
        );

    \I__7706\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35711\
        );

    \I__7705\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35711\
        );

    \I__7704\ : InMux
    port map (
            O => \N__35754\,
            I => \N__35711\
        );

    \I__7703\ : InMux
    port map (
            O => \N__35753\,
            I => \N__35711\
        );

    \I__7702\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35711\
        );

    \I__7701\ : InMux
    port map (
            O => \N__35749\,
            I => \N__35711\
        );

    \I__7700\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35711\
        );

    \I__7699\ : InMux
    port map (
            O => \N__35747\,
            I => \N__35711\
        );

    \I__7698\ : InMux
    port map (
            O => \N__35746\,
            I => \N__35708\
        );

    \I__7697\ : Span4Mux_h
    port map (
            O => \N__35743\,
            I => \N__35705\
        );

    \I__7696\ : InMux
    port map (
            O => \N__35742\,
            I => \N__35688\
        );

    \I__7695\ : InMux
    port map (
            O => \N__35741\,
            I => \N__35688\
        );

    \I__7694\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35688\
        );

    \I__7693\ : InMux
    port map (
            O => \N__35737\,
            I => \N__35688\
        );

    \I__7692\ : InMux
    port map (
            O => \N__35736\,
            I => \N__35688\
        );

    \I__7691\ : InMux
    port map (
            O => \N__35735\,
            I => \N__35688\
        );

    \I__7690\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35688\
        );

    \I__7689\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35688\
        );

    \I__7688\ : InMux
    port map (
            O => \N__35732\,
            I => \N__35677\
        );

    \I__7687\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35677\
        );

    \I__7686\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35677\
        );

    \I__7685\ : InMux
    port map (
            O => \N__35729\,
            I => \N__35677\
        );

    \I__7684\ : InMux
    port map (
            O => \N__35728\,
            I => \N__35677\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__35711\,
            I => \N__35674\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__35708\,
            I => \N__35671\
        );

    \I__7681\ : Span4Mux_h
    port map (
            O => \N__35705\,
            I => \N__35662\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__35688\,
            I => \N__35662\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__35677\,
            I => \N__35662\
        );

    \I__7678\ : Span12Mux_v
    port map (
            O => \N__35674\,
            I => \N__35659\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__35671\,
            I => \N__35656\
        );

    \I__7676\ : InMux
    port map (
            O => \N__35670\,
            I => \N__35653\
        );

    \I__7675\ : InMux
    port map (
            O => \N__35669\,
            I => \N__35650\
        );

    \I__7674\ : Sp12to4
    port map (
            O => \N__35662\,
            I => \N__35647\
        );

    \I__7673\ : Odrv12
    port map (
            O => \N__35659\,
            I => dds_state_2
        );

    \I__7672\ : Odrv4
    port map (
            O => \N__35656\,
            I => dds_state_2
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__35653\,
            I => dds_state_2
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__35650\,
            I => dds_state_2
        );

    \I__7669\ : Odrv12
    port map (
            O => \N__35647\,
            I => dds_state_2
        );

    \I__7668\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35633\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__35633\,
            I => \N__35630\
        );

    \I__7666\ : Span4Mux_h
    port map (
            O => \N__35630\,
            I => \N__35627\
        );

    \I__7665\ : Span4Mux_v
    port map (
            O => \N__35627\,
            I => \N__35624\
        );

    \I__7664\ : Span4Mux_v
    port map (
            O => \N__35624\,
            I => \N__35621\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__35621\,
            I => \ADC_VAC2.n15280\
        );

    \I__7662\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35613\
        );

    \I__7661\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35610\
        );

    \I__7660\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35605\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__35613\,
            I => \N__35600\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__35610\,
            I => \N__35600\
        );

    \I__7657\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35592\
        );

    \I__7656\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35589\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__35605\,
            I => \N__35586\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__35600\,
            I => \N__35583\
        );

    \I__7653\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35572\
        );

    \I__7652\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35572\
        );

    \I__7651\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35572\
        );

    \I__7650\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35572\
        );

    \I__7649\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35572\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__35592\,
            I => \N__35569\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__35589\,
            I => \N__35565\
        );

    \I__7646\ : Span4Mux_h
    port map (
            O => \N__35586\,
            I => \N__35562\
        );

    \I__7645\ : Span4Mux_h
    port map (
            O => \N__35583\,
            I => \N__35557\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__35572\,
            I => \N__35557\
        );

    \I__7643\ : Span4Mux_v
    port map (
            O => \N__35569\,
            I => \N__35554\
        );

    \I__7642\ : InMux
    port map (
            O => \N__35568\,
            I => \N__35551\
        );

    \I__7641\ : Span12Mux_s8_h
    port map (
            O => \N__35565\,
            I => \N__35546\
        );

    \I__7640\ : Sp12to4
    port map (
            O => \N__35562\,
            I => \N__35546\
        );

    \I__7639\ : Span4Mux_h
    port map (
            O => \N__35557\,
            I => \N__35543\
        );

    \I__7638\ : Sp12to4
    port map (
            O => \N__35554\,
            I => \N__35540\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__35551\,
            I => \N__35536\
        );

    \I__7636\ : Span12Mux_v
    port map (
            O => \N__35546\,
            I => \N__35533\
        );

    \I__7635\ : Span4Mux_h
    port map (
            O => \N__35543\,
            I => \N__35530\
        );

    \I__7634\ : Span12Mux_h
    port map (
            O => \N__35540\,
            I => \N__35527\
        );

    \I__7633\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35524\
        );

    \I__7632\ : Span12Mux_h
    port map (
            O => \N__35536\,
            I => \N__35517\
        );

    \I__7631\ : Span12Mux_h
    port map (
            O => \N__35533\,
            I => \N__35517\
        );

    \I__7630\ : Sp12to4
    port map (
            O => \N__35530\,
            I => \N__35517\
        );

    \I__7629\ : Odrv12
    port map (
            O => \N__35527\,
            I => adc_state_1_adj_1043
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__35524\,
            I => adc_state_1_adj_1043
        );

    \I__7627\ : Odrv12
    port map (
            O => \N__35517\,
            I => adc_state_1_adj_1043
        );

    \I__7626\ : CEMux
    port map (
            O => \N__35510\,
            I => \N__35507\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__35507\,
            I => \N__35504\
        );

    \I__7624\ : Span4Mux_h
    port map (
            O => \N__35504\,
            I => \N__35500\
        );

    \I__7623\ : CEMux
    port map (
            O => \N__35503\,
            I => \N__35497\
        );

    \I__7622\ : Span4Mux_v
    port map (
            O => \N__35500\,
            I => \N__35494\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__35497\,
            I => \N__35491\
        );

    \I__7620\ : Span4Mux_v
    port map (
            O => \N__35494\,
            I => \N__35488\
        );

    \I__7619\ : Span4Mux_h
    port map (
            O => \N__35491\,
            I => \N__35485\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__35488\,
            I => \N__35480\
        );

    \I__7617\ : Span4Mux_h
    port map (
            O => \N__35485\,
            I => \N__35480\
        );

    \I__7616\ : Odrv4
    port map (
            O => \N__35480\,
            I => \ADC_VAC2.n12\
        );

    \I__7615\ : CascadeMux
    port map (
            O => \N__35477\,
            I => \N__35474\
        );

    \I__7614\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35471\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35467\
        );

    \I__7612\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35464\
        );

    \I__7611\ : Span4Mux_h
    port map (
            O => \N__35467\,
            I => \N__35461\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__35464\,
            I => data_cntvec_12
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__35461\,
            I => data_cntvec_12
        );

    \I__7608\ : InMux
    port map (
            O => \N__35456\,
            I => n13962
        );

    \I__7607\ : CascadeMux
    port map (
            O => \N__35453\,
            I => \N__35450\
        );

    \I__7606\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35447\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__35447\,
            I => \N__35443\
        );

    \I__7604\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35440\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__35443\,
            I => \N__35437\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__35440\,
            I => data_cntvec_13
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__35437\,
            I => data_cntvec_13
        );

    \I__7600\ : InMux
    port map (
            O => \N__35432\,
            I => n13963
        );

    \I__7599\ : CascadeMux
    port map (
            O => \N__35429\,
            I => \N__35426\
        );

    \I__7598\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35423\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__35423\,
            I => \N__35419\
        );

    \I__7596\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35416\
        );

    \I__7595\ : Span4Mux_h
    port map (
            O => \N__35419\,
            I => \N__35413\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__35416\,
            I => data_cntvec_14
        );

    \I__7593\ : Odrv4
    port map (
            O => \N__35413\,
            I => data_cntvec_14
        );

    \I__7592\ : InMux
    port map (
            O => \N__35408\,
            I => n13964
        );

    \I__7591\ : InMux
    port map (
            O => \N__35405\,
            I => n13965
        );

    \I__7590\ : CascadeMux
    port map (
            O => \N__35402\,
            I => \N__35399\
        );

    \I__7589\ : InMux
    port map (
            O => \N__35399\,
            I => \N__35396\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__35396\,
            I => \N__35392\
        );

    \I__7587\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35389\
        );

    \I__7586\ : Span4Mux_h
    port map (
            O => \N__35392\,
            I => \N__35386\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__35389\,
            I => \N__35381\
        );

    \I__7584\ : Span4Mux_v
    port map (
            O => \N__35386\,
            I => \N__35381\
        );

    \I__7583\ : Odrv4
    port map (
            O => \N__35381\,
            I => data_cntvec_15
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__35378\,
            I => \N__35375\
        );

    \I__7581\ : CascadeBuf
    port map (
            O => \N__35375\,
            I => \N__35372\
        );

    \I__7580\ : CascadeMux
    port map (
            O => \N__35372\,
            I => \N__35369\
        );

    \I__7579\ : CascadeBuf
    port map (
            O => \N__35369\,
            I => \N__35366\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__35366\,
            I => \N__35363\
        );

    \I__7577\ : CascadeBuf
    port map (
            O => \N__35363\,
            I => \N__35360\
        );

    \I__7576\ : CascadeMux
    port map (
            O => \N__35360\,
            I => \N__35357\
        );

    \I__7575\ : CascadeBuf
    port map (
            O => \N__35357\,
            I => \N__35354\
        );

    \I__7574\ : CascadeMux
    port map (
            O => \N__35354\,
            I => \N__35351\
        );

    \I__7573\ : CascadeBuf
    port map (
            O => \N__35351\,
            I => \N__35348\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__35348\,
            I => \N__35345\
        );

    \I__7571\ : CascadeBuf
    port map (
            O => \N__35345\,
            I => \N__35342\
        );

    \I__7570\ : CascadeMux
    port map (
            O => \N__35342\,
            I => \N__35339\
        );

    \I__7569\ : CascadeBuf
    port map (
            O => \N__35339\,
            I => \N__35336\
        );

    \I__7568\ : CascadeMux
    port map (
            O => \N__35336\,
            I => \N__35333\
        );

    \I__7567\ : CascadeBuf
    port map (
            O => \N__35333\,
            I => \N__35329\
        );

    \I__7566\ : CascadeMux
    port map (
            O => \N__35332\,
            I => \N__35326\
        );

    \I__7565\ : CascadeMux
    port map (
            O => \N__35329\,
            I => \N__35323\
        );

    \I__7564\ : CascadeBuf
    port map (
            O => \N__35326\,
            I => \N__35320\
        );

    \I__7563\ : CascadeBuf
    port map (
            O => \N__35323\,
            I => \N__35317\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__35320\,
            I => \N__35314\
        );

    \I__7561\ : CascadeMux
    port map (
            O => \N__35317\,
            I => \N__35311\
        );

    \I__7560\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35308\
        );

    \I__7559\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35305\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__35308\,
            I => \N__35302\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__35305\,
            I => \N__35299\
        );

    \I__7556\ : Span12Mux_v
    port map (
            O => \N__35302\,
            I => \N__35295\
        );

    \I__7555\ : Span4Mux_h
    port map (
            O => \N__35299\,
            I => \N__35292\
        );

    \I__7554\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35289\
        );

    \I__7553\ : Span12Mux_h
    port map (
            O => \N__35295\,
            I => \N__35286\
        );

    \I__7552\ : Span4Mux_h
    port map (
            O => \N__35292\,
            I => \N__35283\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__35289\,
            I => data_count_0
        );

    \I__7550\ : Odrv12
    port map (
            O => \N__35286\,
            I => data_count_0
        );

    \I__7549\ : Odrv4
    port map (
            O => \N__35283\,
            I => data_count_0
        );

    \I__7548\ : InMux
    port map (
            O => \N__35276\,
            I => \bfn_16_18_0_\
        );

    \I__7547\ : CascadeMux
    port map (
            O => \N__35273\,
            I => \N__35270\
        );

    \I__7546\ : CascadeBuf
    port map (
            O => \N__35270\,
            I => \N__35267\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__35267\,
            I => \N__35264\
        );

    \I__7544\ : CascadeBuf
    port map (
            O => \N__35264\,
            I => \N__35261\
        );

    \I__7543\ : CascadeMux
    port map (
            O => \N__35261\,
            I => \N__35258\
        );

    \I__7542\ : CascadeBuf
    port map (
            O => \N__35258\,
            I => \N__35255\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__35255\,
            I => \N__35252\
        );

    \I__7540\ : CascadeBuf
    port map (
            O => \N__35252\,
            I => \N__35249\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__35249\,
            I => \N__35246\
        );

    \I__7538\ : CascadeBuf
    port map (
            O => \N__35246\,
            I => \N__35243\
        );

    \I__7537\ : CascadeMux
    port map (
            O => \N__35243\,
            I => \N__35240\
        );

    \I__7536\ : CascadeBuf
    port map (
            O => \N__35240\,
            I => \N__35237\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__35237\,
            I => \N__35234\
        );

    \I__7534\ : CascadeBuf
    port map (
            O => \N__35234\,
            I => \N__35231\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__35231\,
            I => \N__35228\
        );

    \I__7532\ : CascadeBuf
    port map (
            O => \N__35228\,
            I => \N__35224\
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__35227\,
            I => \N__35221\
        );

    \I__7530\ : CascadeMux
    port map (
            O => \N__35224\,
            I => \N__35218\
        );

    \I__7529\ : CascadeBuf
    port map (
            O => \N__35221\,
            I => \N__35215\
        );

    \I__7528\ : CascadeBuf
    port map (
            O => \N__35218\,
            I => \N__35212\
        );

    \I__7527\ : CascadeMux
    port map (
            O => \N__35215\,
            I => \N__35209\
        );

    \I__7526\ : CascadeMux
    port map (
            O => \N__35212\,
            I => \N__35206\
        );

    \I__7525\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35203\
        );

    \I__7524\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35200\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35197\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__35200\,
            I => \N__35194\
        );

    \I__7521\ : Span12Mux_v
    port map (
            O => \N__35197\,
            I => \N__35190\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__35194\,
            I => \N__35187\
        );

    \I__7519\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35184\
        );

    \I__7518\ : Span12Mux_h
    port map (
            O => \N__35190\,
            I => \N__35181\
        );

    \I__7517\ : Span4Mux_h
    port map (
            O => \N__35187\,
            I => \N__35178\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__35184\,
            I => data_count_1
        );

    \I__7515\ : Odrv12
    port map (
            O => \N__35181\,
            I => data_count_1
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__35178\,
            I => data_count_1
        );

    \I__7513\ : InMux
    port map (
            O => \N__35171\,
            I => n13942
        );

    \I__7512\ : CascadeMux
    port map (
            O => \N__35168\,
            I => \N__35165\
        );

    \I__7511\ : CascadeBuf
    port map (
            O => \N__35165\,
            I => \N__35162\
        );

    \I__7510\ : CascadeMux
    port map (
            O => \N__35162\,
            I => \N__35159\
        );

    \I__7509\ : CascadeBuf
    port map (
            O => \N__35159\,
            I => \N__35156\
        );

    \I__7508\ : CascadeMux
    port map (
            O => \N__35156\,
            I => \N__35153\
        );

    \I__7507\ : CascadeBuf
    port map (
            O => \N__35153\,
            I => \N__35150\
        );

    \I__7506\ : CascadeMux
    port map (
            O => \N__35150\,
            I => \N__35147\
        );

    \I__7505\ : CascadeBuf
    port map (
            O => \N__35147\,
            I => \N__35144\
        );

    \I__7504\ : CascadeMux
    port map (
            O => \N__35144\,
            I => \N__35141\
        );

    \I__7503\ : CascadeBuf
    port map (
            O => \N__35141\,
            I => \N__35138\
        );

    \I__7502\ : CascadeMux
    port map (
            O => \N__35138\,
            I => \N__35135\
        );

    \I__7501\ : CascadeBuf
    port map (
            O => \N__35135\,
            I => \N__35132\
        );

    \I__7500\ : CascadeMux
    port map (
            O => \N__35132\,
            I => \N__35129\
        );

    \I__7499\ : CascadeBuf
    port map (
            O => \N__35129\,
            I => \N__35126\
        );

    \I__7498\ : CascadeMux
    port map (
            O => \N__35126\,
            I => \N__35123\
        );

    \I__7497\ : CascadeBuf
    port map (
            O => \N__35123\,
            I => \N__35119\
        );

    \I__7496\ : CascadeMux
    port map (
            O => \N__35122\,
            I => \N__35116\
        );

    \I__7495\ : CascadeMux
    port map (
            O => \N__35119\,
            I => \N__35113\
        );

    \I__7494\ : CascadeBuf
    port map (
            O => \N__35116\,
            I => \N__35110\
        );

    \I__7493\ : CascadeBuf
    port map (
            O => \N__35113\,
            I => \N__35107\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__35110\,
            I => \N__35104\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__35107\,
            I => \N__35101\
        );

    \I__7490\ : InMux
    port map (
            O => \N__35104\,
            I => \N__35098\
        );

    \I__7489\ : InMux
    port map (
            O => \N__35101\,
            I => \N__35095\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__35098\,
            I => \N__35092\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__35095\,
            I => \N__35089\
        );

    \I__7486\ : Span12Mux_v
    port map (
            O => \N__35092\,
            I => \N__35085\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__35089\,
            I => \N__35082\
        );

    \I__7484\ : InMux
    port map (
            O => \N__35088\,
            I => \N__35079\
        );

    \I__7483\ : Span12Mux_h
    port map (
            O => \N__35085\,
            I => \N__35076\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__35082\,
            I => \N__35073\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__35079\,
            I => data_count_2
        );

    \I__7480\ : Odrv12
    port map (
            O => \N__35076\,
            I => data_count_2
        );

    \I__7479\ : Odrv4
    port map (
            O => \N__35073\,
            I => data_count_2
        );

    \I__7478\ : InMux
    port map (
            O => \N__35066\,
            I => n13943
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__35063\,
            I => \N__35060\
        );

    \I__7476\ : CascadeBuf
    port map (
            O => \N__35060\,
            I => \N__35057\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__35057\,
            I => \N__35054\
        );

    \I__7474\ : CascadeBuf
    port map (
            O => \N__35054\,
            I => \N__35051\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__35051\,
            I => \N__35048\
        );

    \I__7472\ : CascadeBuf
    port map (
            O => \N__35048\,
            I => \N__35045\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__35045\,
            I => \N__35042\
        );

    \I__7470\ : CascadeBuf
    port map (
            O => \N__35042\,
            I => \N__35039\
        );

    \I__7469\ : CascadeMux
    port map (
            O => \N__35039\,
            I => \N__35036\
        );

    \I__7468\ : CascadeBuf
    port map (
            O => \N__35036\,
            I => \N__35033\
        );

    \I__7467\ : CascadeMux
    port map (
            O => \N__35033\,
            I => \N__35030\
        );

    \I__7466\ : CascadeBuf
    port map (
            O => \N__35030\,
            I => \N__35027\
        );

    \I__7465\ : CascadeMux
    port map (
            O => \N__35027\,
            I => \N__35024\
        );

    \I__7464\ : CascadeBuf
    port map (
            O => \N__35024\,
            I => \N__35021\
        );

    \I__7463\ : CascadeMux
    port map (
            O => \N__35021\,
            I => \N__35017\
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__35020\,
            I => \N__35014\
        );

    \I__7461\ : CascadeBuf
    port map (
            O => \N__35017\,
            I => \N__35011\
        );

    \I__7460\ : CascadeBuf
    port map (
            O => \N__35014\,
            I => \N__35008\
        );

    \I__7459\ : CascadeMux
    port map (
            O => \N__35011\,
            I => \N__35005\
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__35008\,
            I => \N__35002\
        );

    \I__7457\ : CascadeBuf
    port map (
            O => \N__35005\,
            I => \N__34999\
        );

    \I__7456\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34996\
        );

    \I__7455\ : CascadeMux
    port map (
            O => \N__34999\,
            I => \N__34993\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34990\
        );

    \I__7453\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34987\
        );

    \I__7452\ : Sp12to4
    port map (
            O => \N__34990\,
            I => \N__34984\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34981\
        );

    \I__7450\ : Span12Mux_v
    port map (
            O => \N__34984\,
            I => \N__34977\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__34981\,
            I => \N__34974\
        );

    \I__7448\ : InMux
    port map (
            O => \N__34980\,
            I => \N__34971\
        );

    \I__7447\ : Span12Mux_h
    port map (
            O => \N__34977\,
            I => \N__34968\
        );

    \I__7446\ : Span4Mux_h
    port map (
            O => \N__34974\,
            I => \N__34965\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__34971\,
            I => data_count_3
        );

    \I__7444\ : Odrv12
    port map (
            O => \N__34968\,
            I => data_count_3
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__34965\,
            I => data_count_3
        );

    \I__7442\ : InMux
    port map (
            O => \N__34958\,
            I => n13944
        );

    \I__7441\ : InMux
    port map (
            O => \N__34955\,
            I => n13953
        );

    \I__7440\ : InMux
    port map (
            O => \N__34952\,
            I => n13954
        );

    \I__7439\ : InMux
    port map (
            O => \N__34949\,
            I => n13955
        );

    \I__7438\ : InMux
    port map (
            O => \N__34946\,
            I => \N__34941\
        );

    \I__7437\ : InMux
    port map (
            O => \N__34945\,
            I => \N__34938\
        );

    \I__7436\ : InMux
    port map (
            O => \N__34944\,
            I => \N__34935\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__34941\,
            I => data_cntvec_6
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__34938\,
            I => data_cntvec_6
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__34935\,
            I => data_cntvec_6
        );

    \I__7432\ : InMux
    port map (
            O => \N__34928\,
            I => n13956
        );

    \I__7431\ : InMux
    port map (
            O => \N__34925\,
            I => \N__34922\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__34922\,
            I => \N__34917\
        );

    \I__7429\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34914\
        );

    \I__7428\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34911\
        );

    \I__7427\ : Span4Mux_h
    port map (
            O => \N__34917\,
            I => \N__34908\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__34914\,
            I => \N__34905\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__34911\,
            I => \N__34900\
        );

    \I__7424\ : Span4Mux_v
    port map (
            O => \N__34908\,
            I => \N__34900\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__34905\,
            I => \N__34897\
        );

    \I__7422\ : Odrv4
    port map (
            O => \N__34900\,
            I => data_cntvec_7
        );

    \I__7421\ : Odrv4
    port map (
            O => \N__34897\,
            I => data_cntvec_7
        );

    \I__7420\ : InMux
    port map (
            O => \N__34892\,
            I => n13957
        );

    \I__7419\ : InMux
    port map (
            O => \N__34889\,
            I => \N__34885\
        );

    \I__7418\ : InMux
    port map (
            O => \N__34888\,
            I => \N__34882\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__34885\,
            I => \N__34878\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__34882\,
            I => \N__34875\
        );

    \I__7415\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34872\
        );

    \I__7414\ : Span4Mux_v
    port map (
            O => \N__34878\,
            I => \N__34869\
        );

    \I__7413\ : Span4Mux_h
    port map (
            O => \N__34875\,
            I => \N__34866\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__34872\,
            I => data_cntvec_8
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__34869\,
            I => data_cntvec_8
        );

    \I__7410\ : Odrv4
    port map (
            O => \N__34866\,
            I => data_cntvec_8
        );

    \I__7409\ : InMux
    port map (
            O => \N__34859\,
            I => \bfn_16_17_0_\
        );

    \I__7408\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34852\
        );

    \I__7407\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34849\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__34852\,
            I => \N__34846\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__34849\,
            I => \N__34842\
        );

    \I__7404\ : Span4Mux_h
    port map (
            O => \N__34846\,
            I => \N__34839\
        );

    \I__7403\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34836\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__34842\,
            I => \N__34833\
        );

    \I__7401\ : Span4Mux_v
    port map (
            O => \N__34839\,
            I => \N__34830\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__34836\,
            I => data_cntvec_9
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__34833\,
            I => data_cntvec_9
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__34830\,
            I => data_cntvec_9
        );

    \I__7397\ : InMux
    port map (
            O => \N__34823\,
            I => n13959
        );

    \I__7396\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34816\
        );

    \I__7395\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34813\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34809\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__34813\,
            I => \N__34806\
        );

    \I__7392\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34803\
        );

    \I__7391\ : Span4Mux_h
    port map (
            O => \N__34809\,
            I => \N__34800\
        );

    \I__7390\ : Span12Mux_v
    port map (
            O => \N__34806\,
            I => \N__34797\
        );

    \I__7389\ : LocalMux
    port map (
            O => \N__34803\,
            I => data_cntvec_10
        );

    \I__7388\ : Odrv4
    port map (
            O => \N__34800\,
            I => data_cntvec_10
        );

    \I__7387\ : Odrv12
    port map (
            O => \N__34797\,
            I => data_cntvec_10
        );

    \I__7386\ : InMux
    port map (
            O => \N__34790\,
            I => n13960
        );

    \I__7385\ : InMux
    port map (
            O => \N__34787\,
            I => \N__34783\
        );

    \I__7384\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34779\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__34783\,
            I => \N__34776\
        );

    \I__7382\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34773\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__34779\,
            I => \N__34768\
        );

    \I__7380\ : Span4Mux_h
    port map (
            O => \N__34776\,
            I => \N__34768\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__34773\,
            I => data_cntvec_11
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__34768\,
            I => data_cntvec_11
        );

    \I__7377\ : InMux
    port map (
            O => \N__34763\,
            I => n13961
        );

    \I__7376\ : InMux
    port map (
            O => \N__34760\,
            I => \N__34755\
        );

    \I__7375\ : InMux
    port map (
            O => \N__34759\,
            I => \N__34752\
        );

    \I__7374\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34749\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__34755\,
            I => \N__34746\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__34752\,
            I => \acadc_skipCount_6\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__34749\,
            I => \acadc_skipCount_6\
        );

    \I__7370\ : Odrv4
    port map (
            O => \N__34746\,
            I => \acadc_skipCount_6\
        );

    \I__7369\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34736\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__34736\,
            I => \N__34733\
        );

    \I__7367\ : Span4Mux_h
    port map (
            O => \N__34733\,
            I => \N__34730\
        );

    \I__7366\ : Span4Mux_h
    port map (
            O => \N__34730\,
            I => \N__34727\
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__34727\,
            I => buf_data1_14
        );

    \I__7364\ : CascadeMux
    port map (
            O => \N__34724\,
            I => \n4191_cascade_\
        );

    \I__7363\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34718\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__34718\,
            I => n4215
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__34715\,
            I => \n4228_cascade_\
        );

    \I__7360\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34709\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__34709\,
            I => n4203
        );

    \I__7358\ : CascadeMux
    port map (
            O => \N__34706\,
            I => \n4248_cascade_\
        );

    \I__7357\ : InMux
    port map (
            O => \N__34703\,
            I => \N__34700\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__34700\,
            I => \N__34697\
        );

    \I__7355\ : Odrv12
    port map (
            O => \N__34697\,
            I => n4258
        );

    \I__7354\ : InMux
    port map (
            O => \N__34694\,
            I => \bfn_16_16_0_\
        );

    \I__7353\ : InMux
    port map (
            O => \N__34691\,
            I => n13951
        );

    \I__7352\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34685\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__34685\,
            I => \N__34680\
        );

    \I__7350\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34677\
        );

    \I__7349\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34674\
        );

    \I__7348\ : Span4Mux_h
    port map (
            O => \N__34680\,
            I => \N__34671\
        );

    \I__7347\ : LocalMux
    port map (
            O => \N__34677\,
            I => \N__34668\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__34674\,
            I => data_cntvec_2
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__34671\,
            I => data_cntvec_2
        );

    \I__7344\ : Odrv4
    port map (
            O => \N__34668\,
            I => data_cntvec_2
        );

    \I__7343\ : InMux
    port map (
            O => \N__34661\,
            I => n13952
        );

    \I__7342\ : InMux
    port map (
            O => \N__34658\,
            I => \N__34654\
        );

    \I__7341\ : CascadeMux
    port map (
            O => \N__34657\,
            I => \N__34650\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__34654\,
            I => \N__34647\
        );

    \I__7339\ : InMux
    port map (
            O => \N__34653\,
            I => \N__34644\
        );

    \I__7338\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34641\
        );

    \I__7337\ : Odrv4
    port map (
            O => \N__34647\,
            I => req_data_cnt_4
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__34644\,
            I => req_data_cnt_4
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__34641\,
            I => req_data_cnt_4
        );

    \I__7334\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34631\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__34631\,
            I => n18_adj_1217
        );

    \I__7332\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34625\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__34625\,
            I => \N__34621\
        );

    \I__7330\ : CascadeMux
    port map (
            O => \N__34624\,
            I => \N__34618\
        );

    \I__7329\ : Span4Mux_h
    port map (
            O => \N__34621\,
            I => \N__34614\
        );

    \I__7328\ : InMux
    port map (
            O => \N__34618\,
            I => \N__34611\
        );

    \I__7327\ : InMux
    port map (
            O => \N__34617\,
            I => \N__34608\
        );

    \I__7326\ : Span4Mux_v
    port map (
            O => \N__34614\,
            I => \N__34605\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__34611\,
            I => \N__34602\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__34608\,
            I => buf_dds_6
        );

    \I__7323\ : Odrv4
    port map (
            O => \N__34605\,
            I => buf_dds_6
        );

    \I__7322\ : Odrv12
    port map (
            O => \N__34602\,
            I => buf_dds_6
        );

    \I__7321\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34587\
        );

    \I__7320\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34584\
        );

    \I__7319\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34581\
        );

    \I__7318\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34578\
        );

    \I__7317\ : InMux
    port map (
            O => \N__34591\,
            I => \N__34575\
        );

    \I__7316\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34572\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__34587\,
            I => \N__34567\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__34584\,
            I => \N__34567\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__34581\,
            I => \N__34564\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__34578\,
            I => \N__34561\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34551\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__34572\,
            I => \N__34551\
        );

    \I__7309\ : Span4Mux_h
    port map (
            O => \N__34567\,
            I => \N__34551\
        );

    \I__7308\ : Span4Mux_h
    port map (
            O => \N__34564\,
            I => \N__34551\
        );

    \I__7307\ : Span4Mux_v
    port map (
            O => \N__34561\,
            I => \N__34547\
        );

    \I__7306\ : InMux
    port map (
            O => \N__34560\,
            I => \N__34544\
        );

    \I__7305\ : Span4Mux_h
    port map (
            O => \N__34551\,
            I => \N__34541\
        );

    \I__7304\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34538\
        );

    \I__7303\ : Span4Mux_h
    port map (
            O => \N__34547\,
            I => \N__34535\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34532\
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__34541\,
            I => comm_buf_0_1
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__34538\,
            I => comm_buf_0_1
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__34535\,
            I => comm_buf_0_1
        );

    \I__7298\ : Odrv12
    port map (
            O => \N__34532\,
            I => comm_buf_0_1
        );

    \I__7297\ : InMux
    port map (
            O => \N__34523\,
            I => \N__34520\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__34520\,
            I => \N__34516\
        );

    \I__7295\ : InMux
    port map (
            O => \N__34519\,
            I => \N__34513\
        );

    \I__7294\ : Odrv4
    port map (
            O => \N__34516\,
            I => n7485
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__34513\,
            I => n7485
        );

    \I__7292\ : InMux
    port map (
            O => \N__34508\,
            I => \N__34503\
        );

    \I__7291\ : InMux
    port map (
            O => \N__34507\,
            I => \N__34499\
        );

    \I__7290\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34496\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__34503\,
            I => \N__34493\
        );

    \I__7288\ : InMux
    port map (
            O => \N__34502\,
            I => \N__34490\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__34499\,
            I => \N__34487\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34480\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__34493\,
            I => \N__34480\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__34490\,
            I => \N__34480\
        );

    \I__7283\ : Odrv12
    port map (
            O => \N__34487\,
            I => eis_stop
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__34480\,
            I => eis_stop
        );

    \I__7281\ : InMux
    port map (
            O => \N__34475\,
            I => \N__34471\
        );

    \I__7280\ : CascadeMux
    port map (
            O => \N__34474\,
            I => \N__34467\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__34471\,
            I => \N__34464\
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__34470\,
            I => \N__34461\
        );

    \I__7277\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34458\
        );

    \I__7276\ : Span4Mux_h
    port map (
            O => \N__34464\,
            I => \N__34455\
        );

    \I__7275\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34452\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__34458\,
            I => cmd_rdadctmp_23_adj_1053
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__34455\,
            I => cmd_rdadctmp_23_adj_1053
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__34452\,
            I => cmd_rdadctmp_23_adj_1053
        );

    \I__7271\ : InMux
    port map (
            O => \N__34445\,
            I => \N__34442\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__34442\,
            I => \N__34438\
        );

    \I__7269\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34435\
        );

    \I__7268\ : Span4Mux_v
    port map (
            O => \N__34438\,
            I => \N__34432\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__34435\,
            I => \N__34427\
        );

    \I__7266\ : Sp12to4
    port map (
            O => \N__34432\,
            I => \N__34427\
        );

    \I__7265\ : Odrv12
    port map (
            O => \N__34427\,
            I => buf_adcdata2_15
        );

    \I__7264\ : InMux
    port map (
            O => \N__34424\,
            I => \N__34420\
        );

    \I__7263\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34416\
        );

    \I__7262\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34413\
        );

    \I__7261\ : InMux
    port map (
            O => \N__34419\,
            I => \N__34410\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__34416\,
            I => \N__34400\
        );

    \I__7259\ : Span4Mux_v
    port map (
            O => \N__34413\,
            I => \N__34400\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__34410\,
            I => \N__34400\
        );

    \I__7257\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34397\
        );

    \I__7256\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34393\
        );

    \I__7255\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34390\
        );

    \I__7254\ : Span4Mux_v
    port map (
            O => \N__34400\,
            I => \N__34385\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__34397\,
            I => \N__34385\
        );

    \I__7252\ : InMux
    port map (
            O => \N__34396\,
            I => \N__34382\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__34393\,
            I => \N__34377\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__34390\,
            I => \N__34377\
        );

    \I__7249\ : Span4Mux_v
    port map (
            O => \N__34385\,
            I => \N__34374\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34370\
        );

    \I__7247\ : Span4Mux_v
    port map (
            O => \N__34377\,
            I => \N__34365\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__34374\,
            I => \N__34365\
        );

    \I__7245\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34362\
        );

    \I__7244\ : Span4Mux_h
    port map (
            O => \N__34370\,
            I => \N__34359\
        );

    \I__7243\ : Odrv4
    port map (
            O => \N__34365\,
            I => comm_buf_0_2
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__34362\,
            I => comm_buf_0_2
        );

    \I__7241\ : Odrv4
    port map (
            O => \N__34359\,
            I => comm_buf_0_2
        );

    \I__7240\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34349\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__34349\,
            I => \N__34345\
        );

    \I__7238\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34342\
        );

    \I__7237\ : Span4Mux_v
    port map (
            O => \N__34345\,
            I => \N__34338\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34335\
        );

    \I__7235\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34332\
        );

    \I__7234\ : Span4Mux_v
    port map (
            O => \N__34338\,
            I => \N__34327\
        );

    \I__7233\ : Span4Mux_v
    port map (
            O => \N__34335\,
            I => \N__34327\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__34332\,
            I => buf_dds_10
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__34327\,
            I => buf_dds_10
        );

    \I__7230\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34319\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__34319\,
            I => \N__34315\
        );

    \I__7228\ : InMux
    port map (
            O => \N__34318\,
            I => \N__34311\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__34315\,
            I => \N__34308\
        );

    \I__7226\ : InMux
    port map (
            O => \N__34314\,
            I => \N__34305\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__34311\,
            I => \acadc_skipCount_0\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__34308\,
            I => \acadc_skipCount_0\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__34305\,
            I => \acadc_skipCount_0\
        );

    \I__7222\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34295\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__34295\,
            I => n17_adj_1214
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__34292\,
            I => \N__34289\
        );

    \I__7219\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34286\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__34286\,
            I => \N__34281\
        );

    \I__7217\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34278\
        );

    \I__7216\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34275\
        );

    \I__7215\ : Odrv4
    port map (
            O => \N__34281\,
            I => req_data_cnt_0
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__34278\,
            I => req_data_cnt_0
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__34275\,
            I => req_data_cnt_0
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__34268\,
            I => \N__34265\
        );

    \I__7211\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34262\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__34262\,
            I => \N__34259\
        );

    \I__7209\ : Span12Mux_v
    port map (
            O => \N__34259\,
            I => \N__34256\
        );

    \I__7208\ : Odrv12
    port map (
            O => \N__34256\,
            I => buf_data1_21
        );

    \I__7207\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34250\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__34250\,
            I => \N__34247\
        );

    \I__7205\ : Span4Mux_v
    port map (
            O => \N__34247\,
            I => \N__34244\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__34244\,
            I => \N__34241\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__34241\,
            I => n66_adj_1158
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__34238\,
            I => \N__34235\
        );

    \I__7201\ : InMux
    port map (
            O => \N__34235\,
            I => \N__34230\
        );

    \I__7200\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34227\
        );

    \I__7199\ : InMux
    port map (
            O => \N__34233\,
            I => \N__34224\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__34230\,
            I => \N__34221\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__34227\,
            I => buf_dds_5
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__34224\,
            I => buf_dds_5
        );

    \I__7195\ : Odrv12
    port map (
            O => \N__34221\,
            I => buf_dds_5
        );

    \I__7194\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34211\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__34211\,
            I => \N__34207\
        );

    \I__7192\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34203\
        );

    \I__7191\ : Span4Mux_h
    port map (
            O => \N__34207\,
            I => \N__34200\
        );

    \I__7190\ : InMux
    port map (
            O => \N__34206\,
            I => \N__34197\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__34203\,
            I => \acadc_skipCount_10\
        );

    \I__7188\ : Odrv4
    port map (
            O => \N__34200\,
            I => \acadc_skipCount_10\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__34197\,
            I => \acadc_skipCount_10\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__34190\,
            I => \n7485_cascade_\
        );

    \I__7185\ : InMux
    port map (
            O => \N__34187\,
            I => \N__34181\
        );

    \I__7184\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34181\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__34181\,
            I => tacadc_rst
        );

    \I__7182\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34173\
        );

    \I__7181\ : InMux
    port map (
            O => \N__34177\,
            I => \N__34168\
        );

    \I__7180\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34168\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__34173\,
            I => req_data_cnt_10
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__34168\,
            I => req_data_cnt_10
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__34163\,
            I => \N__34160\
        );

    \I__7176\ : InMux
    port map (
            O => \N__34160\,
            I => \N__34157\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__34157\,
            I => n90_adj_1167
        );

    \I__7174\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34151\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__34151\,
            I => \N__34148\
        );

    \I__7172\ : Span4Mux_h
    port map (
            O => \N__34148\,
            I => \N__34145\
        );

    \I__7171\ : Odrv4
    port map (
            O => \N__34145\,
            I => n72_adj_1162
        );

    \I__7170\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34138\
        );

    \I__7169\ : CascadeMux
    port map (
            O => \N__34141\,
            I => \N__34135\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34130\
        );

    \I__7167\ : InMux
    port map (
            O => \N__34135\,
            I => \N__34125\
        );

    \I__7166\ : InMux
    port map (
            O => \N__34134\,
            I => \N__34125\
        );

    \I__7165\ : InMux
    port map (
            O => \N__34133\,
            I => \N__34121\
        );

    \I__7164\ : Span4Mux_h
    port map (
            O => \N__34130\,
            I => \N__34113\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__34125\,
            I => \N__34113\
        );

    \I__7162\ : InMux
    port map (
            O => \N__34124\,
            I => \N__34110\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__34121\,
            I => \N__34107\
        );

    \I__7160\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34102\
        );

    \I__7159\ : InMux
    port map (
            O => \N__34119\,
            I => \N__34102\
        );

    \I__7158\ : InMux
    port map (
            O => \N__34118\,
            I => \N__34099\
        );

    \I__7157\ : Span4Mux_v
    port map (
            O => \N__34113\,
            I => \N__34094\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__34110\,
            I => \N__34094\
        );

    \I__7155\ : Span4Mux_v
    port map (
            O => \N__34107\,
            I => \N__34089\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__34089\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__34099\,
            I => \N__34084\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__34094\,
            I => \N__34084\
        );

    \I__7151\ : Span4Mux_h
    port map (
            O => \N__34089\,
            I => \N__34081\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__34084\,
            I => \N__34078\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__34081\,
            I => \N__34075\
        );

    \I__7148\ : Odrv4
    port map (
            O => \N__34078\,
            I => comm_buf_0_0
        );

    \I__7147\ : Odrv4
    port map (
            O => \N__34075\,
            I => comm_buf_0_0
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__34070\,
            I => \n14_adj_1202_cascade_\
        );

    \I__7145\ : InMux
    port map (
            O => \N__34067\,
            I => \N__34064\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__34064\,
            I => \N__34061\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__34061\,
            I => \N__34056\
        );

    \I__7142\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34051\
        );

    \I__7141\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34051\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__34056\,
            I => buf_dds_13
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__34051\,
            I => buf_dds_13
        );

    \I__7138\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34043\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34040\
        );

    \I__7136\ : Odrv12
    port map (
            O => \N__34040\,
            I => n15690
        );

    \I__7135\ : InMux
    port map (
            O => \N__34037\,
            I => \N__34034\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__34034\,
            I => \N__34031\
        );

    \I__7133\ : Span4Mux_h
    port map (
            O => \N__34031\,
            I => \N__34026\
        );

    \I__7132\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34023\
        );

    \I__7131\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34020\
        );

    \I__7130\ : Span4Mux_h
    port map (
            O => \N__34026\,
            I => \N__34015\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__34015\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__34020\,
            I => req_data_cnt_12
        );

    \I__7127\ : Odrv4
    port map (
            O => \N__34015\,
            I => req_data_cnt_12
        );

    \I__7126\ : InMux
    port map (
            O => \N__34010\,
            I => \N__34007\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__34007\,
            I => \N__34004\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__34004\,
            I => n13_adj_1026
        );

    \I__7123\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33998\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__33998\,
            I => \N__33995\
        );

    \I__7121\ : Odrv12
    port map (
            O => \N__33995\,
            I => buf_data1_17
        );

    \I__7120\ : CascadeMux
    port map (
            O => \N__33992\,
            I => \n78_cascade_\
        );

    \I__7119\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33986\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__33986\,
            I => \N__33983\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__33983\,
            I => \N__33980\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__33980\,
            I => n99_adj_1024
        );

    \I__7115\ : InMux
    port map (
            O => \N__33977\,
            I => \N__33974\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__33974\,
            I => n4257
        );

    \I__7113\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33966\
        );

    \I__7112\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33963\
        );

    \I__7111\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33958\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__33966\,
            I => \N__33953\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__33963\,
            I => \N__33953\
        );

    \I__7108\ : InMux
    port map (
            O => \N__33962\,
            I => \N__33950\
        );

    \I__7107\ : InMux
    port map (
            O => \N__33961\,
            I => \N__33947\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__33958\,
            I => \N__33944\
        );

    \I__7105\ : Span4Mux_v
    port map (
            O => \N__33953\,
            I => \N__33941\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__33950\,
            I => \N__33938\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__33947\,
            I => \N__33933\
        );

    \I__7102\ : Span4Mux_h
    port map (
            O => \N__33944\,
            I => \N__33933\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__33941\,
            I => \N__33930\
        );

    \I__7100\ : Span12Mux_h
    port map (
            O => \N__33938\,
            I => \N__33927\
        );

    \I__7099\ : Sp12to4
    port map (
            O => \N__33933\,
            I => \N__33924\
        );

    \I__7098\ : Span4Mux_h
    port map (
            O => \N__33930\,
            I => \N__33921\
        );

    \I__7097\ : Odrv12
    port map (
            O => \N__33927\,
            I => comm_buf_1_6
        );

    \I__7096\ : Odrv12
    port map (
            O => \N__33924\,
            I => comm_buf_1_6
        );

    \I__7095\ : Odrv4
    port map (
            O => \N__33921\,
            I => comm_buf_1_6
        );

    \I__7094\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33911\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__33911\,
            I => n8133
        );

    \I__7092\ : CascadeMux
    port map (
            O => \N__33908\,
            I => \N__33904\
        );

    \I__7091\ : CascadeMux
    port map (
            O => \N__33907\,
            I => \N__33900\
        );

    \I__7090\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33897\
        );

    \I__7089\ : CascadeMux
    port map (
            O => \N__33903\,
            I => \N__33893\
        );

    \I__7088\ : InMux
    port map (
            O => \N__33900\,
            I => \N__33890\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__33897\,
            I => \N__33887\
        );

    \I__7086\ : InMux
    port map (
            O => \N__33896\,
            I => \N__33882\
        );

    \I__7085\ : InMux
    port map (
            O => \N__33893\,
            I => \N__33882\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__33890\,
            I => trig_dds
        );

    \I__7083\ : Odrv12
    port map (
            O => \N__33887\,
            I => trig_dds
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__33882\,
            I => trig_dds
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__33875\,
            I => \N__33872\
        );

    \I__7080\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33867\
        );

    \I__7079\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33864\
        );

    \I__7078\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33861\
        );

    \I__7077\ : LocalMux
    port map (
            O => \N__33867\,
            I => \N__33856\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__33864\,
            I => \N__33856\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__33861\,
            I => buf_dds_0
        );

    \I__7074\ : Odrv12
    port map (
            O => \N__33856\,
            I => buf_dds_0
        );

    \I__7073\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33846\
        );

    \I__7072\ : CascadeMux
    port map (
            O => \N__33850\,
            I => \N__33843\
        );

    \I__7071\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33840\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33837\
        );

    \I__7069\ : InMux
    port map (
            O => \N__33843\,
            I => \N__33834\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__33840\,
            I => \N__33831\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__33837\,
            I => \N__33828\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__33834\,
            I => buf_dds_8
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__33831\,
            I => buf_dds_8
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__33828\,
            I => buf_dds_8
        );

    \I__7063\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33818\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__33818\,
            I => \N__33815\
        );

    \I__7061\ : Span12Mux_v
    port map (
            O => \N__33815\,
            I => \N__33812\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__33812\,
            I => buf_data1_15
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__33809\,
            I => \n4190_cascade_\
        );

    \I__7058\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33803\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__33803\,
            I => n4227
        );

    \I__7056\ : InMux
    port map (
            O => \N__33800\,
            I => \N__33797\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__33797\,
            I => n4262
        );

    \I__7054\ : CascadeMux
    port map (
            O => \N__33794\,
            I => \N__33790\
        );

    \I__7053\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33786\
        );

    \I__7052\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33782\
        );

    \I__7051\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33779\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33776\
        );

    \I__7049\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33772\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__33782\,
            I => \N__33765\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__33779\,
            I => \N__33765\
        );

    \I__7046\ : Span4Mux_v
    port map (
            O => \N__33776\,
            I => \N__33765\
        );

    \I__7045\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33762\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__33772\,
            I => \N__33759\
        );

    \I__7043\ : Span4Mux_v
    port map (
            O => \N__33765\,
            I => \N__33756\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33753\
        );

    \I__7041\ : Span4Mux_v
    port map (
            O => \N__33759\,
            I => \N__33749\
        );

    \I__7040\ : Span4Mux_h
    port map (
            O => \N__33756\,
            I => \N__33744\
        );

    \I__7039\ : Span4Mux_h
    port map (
            O => \N__33753\,
            I => \N__33744\
        );

    \I__7038\ : InMux
    port map (
            O => \N__33752\,
            I => \N__33741\
        );

    \I__7037\ : Span4Mux_v
    port map (
            O => \N__33749\,
            I => \N__33736\
        );

    \I__7036\ : Span4Mux_h
    port map (
            O => \N__33744\,
            I => \N__33736\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__33741\,
            I => comm_buf_0_5
        );

    \I__7034\ : Odrv4
    port map (
            O => \N__33736\,
            I => comm_buf_0_5
        );

    \I__7033\ : CascadeMux
    port map (
            O => \N__33731\,
            I => \n13_cascade_\
        );

    \I__7032\ : InMux
    port map (
            O => \N__33728\,
            I => \N__33725\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__33725\,
            I => n6_adj_1273
        );

    \I__7030\ : InMux
    port map (
            O => \N__33722\,
            I => \N__33719\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__33719\,
            I => n5_adj_1282
        );

    \I__7028\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33712\
        );

    \I__7027\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33709\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__33712\,
            I => comm_length_0
        );

    \I__7025\ : LocalMux
    port map (
            O => \N__33709\,
            I => comm_length_0
        );

    \I__7024\ : SRMux
    port map (
            O => \N__33704\,
            I => \N__33701\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__33701\,
            I => \N__33697\
        );

    \I__7022\ : SRMux
    port map (
            O => \N__33700\,
            I => \N__33694\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__33697\,
            I => \N__33689\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33686\
        );

    \I__7019\ : SRMux
    port map (
            O => \N__33693\,
            I => \N__33683\
        );

    \I__7018\ : SRMux
    port map (
            O => \N__33692\,
            I => \N__33680\
        );

    \I__7017\ : Span4Mux_h
    port map (
            O => \N__33689\,
            I => \N__33677\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__33686\,
            I => \N__33674\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__33683\,
            I => \N__33669\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__33680\,
            I => \N__33669\
        );

    \I__7013\ : Span4Mux_h
    port map (
            O => \N__33677\,
            I => \N__33666\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__33674\,
            I => \N__33661\
        );

    \I__7011\ : Span4Mux_v
    port map (
            O => \N__33669\,
            I => \N__33661\
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__33666\,
            I => n10566
        );

    \I__7009\ : Odrv4
    port map (
            O => \N__33661\,
            I => n10566
        );

    \I__7008\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33653\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__33653\,
            I => n13
        );

    \I__7006\ : CascadeMux
    port map (
            O => \N__33650\,
            I => \N__33646\
        );

    \I__7005\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33641\
        );

    \I__7004\ : InMux
    port map (
            O => \N__33646\,
            I => \N__33641\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__33641\,
            I => \N__33638\
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__33638\,
            I => n12649
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__33635\,
            I => \n8525_cascade_\
        );

    \I__7000\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33629\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__33629\,
            I => \N__33622\
        );

    \I__6998\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33617\
        );

    \I__6997\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33617\
        );

    \I__6996\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33614\
        );

    \I__6995\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33611\
        );

    \I__6994\ : Span4Mux_v
    port map (
            O => \N__33622\,
            I => \N__33608\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__33617\,
            I => \N__33603\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__33614\,
            I => \N__33603\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__33611\,
            I => n4075
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__33608\,
            I => n4075
        );

    \I__6989\ : Odrv12
    port map (
            O => \N__33603\,
            I => n4075
        );

    \I__6988\ : CascadeMux
    port map (
            O => \N__33596\,
            I => \n15460_cascade_\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__33593\,
            I => \n19_cascade_\
        );

    \I__6986\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33587\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__33587\,
            I => n15463
        );

    \I__6984\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33581\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__33581\,
            I => \N__33578\
        );

    \I__6982\ : Span4Mux_v
    port map (
            O => \N__33578\,
            I => \N__33575\
        );

    \I__6981\ : Span4Mux_h
    port map (
            O => \N__33575\,
            I => \N__33572\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__33572\,
            I => n23
        );

    \I__6979\ : CascadeMux
    port map (
            O => \N__33569\,
            I => \n19_adj_1151_cascade_\
        );

    \I__6978\ : InMux
    port map (
            O => \N__33566\,
            I => \N__33563\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__33563\,
            I => \N__33560\
        );

    \I__6976\ : Span4Mux_v
    port map (
            O => \N__33560\,
            I => \N__33556\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__33559\,
            I => \N__33552\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__33556\,
            I => \N__33548\
        );

    \I__6973\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33541\
        );

    \I__6972\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33541\
        );

    \I__6971\ : InMux
    port map (
            O => \N__33551\,
            I => \N__33541\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__33548\,
            I => comm_length_2
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__33541\,
            I => comm_length_2
        );

    \I__6968\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33526\
        );

    \I__6967\ : InMux
    port map (
            O => \N__33535\,
            I => \N__33526\
        );

    \I__6966\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33513\
        );

    \I__6965\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33513\
        );

    \I__6964\ : InMux
    port map (
            O => \N__33532\,
            I => \N__33513\
        );

    \I__6963\ : InMux
    port map (
            O => \N__33531\,
            I => \N__33510\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__33526\,
            I => \N__33507\
        );

    \I__6961\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33502\
        );

    \I__6960\ : InMux
    port map (
            O => \N__33524\,
            I => \N__33502\
        );

    \I__6959\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33495\
        );

    \I__6958\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33495\
        );

    \I__6957\ : InMux
    port map (
            O => \N__33521\,
            I => \N__33495\
        );

    \I__6956\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33492\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__33513\,
            I => \N__33480\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__33510\,
            I => \N__33471\
        );

    \I__6953\ : Span4Mux_h
    port map (
            O => \N__33507\,
            I => \N__33471\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33471\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33471\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__33492\,
            I => \N__33468\
        );

    \I__6949\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33461\
        );

    \I__6948\ : InMux
    port map (
            O => \N__33490\,
            I => \N__33461\
        );

    \I__6947\ : InMux
    port map (
            O => \N__33489\,
            I => \N__33461\
        );

    \I__6946\ : CascadeMux
    port map (
            O => \N__33488\,
            I => \N__33456\
        );

    \I__6945\ : InMux
    port map (
            O => \N__33487\,
            I => \N__33453\
        );

    \I__6944\ : InMux
    port map (
            O => \N__33486\,
            I => \N__33450\
        );

    \I__6943\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33441\
        );

    \I__6942\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33441\
        );

    \I__6941\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33441\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__33480\,
            I => \N__33436\
        );

    \I__6939\ : Span4Mux_v
    port map (
            O => \N__33471\,
            I => \N__33436\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__33468\,
            I => \N__33431\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__33461\,
            I => \N__33431\
        );

    \I__6936\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33424\
        );

    \I__6935\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33424\
        );

    \I__6934\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33424\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33419\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__33450\,
            I => \N__33419\
        );

    \I__6931\ : CascadeMux
    port map (
            O => \N__33449\,
            I => \N__33416\
        );

    \I__6930\ : InMux
    port map (
            O => \N__33448\,
            I => \N__33411\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__33441\,
            I => \N__33408\
        );

    \I__6928\ : Span4Mux_h
    port map (
            O => \N__33436\,
            I => \N__33405\
        );

    \I__6927\ : Span4Mux_h
    port map (
            O => \N__33431\,
            I => \N__33400\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__33424\,
            I => \N__33400\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__33419\,
            I => \N__33397\
        );

    \I__6924\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33394\
        );

    \I__6923\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33389\
        );

    \I__6922\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33389\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__33411\,
            I => comm_index_2
        );

    \I__6920\ : Odrv12
    port map (
            O => \N__33408\,
            I => comm_index_2
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__33405\,
            I => comm_index_2
        );

    \I__6918\ : Odrv4
    port map (
            O => \N__33400\,
            I => comm_index_2
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__33397\,
            I => comm_index_2
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__33394\,
            I => comm_index_2
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__33389\,
            I => comm_index_2
        );

    \I__6914\ : CascadeMux
    port map (
            O => \N__33374\,
            I => \N__33368\
        );

    \I__6913\ : InMux
    port map (
            O => \N__33373\,
            I => \N__33363\
        );

    \I__6912\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33363\
        );

    \I__6911\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33358\
        );

    \I__6910\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33358\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__33363\,
            I => comm_length_3
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__33358\,
            I => comm_length_3
        );

    \I__6907\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33343\
        );

    \I__6906\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33340\
        );

    \I__6905\ : InMux
    port map (
            O => \N__33351\,
            I => \N__33337\
        );

    \I__6904\ : InMux
    port map (
            O => \N__33350\,
            I => \N__33332\
        );

    \I__6903\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33332\
        );

    \I__6902\ : InMux
    port map (
            O => \N__33348\,
            I => \N__33325\
        );

    \I__6901\ : InMux
    port map (
            O => \N__33347\,
            I => \N__33322\
        );

    \I__6900\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33317\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__33343\,
            I => \N__33312\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__33340\,
            I => \N__33312\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__33337\,
            I => \N__33307\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33307\
        );

    \I__6895\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33302\
        );

    \I__6894\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33302\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__33329\,
            I => \N__33299\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__33328\,
            I => \N__33296\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__33325\,
            I => \N__33291\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__33322\,
            I => \N__33288\
        );

    \I__6889\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33285\
        );

    \I__6888\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33282\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__33317\,
            I => \N__33279\
        );

    \I__6886\ : Span4Mux_h
    port map (
            O => \N__33312\,
            I => \N__33272\
        );

    \I__6885\ : Span4Mux_v
    port map (
            O => \N__33307\,
            I => \N__33272\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__33302\,
            I => \N__33272\
        );

    \I__6883\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33269\
        );

    \I__6882\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33262\
        );

    \I__6881\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33262\
        );

    \I__6880\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33262\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__33291\,
            I => \N__33255\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__33288\,
            I => \N__33255\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__33285\,
            I => \N__33255\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33252\
        );

    \I__6875\ : Span4Mux_v
    port map (
            O => \N__33279\,
            I => \N__33246\
        );

    \I__6874\ : Span4Mux_h
    port map (
            O => \N__33272\,
            I => \N__33239\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__33269\,
            I => \N__33239\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__33262\,
            I => \N__33239\
        );

    \I__6871\ : Span4Mux_h
    port map (
            O => \N__33255\,
            I => \N__33234\
        );

    \I__6870\ : Span4Mux_v
    port map (
            O => \N__33252\,
            I => \N__33234\
        );

    \I__6869\ : InMux
    port map (
            O => \N__33251\,
            I => \N__33229\
        );

    \I__6868\ : InMux
    port map (
            O => \N__33250\,
            I => \N__33229\
        );

    \I__6867\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33226\
        );

    \I__6866\ : Odrv4
    port map (
            O => \N__33246\,
            I => comm_index_3
        );

    \I__6865\ : Odrv4
    port map (
            O => \N__33239\,
            I => comm_index_3
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__33234\,
            I => comm_index_3
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__33229\,
            I => comm_index_3
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__33226\,
            I => comm_index_3
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__33215\,
            I => \n6_adj_1281_cascade_\
        );

    \I__6860\ : InMux
    port map (
            O => \N__33212\,
            I => \N__33202\
        );

    \I__6859\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33195\
        );

    \I__6858\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33195\
        );

    \I__6857\ : InMux
    port map (
            O => \N__33209\,
            I => \N__33195\
        );

    \I__6856\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33188\
        );

    \I__6855\ : InMux
    port map (
            O => \N__33207\,
            I => \N__33188\
        );

    \I__6854\ : InMux
    port map (
            O => \N__33206\,
            I => \N__33188\
        );

    \I__6853\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33185\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__33202\,
            I => \N__33163\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33163\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__33188\,
            I => \N__33160\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__33185\,
            I => \N__33157\
        );

    \I__6848\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33146\
        );

    \I__6847\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33146\
        );

    \I__6846\ : InMux
    port map (
            O => \N__33182\,
            I => \N__33146\
        );

    \I__6845\ : InMux
    port map (
            O => \N__33181\,
            I => \N__33146\
        );

    \I__6844\ : InMux
    port map (
            O => \N__33180\,
            I => \N__33146\
        );

    \I__6843\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33141\
        );

    \I__6842\ : InMux
    port map (
            O => \N__33178\,
            I => \N__33141\
        );

    \I__6841\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33138\
        );

    \I__6840\ : InMux
    port map (
            O => \N__33176\,
            I => \N__33133\
        );

    \I__6839\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33133\
        );

    \I__6838\ : InMux
    port map (
            O => \N__33174\,
            I => \N__33121\
        );

    \I__6837\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33121\
        );

    \I__6836\ : InMux
    port map (
            O => \N__33172\,
            I => \N__33121\
        );

    \I__6835\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33121\
        );

    \I__6834\ : InMux
    port map (
            O => \N__33170\,
            I => \N__33118\
        );

    \I__6833\ : CascadeMux
    port map (
            O => \N__33169\,
            I => \N__33113\
        );

    \I__6832\ : CascadeMux
    port map (
            O => \N__33168\,
            I => \N__33107\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__33163\,
            I => \N__33091\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__33160\,
            I => \N__33091\
        );

    \I__6829\ : Span4Mux_v
    port map (
            O => \N__33157\,
            I => \N__33086\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__33146\,
            I => \N__33086\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__33141\,
            I => \N__33080\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__33138\,
            I => \N__33080\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__33133\,
            I => \N__33077\
        );

    \I__6824\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33070\
        );

    \I__6823\ : InMux
    port map (
            O => \N__33131\,
            I => \N__33070\
        );

    \I__6822\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33070\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__33121\,
            I => \N__33065\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__33118\,
            I => \N__33065\
        );

    \I__6819\ : InMux
    port map (
            O => \N__33117\,
            I => \N__33062\
        );

    \I__6818\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33059\
        );

    \I__6817\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33052\
        );

    \I__6816\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33052\
        );

    \I__6815\ : InMux
    port map (
            O => \N__33111\,
            I => \N__33052\
        );

    \I__6814\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33041\
        );

    \I__6813\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33041\
        );

    \I__6812\ : InMux
    port map (
            O => \N__33106\,
            I => \N__33041\
        );

    \I__6811\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33041\
        );

    \I__6810\ : InMux
    port map (
            O => \N__33104\,
            I => \N__33041\
        );

    \I__6809\ : InMux
    port map (
            O => \N__33103\,
            I => \N__33038\
        );

    \I__6808\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33031\
        );

    \I__6807\ : InMux
    port map (
            O => \N__33101\,
            I => \N__33031\
        );

    \I__6806\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33031\
        );

    \I__6805\ : InMux
    port map (
            O => \N__33099\,
            I => \N__33028\
        );

    \I__6804\ : InMux
    port map (
            O => \N__33098\,
            I => \N__33021\
        );

    \I__6803\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33021\
        );

    \I__6802\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33021\
        );

    \I__6801\ : Span4Mux_h
    port map (
            O => \N__33091\,
            I => \N__33015\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__33086\,
            I => \N__33015\
        );

    \I__6799\ : InMux
    port map (
            O => \N__33085\,
            I => \N__33012\
        );

    \I__6798\ : Span4Mux_v
    port map (
            O => \N__33080\,
            I => \N__33007\
        );

    \I__6797\ : Span4Mux_v
    port map (
            O => \N__33077\,
            I => \N__33007\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33002\
        );

    \I__6795\ : Span4Mux_v
    port map (
            O => \N__33065\,
            I => \N__33002\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__32997\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__33059\,
            I => \N__32997\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__33052\,
            I => \N__32994\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__33041\,
            I => \N__32991\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__33038\,
            I => \N__32982\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__33031\,
            I => \N__32982\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__32982\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__33021\,
            I => \N__32982\
        );

    \I__6786\ : InMux
    port map (
            O => \N__33020\,
            I => \N__32979\
        );

    \I__6785\ : Span4Mux_h
    port map (
            O => \N__33015\,
            I => \N__32976\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__32973\
        );

    \I__6783\ : Span4Mux_h
    port map (
            O => \N__33007\,
            I => \N__32964\
        );

    \I__6782\ : Span4Mux_h
    port map (
            O => \N__33002\,
            I => \N__32964\
        );

    \I__6781\ : Span4Mux_v
    port map (
            O => \N__32997\,
            I => \N__32964\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__32994\,
            I => \N__32964\
        );

    \I__6779\ : Span12Mux_h
    port map (
            O => \N__32991\,
            I => \N__32959\
        );

    \I__6778\ : Span12Mux_v
    port map (
            O => \N__32982\,
            I => \N__32959\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__32979\,
            I => comm_index_1
        );

    \I__6776\ : Odrv4
    port map (
            O => \N__32976\,
            I => comm_index_1
        );

    \I__6775\ : Odrv4
    port map (
            O => \N__32973\,
            I => comm_index_1
        );

    \I__6774\ : Odrv4
    port map (
            O => \N__32964\,
            I => comm_index_1
        );

    \I__6773\ : Odrv12
    port map (
            O => \N__32959\,
            I => comm_index_1
        );

    \I__6772\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32945\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__32945\,
            I => n2
        );

    \I__6770\ : CascadeMux
    port map (
            O => \N__32942\,
            I => \n15119_cascade_\
        );

    \I__6769\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32933\
        );

    \I__6768\ : InMux
    port map (
            O => \N__32938\,
            I => \N__32933\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__32933\,
            I => comm_length_1
        );

    \I__6766\ : InMux
    port map (
            O => \N__32930\,
            I => \N__32927\
        );

    \I__6765\ : LocalMux
    port map (
            O => \N__32927\,
            I => \N__32920\
        );

    \I__6764\ : InMux
    port map (
            O => \N__32926\,
            I => \N__32917\
        );

    \I__6763\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32913\
        );

    \I__6762\ : CascadeMux
    port map (
            O => \N__32924\,
            I => \N__32908\
        );

    \I__6761\ : CascadeMux
    port map (
            O => \N__32923\,
            I => \N__32905\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__32920\,
            I => \N__32900\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__32917\,
            I => \N__32900\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__32916\,
            I => \N__32896\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__32913\,
            I => \N__32893\
        );

    \I__6756\ : CascadeMux
    port map (
            O => \N__32912\,
            I => \N__32890\
        );

    \I__6755\ : InMux
    port map (
            O => \N__32911\,
            I => \N__32882\
        );

    \I__6754\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32882\
        );

    \I__6753\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32882\
        );

    \I__6752\ : Span4Mux_h
    port map (
            O => \N__32900\,
            I => \N__32879\
        );

    \I__6751\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32872\
        );

    \I__6750\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32872\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__32893\,
            I => \N__32869\
        );

    \I__6748\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32866\
        );

    \I__6747\ : InMux
    port map (
            O => \N__32889\,
            I => \N__32863\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__32882\,
            I => \N__32858\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__32879\,
            I => \N__32858\
        );

    \I__6744\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32853\
        );

    \I__6743\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32853\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__32872\,
            I => eis_state_0
        );

    \I__6741\ : Odrv4
    port map (
            O => \N__32869\,
            I => eis_state_0
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__32866\,
            I => eis_state_0
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__32863\,
            I => eis_state_0
        );

    \I__6738\ : Odrv4
    port map (
            O => \N__32858\,
            I => eis_state_0
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__32853\,
            I => eis_state_0
        );

    \I__6736\ : CascadeMux
    port map (
            O => \N__32840\,
            I => \N__32837\
        );

    \I__6735\ : InMux
    port map (
            O => \N__32837\,
            I => \N__32826\
        );

    \I__6734\ : InMux
    port map (
            O => \N__32836\,
            I => \N__32826\
        );

    \I__6733\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32826\
        );

    \I__6732\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32823\
        );

    \I__6731\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32820\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__32826\,
            I => \N__32815\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__32823\,
            I => \N__32815\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__32820\,
            I => \N__32803\
        );

    \I__6727\ : Span4Mux_v
    port map (
            O => \N__32815\,
            I => \N__32803\
        );

    \I__6726\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32798\
        );

    \I__6725\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32798\
        );

    \I__6724\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32795\
        );

    \I__6723\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32790\
        );

    \I__6722\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32790\
        );

    \I__6721\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32785\
        );

    \I__6720\ : InMux
    port map (
            O => \N__32808\,
            I => \N__32785\
        );

    \I__6719\ : Span4Mux_v
    port map (
            O => \N__32803\,
            I => \N__32782\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__32798\,
            I => \eis_end_N_770\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__32795\,
            I => \eis_end_N_770\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__32790\,
            I => \eis_end_N_770\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__32785\,
            I => \eis_end_N_770\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__32782\,
            I => \eis_end_N_770\
        );

    \I__6713\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32768\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__32768\,
            I => \N__32764\
        );

    \I__6711\ : CascadeMux
    port map (
            O => \N__32767\,
            I => \N__32760\
        );

    \I__6710\ : Span4Mux_v
    port map (
            O => \N__32764\,
            I => \N__32757\
        );

    \I__6709\ : CascadeMux
    port map (
            O => \N__32763\,
            I => \N__32754\
        );

    \I__6708\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32750\
        );

    \I__6707\ : Span4Mux_h
    port map (
            O => \N__32757\,
            I => \N__32747\
        );

    \I__6706\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32744\
        );

    \I__6705\ : SRMux
    port map (
            O => \N__32753\,
            I => \N__32741\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__32750\,
            I => \N__32738\
        );

    \I__6703\ : Span4Mux_h
    port map (
            O => \N__32747\,
            I => \N__32730\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__32744\,
            I => \N__32730\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32725\
        );

    \I__6700\ : Span4Mux_h
    port map (
            O => \N__32738\,
            I => \N__32722\
        );

    \I__6699\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32715\
        );

    \I__6698\ : InMux
    port map (
            O => \N__32736\,
            I => \N__32715\
        );

    \I__6697\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32715\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__32730\,
            I => \N__32712\
        );

    \I__6695\ : InMux
    port map (
            O => \N__32729\,
            I => \N__32707\
        );

    \I__6694\ : InMux
    port map (
            O => \N__32728\,
            I => \N__32707\
        );

    \I__6693\ : Span4Mux_v
    port map (
            O => \N__32725\,
            I => \N__32704\
        );

    \I__6692\ : Span4Mux_v
    port map (
            O => \N__32722\,
            I => \N__32699\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32699\
        );

    \I__6690\ : Sp12to4
    port map (
            O => \N__32712\,
            I => \N__32696\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__32707\,
            I => \N__32693\
        );

    \I__6688\ : Span4Mux_v
    port map (
            O => \N__32704\,
            I => \N__32688\
        );

    \I__6687\ : Span4Mux_v
    port map (
            O => \N__32699\,
            I => \N__32688\
        );

    \I__6686\ : Span12Mux_h
    port map (
            O => \N__32696\,
            I => \N__32685\
        );

    \I__6685\ : Span12Mux_v
    port map (
            O => \N__32693\,
            I => \N__32682\
        );

    \I__6684\ : Sp12to4
    port map (
            O => \N__32688\,
            I => \N__32679\
        );

    \I__6683\ : Span12Mux_v
    port map (
            O => \N__32685\,
            I => \N__32676\
        );

    \I__6682\ : Span12Mux_v
    port map (
            O => \N__32682\,
            I => \N__32673\
        );

    \I__6681\ : Span12Mux_h
    port map (
            O => \N__32679\,
            I => \N__32670\
        );

    \I__6680\ : Span12Mux_v
    port map (
            O => \N__32676\,
            I => \N__32667\
        );

    \I__6679\ : Span12Mux_h
    port map (
            O => \N__32673\,
            I => \N__32662\
        );

    \I__6678\ : Span12Mux_v
    port map (
            O => \N__32670\,
            I => \N__32662\
        );

    \I__6677\ : Odrv12
    port map (
            O => \N__32667\,
            I => \ICE_GPMO_0\
        );

    \I__6676\ : Odrv12
    port map (
            O => \N__32662\,
            I => \ICE_GPMO_0\
        );

    \I__6675\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32652\
        );

    \I__6674\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32647\
        );

    \I__6673\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32647\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__32652\,
            I => \N__32644\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__32647\,
            I => \N__32641\
        );

    \I__6670\ : Span4Mux_h
    port map (
            O => \N__32644\,
            I => \N__32636\
        );

    \I__6669\ : Span4Mux_h
    port map (
            O => \N__32641\,
            I => \N__32636\
        );

    \I__6668\ : Odrv4
    port map (
            O => \N__32636\,
            I => data_index_8
        );

    \I__6667\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32630\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__32630\,
            I => \N__32627\
        );

    \I__6665\ : Odrv12
    port map (
            O => \N__32627\,
            I => buf_data1_3
        );

    \I__6664\ : InMux
    port map (
            O => \N__32624\,
            I => \N__32620\
        );

    \I__6663\ : InMux
    port map (
            O => \N__32623\,
            I => \N__32616\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__32620\,
            I => \N__32613\
        );

    \I__6661\ : CascadeMux
    port map (
            O => \N__32619\,
            I => \N__32610\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__32616\,
            I => \N__32607\
        );

    \I__6659\ : Span12Mux_v
    port map (
            O => \N__32613\,
            I => \N__32604\
        );

    \I__6658\ : InMux
    port map (
            O => \N__32610\,
            I => \N__32601\
        );

    \I__6657\ : Sp12to4
    port map (
            O => \N__32607\,
            I => \N__32598\
        );

    \I__6656\ : Span12Mux_h
    port map (
            O => \N__32604\,
            I => \N__32595\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__32601\,
            I => \N__32590\
        );

    \I__6654\ : Span12Mux_v
    port map (
            O => \N__32598\,
            I => \N__32590\
        );

    \I__6653\ : Span12Mux_v
    port map (
            O => \N__32595\,
            I => \N__32587\
        );

    \I__6652\ : Odrv12
    port map (
            O => \N__32590\,
            I => buf_adcdata3_3
        );

    \I__6651\ : Odrv12
    port map (
            O => \N__32587\,
            I => buf_adcdata3_3
        );

    \I__6650\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32579\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__32579\,
            I => \N__32576\
        );

    \I__6648\ : Span4Mux_v
    port map (
            O => \N__32576\,
            I => \N__32573\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__32573\,
            I => \N__32570\
        );

    \I__6646\ : Span4Mux_h
    port map (
            O => \N__32570\,
            I => \N__32567\
        );

    \I__6645\ : Odrv4
    port map (
            O => \N__32567\,
            I => n4149
        );

    \I__6644\ : InMux
    port map (
            O => \N__32564\,
            I => \N__32559\
        );

    \I__6643\ : InMux
    port map (
            O => \N__32563\,
            I => \N__32554\
        );

    \I__6642\ : InMux
    port map (
            O => \N__32562\,
            I => \N__32554\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__32559\,
            I => \N__32551\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__32554\,
            I => \N__32548\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__32551\,
            I => \N__32543\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__32548\,
            I => \N__32543\
        );

    \I__6637\ : Span4Mux_h
    port map (
            O => \N__32543\,
            I => \N__32540\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__32540\,
            I => comm_tx_buf_5
        );

    \I__6635\ : SRMux
    port map (
            O => \N__32537\,
            I => \N__32534\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__32534\,
            I => \N__32531\
        );

    \I__6633\ : Span4Mux_v
    port map (
            O => \N__32531\,
            I => \N__32528\
        );

    \I__6632\ : Sp12to4
    port map (
            O => \N__32528\,
            I => \N__32525\
        );

    \I__6631\ : Odrv12
    port map (
            O => \N__32525\,
            I => \comm_spi.data_tx_7__N_819\
        );

    \I__6630\ : CEMux
    port map (
            O => \N__32522\,
            I => \N__32519\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__32519\,
            I => \N__32515\
        );

    \I__6628\ : CEMux
    port map (
            O => \N__32518\,
            I => \N__32512\
        );

    \I__6627\ : Span4Mux_h
    port map (
            O => \N__32515\,
            I => \N__32509\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32506\
        );

    \I__6625\ : Odrv4
    port map (
            O => \N__32509\,
            I => n8561
        );

    \I__6624\ : Odrv4
    port map (
            O => \N__32506\,
            I => n8561
        );

    \I__6623\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32497\
        );

    \I__6622\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32494\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__32497\,
            I => n8_adj_1229
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__32494\,
            I => n8_adj_1229
        );

    \I__6619\ : InMux
    port map (
            O => \N__32489\,
            I => \N__32485\
        );

    \I__6618\ : InMux
    port map (
            O => \N__32488\,
            I => \N__32482\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__32485\,
            I => n7_adj_1228
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__32482\,
            I => n7_adj_1228
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__32477\,
            I => \N__32474\
        );

    \I__6614\ : CascadeBuf
    port map (
            O => \N__32474\,
            I => \N__32471\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__32471\,
            I => \N__32468\
        );

    \I__6612\ : CascadeBuf
    port map (
            O => \N__32468\,
            I => \N__32465\
        );

    \I__6611\ : CascadeMux
    port map (
            O => \N__32465\,
            I => \N__32462\
        );

    \I__6610\ : CascadeBuf
    port map (
            O => \N__32462\,
            I => \N__32459\
        );

    \I__6609\ : CascadeMux
    port map (
            O => \N__32459\,
            I => \N__32456\
        );

    \I__6608\ : CascadeBuf
    port map (
            O => \N__32456\,
            I => \N__32453\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__32453\,
            I => \N__32450\
        );

    \I__6606\ : CascadeBuf
    port map (
            O => \N__32450\,
            I => \N__32447\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__32447\,
            I => \N__32444\
        );

    \I__6604\ : CascadeBuf
    port map (
            O => \N__32444\,
            I => \N__32441\
        );

    \I__6603\ : CascadeMux
    port map (
            O => \N__32441\,
            I => \N__32437\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__32440\,
            I => \N__32434\
        );

    \I__6601\ : CascadeBuf
    port map (
            O => \N__32437\,
            I => \N__32431\
        );

    \I__6600\ : CascadeBuf
    port map (
            O => \N__32434\,
            I => \N__32428\
        );

    \I__6599\ : CascadeMux
    port map (
            O => \N__32431\,
            I => \N__32425\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__32428\,
            I => \N__32422\
        );

    \I__6597\ : CascadeBuf
    port map (
            O => \N__32425\,
            I => \N__32419\
        );

    \I__6596\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32416\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__32419\,
            I => \N__32413\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32410\
        );

    \I__6593\ : CascadeBuf
    port map (
            O => \N__32413\,
            I => \N__32407\
        );

    \I__6592\ : Span4Mux_h
    port map (
            O => \N__32410\,
            I => \N__32404\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__32407\,
            I => \N__32401\
        );

    \I__6590\ : Span4Mux_v
    port map (
            O => \N__32404\,
            I => \N__32398\
        );

    \I__6589\ : InMux
    port map (
            O => \N__32401\,
            I => \N__32395\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__32398\,
            I => \N__32392\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__32395\,
            I => \N__32389\
        );

    \I__6586\ : Span4Mux_h
    port map (
            O => \N__32392\,
            I => \N__32386\
        );

    \I__6585\ : Span4Mux_h
    port map (
            O => \N__32389\,
            I => \N__32383\
        );

    \I__6584\ : Span4Mux_h
    port map (
            O => \N__32386\,
            I => \N__32378\
        );

    \I__6583\ : Span4Mux_h
    port map (
            O => \N__32383\,
            I => \N__32378\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__32378\,
            I => \data_index_9_N_258_3\
        );

    \I__6581\ : CEMux
    port map (
            O => \N__32375\,
            I => \N__32372\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__32372\,
            I => \N__32368\
        );

    \I__6579\ : CEMux
    port map (
            O => \N__32371\,
            I => \N__32364\
        );

    \I__6578\ : Span4Mux_h
    port map (
            O => \N__32368\,
            I => \N__32361\
        );

    \I__6577\ : CEMux
    port map (
            O => \N__32367\,
            I => \N__32358\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32355\
        );

    \I__6575\ : Span4Mux_h
    port map (
            O => \N__32361\,
            I => \N__32352\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__32358\,
            I => \N__32349\
        );

    \I__6573\ : Span4Mux_h
    port map (
            O => \N__32355\,
            I => \N__32346\
        );

    \I__6572\ : Span4Mux_h
    port map (
            O => \N__32352\,
            I => \N__32342\
        );

    \I__6571\ : Span4Mux_h
    port map (
            O => \N__32349\,
            I => \N__32339\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__32346\,
            I => \N__32336\
        );

    \I__6569\ : InMux
    port map (
            O => \N__32345\,
            I => \N__32333\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__32342\,
            I => n8456
        );

    \I__6567\ : Odrv4
    port map (
            O => \N__32339\,
            I => n8456
        );

    \I__6566\ : Odrv4
    port map (
            O => \N__32336\,
            I => n8456
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__32333\,
            I => n8456
        );

    \I__6564\ : InMux
    port map (
            O => \N__32324\,
            I => \N__32320\
        );

    \I__6563\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32317\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__32320\,
            I => \N__32312\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__32317\,
            I => \N__32312\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__32312\,
            I => acadc_skipcnt_3
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__32309\,
            I => \N__32306\
        );

    \I__6558\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32302\
        );

    \I__6557\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32299\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__32302\,
            I => \N__32296\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__32299\,
            I => acadc_skipcnt_5
        );

    \I__6554\ : Odrv4
    port map (
            O => \N__32296\,
            I => acadc_skipcnt_5
        );

    \I__6553\ : InMux
    port map (
            O => \N__32291\,
            I => \N__32287\
        );

    \I__6552\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32284\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__32287\,
            I => \N__32281\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__32284\,
            I => acadc_skipcnt_8
        );

    \I__6549\ : Odrv4
    port map (
            O => \N__32281\,
            I => acadc_skipcnt_8
        );

    \I__6548\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32273\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__32273\,
            I => \N__32268\
        );

    \I__6546\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32265\
        );

    \I__6545\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32262\
        );

    \I__6544\ : Span4Mux_v
    port map (
            O => \N__32268\,
            I => \N__32259\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32256\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__32262\,
            I => \acadc_skipCount_8\
        );

    \I__6541\ : Odrv4
    port map (
            O => \N__32259\,
            I => \acadc_skipCount_8\
        );

    \I__6540\ : Odrv4
    port map (
            O => \N__32256\,
            I => \acadc_skipCount_8\
        );

    \I__6539\ : CascadeMux
    port map (
            O => \N__32249\,
            I => \n20_cascade_\
        );

    \I__6538\ : InMux
    port map (
            O => \N__32246\,
            I => \N__32243\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__32243\,
            I => \N__32240\
        );

    \I__6536\ : Span4Mux_h
    port map (
            O => \N__32240\,
            I => \N__32237\
        );

    \I__6535\ : Odrv4
    port map (
            O => \N__32237\,
            I => n26
        );

    \I__6534\ : InMux
    port map (
            O => \N__32234\,
            I => \N__32231\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__32231\,
            I => \N__32227\
        );

    \I__6532\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32224\
        );

    \I__6531\ : Span4Mux_h
    port map (
            O => \N__32227\,
            I => \N__32221\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__32224\,
            I => acadc_skipcnt_13
        );

    \I__6529\ : Odrv4
    port map (
            O => \N__32221\,
            I => acadc_skipcnt_13
        );

    \I__6528\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32212\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__32215\,
            I => \N__32209\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__32212\,
            I => \N__32206\
        );

    \I__6525\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32202\
        );

    \I__6524\ : Span12Mux_h
    port map (
            O => \N__32206\,
            I => \N__32199\
        );

    \I__6523\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32196\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__32202\,
            I => \acadc_skipCount_13\
        );

    \I__6521\ : Odrv12
    port map (
            O => \N__32199\,
            I => \acadc_skipCount_13\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__32196\,
            I => \acadc_skipCount_13\
        );

    \I__6519\ : InMux
    port map (
            O => \N__32189\,
            I => \N__32186\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__32186\,
            I => n14_adj_1160
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__32183\,
            I => \N__32180\
        );

    \I__6516\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32177\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__32177\,
            I => \N__32174\
        );

    \I__6514\ : Span4Mux_v
    port map (
            O => \N__32174\,
            I => \N__32170\
        );

    \I__6513\ : InMux
    port map (
            O => \N__32173\,
            I => \N__32167\
        );

    \I__6512\ : Span4Mux_h
    port map (
            O => \N__32170\,
            I => \N__32161\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__32167\,
            I => \N__32161\
        );

    \I__6510\ : CascadeMux
    port map (
            O => \N__32166\,
            I => \N__32158\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__32161\,
            I => \N__32155\
        );

    \I__6508\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32152\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__32155\,
            I => cmd_rdadctmp_16
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__32152\,
            I => cmd_rdadctmp_16
        );

    \I__6505\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32144\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__32144\,
            I => \N__32141\
        );

    \I__6503\ : Span4Mux_h
    port map (
            O => \N__32141\,
            I => \N__32137\
        );

    \I__6502\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32134\
        );

    \I__6501\ : Span4Mux_h
    port map (
            O => \N__32137\,
            I => \N__32131\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__32134\,
            I => buf_adcdata1_8
        );

    \I__6499\ : Odrv4
    port map (
            O => \N__32131\,
            I => buf_adcdata1_8
        );

    \I__6498\ : InMux
    port map (
            O => \N__32126\,
            I => \N__32122\
        );

    \I__6497\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32119\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__32122\,
            I => \N__32115\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__32119\,
            I => \N__32112\
        );

    \I__6494\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32109\
        );

    \I__6493\ : Span4Mux_v
    port map (
            O => \N__32115\,
            I => \N__32105\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__32112\,
            I => \N__32101\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__32109\,
            I => \N__32098\
        );

    \I__6490\ : InMux
    port map (
            O => \N__32108\,
            I => \N__32095\
        );

    \I__6489\ : Span4Mux_h
    port map (
            O => \N__32105\,
            I => \N__32091\
        );

    \I__6488\ : InMux
    port map (
            O => \N__32104\,
            I => \N__32088\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__32101\,
            I => \N__32081\
        );

    \I__6486\ : Span4Mux_v
    port map (
            O => \N__32098\,
            I => \N__32081\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__32095\,
            I => \N__32081\
        );

    \I__6484\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32078\
        );

    \I__6483\ : Odrv4
    port map (
            O => \N__32091\,
            I => n84
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__32088\,
            I => n84
        );

    \I__6481\ : Odrv4
    port map (
            O => \N__32081\,
            I => n84
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__32078\,
            I => n84
        );

    \I__6479\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32066\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__32063\
        );

    \I__6477\ : Span4Mux_h
    port map (
            O => \N__32063\,
            I => \N__32060\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__32060\,
            I => n15546
        );

    \I__6475\ : InMux
    port map (
            O => \N__32057\,
            I => \N__32052\
        );

    \I__6474\ : InMux
    port map (
            O => \N__32056\,
            I => \N__32049\
        );

    \I__6473\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32046\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__32052\,
            I => data_index_5
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__32049\,
            I => data_index_5
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__32046\,
            I => data_index_5
        );

    \I__6469\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32035\
        );

    \I__6468\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32032\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__32035\,
            I => \N__32026\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__32032\,
            I => \N__32026\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__32031\,
            I => \N__32023\
        );

    \I__6464\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__32020\
        );

    \I__6463\ : InMux
    port map (
            O => \N__32023\,
            I => \N__32017\
        );

    \I__6462\ : Span4Mux_v
    port map (
            O => \N__32020\,
            I => \N__32014\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__32017\,
            I => buf_dds_12
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__32014\,
            I => buf_dds_12
        );

    \I__6459\ : InMux
    port map (
            O => \N__32009\,
            I => \N__32006\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__32006\,
            I => \N__32002\
        );

    \I__6457\ : InMux
    port map (
            O => \N__32005\,
            I => \N__31999\
        );

    \I__6456\ : Span4Mux_v
    port map (
            O => \N__32002\,
            I => \N__31996\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__31999\,
            I => acadc_skipcnt_2
        );

    \I__6454\ : Odrv4
    port map (
            O => \N__31996\,
            I => acadc_skipcnt_2
        );

    \I__6453\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31988\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31983\
        );

    \I__6451\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31980\
        );

    \I__6450\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31977\
        );

    \I__6449\ : Sp12to4
    port map (
            O => \N__31983\,
            I => \N__31972\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__31980\,
            I => \N__31972\
        );

    \I__6447\ : LocalMux
    port map (
            O => \N__31977\,
            I => \acadc_skipCount_7\
        );

    \I__6446\ : Odrv12
    port map (
            O => \N__31972\,
            I => \acadc_skipCount_7\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__31967\,
            I => \N__31964\
        );

    \I__6444\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31961\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__31961\,
            I => \N__31957\
        );

    \I__6442\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31954\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__31957\,
            I => \N__31951\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__31954\,
            I => acadc_skipcnt_7
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__31951\,
            I => acadc_skipcnt_7
        );

    \I__6438\ : InMux
    port map (
            O => \N__31946\,
            I => \N__31942\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__31945\,
            I => \N__31939\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__31942\,
            I => \N__31936\
        );

    \I__6435\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31932\
        );

    \I__6434\ : Span4Mux_h
    port map (
            O => \N__31936\,
            I => \N__31929\
        );

    \I__6433\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31926\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__31932\,
            I => \acadc_skipCount_2\
        );

    \I__6431\ : Odrv4
    port map (
            O => \N__31929\,
            I => \acadc_skipCount_2\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__31926\,
            I => \acadc_skipCount_2\
        );

    \I__6429\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31916\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__31916\,
            I => n22_adj_1170
        );

    \I__6427\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31908\
        );

    \I__6426\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31903\
        );

    \I__6425\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31903\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31900\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__31903\,
            I => req_data_cnt_14
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__31900\,
            I => req_data_cnt_14
        );

    \I__6421\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31892\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__31892\,
            I => n23_adj_1194
        );

    \I__6419\ : InMux
    port map (
            O => \N__31889\,
            I => \N__31886\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__31886\,
            I => \N__31881\
        );

    \I__6417\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31876\
        );

    \I__6416\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31876\
        );

    \I__6415\ : Odrv4
    port map (
            O => \N__31881\,
            I => \acadc_skipCount_4\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__31876\,
            I => \acadc_skipCount_4\
        );

    \I__6413\ : InMux
    port map (
            O => \N__31871\,
            I => \N__31866\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__31870\,
            I => \N__31863\
        );

    \I__6411\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31859\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31856\
        );

    \I__6409\ : InMux
    port map (
            O => \N__31863\,
            I => \N__31853\
        );

    \I__6408\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31850\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__31859\,
            I => \N__31843\
        );

    \I__6406\ : Span4Mux_h
    port map (
            O => \N__31856\,
            I => \N__31838\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__31853\,
            I => \N__31838\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__31850\,
            I => \N__31835\
        );

    \I__6403\ : InMux
    port map (
            O => \N__31849\,
            I => \N__31832\
        );

    \I__6402\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31829\
        );

    \I__6401\ : InMux
    port map (
            O => \N__31847\,
            I => \N__31824\
        );

    \I__6400\ : InMux
    port map (
            O => \N__31846\,
            I => \N__31824\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__31843\,
            I => \N__31819\
        );

    \I__6398\ : Span4Mux_v
    port map (
            O => \N__31838\,
            I => \N__31819\
        );

    \I__6397\ : Span4Mux_v
    port map (
            O => \N__31835\,
            I => \N__31816\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__31832\,
            I => n9224
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__31829\,
            I => n9224
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__31824\,
            I => n9224
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__31819\,
            I => n9224
        );

    \I__6392\ : Odrv4
    port map (
            O => \N__31816\,
            I => n9224
        );

    \I__6391\ : InMux
    port map (
            O => \N__31805\,
            I => \N__31802\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__31802\,
            I => \N__31799\
        );

    \I__6389\ : Span4Mux_h
    port map (
            O => \N__31799\,
            I => \N__31795\
        );

    \I__6388\ : InMux
    port map (
            O => \N__31798\,
            I => \N__31792\
        );

    \I__6387\ : Span4Mux_v
    port map (
            O => \N__31795\,
            I => \N__31789\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__31792\,
            I => buf_device_acadc_5
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__31789\,
            I => buf_device_acadc_5
        );

    \I__6384\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31775\
        );

    \I__6383\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31775\
        );

    \I__6382\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31775\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__31775\,
            I => \acadc_skipCount_9\
        );

    \I__6380\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31769\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__31769\,
            I => \N__31766\
        );

    \I__6378\ : Span4Mux_h
    port map (
            O => \N__31766\,
            I => \N__31763\
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__31763\,
            I => n15834
        );

    \I__6376\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31757\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__31757\,
            I => \N__31754\
        );

    \I__6374\ : Span4Mux_v
    port map (
            O => \N__31754\,
            I => \N__31751\
        );

    \I__6373\ : Span4Mux_h
    port map (
            O => \N__31751\,
            I => \N__31748\
        );

    \I__6372\ : Odrv4
    port map (
            O => \N__31748\,
            I => n19_adj_1234
        );

    \I__6371\ : CascadeMux
    port map (
            O => \N__31745\,
            I => \n20_adj_1253_cascade_\
        );

    \I__6370\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31739\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__31739\,
            I => \N__31736\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__31736\,
            I => \N__31733\
        );

    \I__6367\ : Odrv4
    port map (
            O => \N__31733\,
            I => n29
        );

    \I__6366\ : InMux
    port map (
            O => \N__31730\,
            I => \N__31723\
        );

    \I__6365\ : InMux
    port map (
            O => \N__31729\,
            I => \N__31723\
        );

    \I__6364\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31720\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31717\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__31720\,
            I => buf_dds_7
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__31717\,
            I => buf_dds_7
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__31712\,
            I => \N__31709\
        );

    \I__6359\ : InMux
    port map (
            O => \N__31709\,
            I => \N__31706\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__31706\,
            I => \N__31696\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__31705\,
            I => \N__31693\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__31704\,
            I => \N__31690\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__31703\,
            I => \N__31687\
        );

    \I__6354\ : CascadeMux
    port map (
            O => \N__31702\,
            I => \N__31684\
        );

    \I__6353\ : CascadeMux
    port map (
            O => \N__31701\,
            I => \N__31681\
        );

    \I__6352\ : CascadeMux
    port map (
            O => \N__31700\,
            I => \N__31678\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__31699\,
            I => \N__31675\
        );

    \I__6350\ : Span4Mux_v
    port map (
            O => \N__31696\,
            I => \N__31670\
        );

    \I__6349\ : InMux
    port map (
            O => \N__31693\,
            I => \N__31663\
        );

    \I__6348\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31663\
        );

    \I__6347\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31663\
        );

    \I__6346\ : InMux
    port map (
            O => \N__31684\,
            I => \N__31654\
        );

    \I__6345\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31654\
        );

    \I__6344\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31654\
        );

    \I__6343\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31654\
        );

    \I__6342\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31651\
        );

    \I__6341\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31648\
        );

    \I__6340\ : Span4Mux_h
    port map (
            O => \N__31670\,
            I => \N__31641\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__31663\,
            I => \N__31641\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__31654\,
            I => \N__31641\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31634\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__31648\,
            I => \N__31634\
        );

    \I__6335\ : Span4Mux_v
    port map (
            O => \N__31641\,
            I => \N__31634\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__31634\,
            I => n7567
        );

    \I__6333\ : InMux
    port map (
            O => \N__31631\,
            I => \N__31628\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__31628\,
            I => n21_adj_1204
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__31625\,
            I => \N__31621\
        );

    \I__6330\ : InMux
    port map (
            O => \N__31624\,
            I => \N__31618\
        );

    \I__6329\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31614\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__31618\,
            I => \N__31611\
        );

    \I__6327\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31608\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__31614\,
            I => \N__31605\
        );

    \I__6325\ : Span4Mux_v
    port map (
            O => \N__31611\,
            I => \N__31602\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__31608\,
            I => \N__31599\
        );

    \I__6323\ : Span4Mux_v
    port map (
            O => \N__31605\,
            I => \N__31594\
        );

    \I__6322\ : Span4Mux_h
    port map (
            O => \N__31602\,
            I => \N__31589\
        );

    \I__6321\ : Span4Mux_v
    port map (
            O => \N__31599\,
            I => \N__31589\
        );

    \I__6320\ : InMux
    port map (
            O => \N__31598\,
            I => \N__31584\
        );

    \I__6319\ : InMux
    port map (
            O => \N__31597\,
            I => \N__31584\
        );

    \I__6318\ : Odrv4
    port map (
            O => \N__31594\,
            I => comm_buf_1_4
        );

    \I__6317\ : Odrv4
    port map (
            O => \N__31589\,
            I => comm_buf_1_4
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__31584\,
            I => comm_buf_1_4
        );

    \I__6315\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31572\
        );

    \I__6314\ : InMux
    port map (
            O => \N__31576\,
            I => \N__31569\
        );

    \I__6313\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31566\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__31572\,
            I => \N__31563\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__31569\,
            I => \N__31560\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__31566\,
            I => buf_dds_4
        );

    \I__6309\ : Odrv12
    port map (
            O => \N__31563\,
            I => buf_dds_4
        );

    \I__6308\ : Odrv4
    port map (
            O => \N__31560\,
            I => buf_dds_4
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__31553\,
            I => \N__31550\
        );

    \I__6306\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31546\
        );

    \I__6305\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31543\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__31546\,
            I => \N__31540\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__31543\,
            I => buf_control_5
        );

    \I__6302\ : Odrv4
    port map (
            O => \N__31540\,
            I => buf_control_5
        );

    \I__6301\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31532\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__31532\,
            I => \N__31529\
        );

    \I__6299\ : Span4Mux_h
    port map (
            O => \N__31529\,
            I => \N__31526\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__31526\,
            I => \N__31523\
        );

    \I__6297\ : Odrv4
    port map (
            O => \N__31523\,
            I => buf_data1_10
        );

    \I__6296\ : CascadeMux
    port map (
            O => \N__31520\,
            I => \n4195_cascade_\
        );

    \I__6295\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31514\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__31514\,
            I => n4232
        );

    \I__6293\ : InMux
    port map (
            O => \N__31511\,
            I => \N__31508\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__31508\,
            I => \N__31504\
        );

    \I__6291\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31501\
        );

    \I__6290\ : Span4Mux_h
    port map (
            O => \N__31504\,
            I => \N__31498\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__31501\,
            I => acadc_skipcnt_9
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__31498\,
            I => acadc_skipcnt_9
        );

    \I__6287\ : CascadeMux
    port map (
            O => \N__31493\,
            I => \N__31490\
        );

    \I__6286\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31487\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__31487\,
            I => \N__31483\
        );

    \I__6284\ : InMux
    port map (
            O => \N__31486\,
            I => \N__31480\
        );

    \I__6283\ : Span12Mux_v
    port map (
            O => \N__31483\,
            I => \N__31477\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__31480\,
            I => acadc_skipcnt_15
        );

    \I__6281\ : Odrv12
    port map (
            O => \N__31477\,
            I => acadc_skipcnt_15
        );

    \I__6280\ : InMux
    port map (
            O => \N__31472\,
            I => \N__31469\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__31469\,
            I => n24_adj_1174
        );

    \I__6278\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31463\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__31463\,
            I => n4247
        );

    \I__6276\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31457\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__31457\,
            I => \N__31453\
        );

    \I__6274\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31449\
        );

    \I__6273\ : Span4Mux_v
    port map (
            O => \N__31453\,
            I => \N__31446\
        );

    \I__6272\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31443\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__31449\,
            I => \N__31440\
        );

    \I__6270\ : Span4Mux_v
    port map (
            O => \N__31446\,
            I => \N__31437\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__31443\,
            I => buf_dds_15
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__31440\,
            I => buf_dds_15
        );

    \I__6267\ : Odrv4
    port map (
            O => \N__31437\,
            I => buf_dds_15
        );

    \I__6266\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31427\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__31427\,
            I => \N__31424\
        );

    \I__6264\ : Span12Mux_v
    port map (
            O => \N__31424\,
            I => \N__31419\
        );

    \I__6263\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31414\
        );

    \I__6262\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31414\
        );

    \I__6261\ : Odrv12
    port map (
            O => \N__31419\,
            I => req_data_cnt_13
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__31414\,
            I => req_data_cnt_13
        );

    \I__6259\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31404\
        );

    \I__6258\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31399\
        );

    \I__6257\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31399\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__31404\,
            I => req_data_cnt_8
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__31399\,
            I => req_data_cnt_8
        );

    \I__6254\ : CascadeMux
    port map (
            O => \N__31394\,
            I => \N__31391\
        );

    \I__6253\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31388\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31385\
        );

    \I__6251\ : Odrv12
    port map (
            O => \N__31385\,
            I => n15812
        );

    \I__6250\ : InMux
    port map (
            O => \N__31382\,
            I => \N__31379\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__31379\,
            I => \N__31375\
        );

    \I__6248\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31372\
        );

    \I__6247\ : Span4Mux_v
    port map (
            O => \N__31375\,
            I => \N__31369\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__31372\,
            I => buf_device_acadc_6
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__31369\,
            I => buf_device_acadc_6
        );

    \I__6244\ : CascadeMux
    port map (
            O => \N__31364\,
            I => \N__31361\
        );

    \I__6243\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31358\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__31358\,
            I => \N__31355\
        );

    \I__6241\ : Span4Mux_h
    port map (
            O => \N__31355\,
            I => \N__31352\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__31352\,
            I => buf_data1_16
        );

    \I__6239\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31346\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__31346\,
            I => \N__31343\
        );

    \I__6237\ : Span4Mux_h
    port map (
            O => \N__31343\,
            I => \N__31340\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__31340\,
            I => n99
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__31337\,
            I => \N__31332\
        );

    \I__6234\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31329\
        );

    \I__6233\ : InMux
    port map (
            O => \N__31335\,
            I => \N__31326\
        );

    \I__6232\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31323\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__31329\,
            I => req_data_cnt_7
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__31326\,
            I => req_data_cnt_7
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__31323\,
            I => req_data_cnt_7
        );

    \I__6228\ : InMux
    port map (
            O => \N__31316\,
            I => \N__31313\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__31313\,
            I => \N__31310\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__31310\,
            I => n4214
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__31307\,
            I => \N__31304\
        );

    \I__6224\ : InMux
    port map (
            O => \N__31304\,
            I => \N__31301\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__31301\,
            I => \N__31298\
        );

    \I__6222\ : Span4Mux_v
    port map (
            O => \N__31298\,
            I => \N__31295\
        );

    \I__6221\ : Odrv4
    port map (
            O => \N__31295\,
            I => n15556
        );

    \I__6220\ : InMux
    port map (
            O => \N__31292\,
            I => \N__31289\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__31289\,
            I => \N__31286\
        );

    \I__6218\ : Span12Mux_h
    port map (
            O => \N__31286\,
            I => \N__31283\
        );

    \I__6217\ : Odrv12
    port map (
            O => \N__31283\,
            I => n60_adj_1157
        );

    \I__6216\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31277\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__31277\,
            I => \N__31274\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__31274\,
            I => n4252
        );

    \I__6213\ : CascadeMux
    port map (
            O => \N__31271\,
            I => \N__31268\
        );

    \I__6212\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31265\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__31265\,
            I => n4202
        );

    \I__6210\ : CascadeMux
    port map (
            O => \N__31262\,
            I => \N__31259\
        );

    \I__6209\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31256\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__31256\,
            I => \CLOCK_DDS.tmp_buf_2\
        );

    \I__6207\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31250\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__31250\,
            I => \N__31247\
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__31247\,
            I => \CLOCK_DDS.tmp_buf_3\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__31244\,
            I => \N__31241\
        );

    \I__6203\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31238\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__31238\,
            I => \CLOCK_DDS.tmp_buf_4\
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__31235\,
            I => \N__31232\
        );

    \I__6200\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31229\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__31229\,
            I => \CLOCK_DDS.tmp_buf_5\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__31226\,
            I => \N__31223\
        );

    \I__6197\ : InMux
    port map (
            O => \N__31223\,
            I => \N__31220\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__31220\,
            I => \CLOCK_DDS.tmp_buf_6\
        );

    \I__6195\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31214\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__31214\,
            I => \CLOCK_DDS.tmp_buf_7\
        );

    \I__6193\ : CEMux
    port map (
            O => \N__31211\,
            I => \N__31206\
        );

    \I__6192\ : CEMux
    port map (
            O => \N__31210\,
            I => \N__31203\
        );

    \I__6191\ : CEMux
    port map (
            O => \N__31209\,
            I => \N__31200\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__31206\,
            I => \CLOCK_DDS.n9759\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__31203\,
            I => \CLOCK_DDS.n9759\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__31200\,
            I => \CLOCK_DDS.n9759\
        );

    \I__6187\ : SRMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__31190\,
            I => \N__31186\
        );

    \I__6185\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31183\
        );

    \I__6184\ : Span4Mux_v
    port map (
            O => \N__31186\,
            I => \N__31180\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31177\
        );

    \I__6182\ : Span4Mux_h
    port map (
            O => \N__31180\,
            I => \N__31174\
        );

    \I__6181\ : Span4Mux_h
    port map (
            O => \N__31177\,
            I => \N__31171\
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__31174\,
            I => n10823
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__31171\,
            I => n10823
        );

    \I__6178\ : CEMux
    port map (
            O => \N__31166\,
            I => \N__31163\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__6176\ : Span4Mux_h
    port map (
            O => \N__31160\,
            I => \N__31157\
        );

    \I__6175\ : Span4Mux_v
    port map (
            O => \N__31157\,
            I => \N__31154\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__31154\,
            I => \CLOCK_DDS.n9_adj_1021\
        );

    \I__6173\ : InMux
    port map (
            O => \N__31151\,
            I => \N__31148\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__31148\,
            I => \N__31145\
        );

    \I__6171\ : Span4Mux_v
    port map (
            O => \N__31145\,
            I => \N__31139\
        );

    \I__6170\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31132\
        );

    \I__6169\ : InMux
    port map (
            O => \N__31143\,
            I => \N__31132\
        );

    \I__6168\ : InMux
    port map (
            O => \N__31142\,
            I => \N__31132\
        );

    \I__6167\ : Span4Mux_h
    port map (
            O => \N__31139\,
            I => \N__31129\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__31132\,
            I => bit_cnt_1
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__31129\,
            I => bit_cnt_1
        );

    \I__6164\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31120\
        );

    \I__6163\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31117\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31112\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__31117\,
            I => \N__31112\
        );

    \I__6160\ : Odrv12
    port map (
            O => \N__31112\,
            I => n15176
        );

    \I__6159\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31106\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__31106\,
            I => \N__31103\
        );

    \I__6157\ : Span4Mux_v
    port map (
            O => \N__31103\,
            I => \N__31100\
        );

    \I__6156\ : Sp12to4
    port map (
            O => \N__31100\,
            I => \N__31097\
        );

    \I__6155\ : Odrv12
    port map (
            O => \N__31097\,
            I => n15396
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__31094\,
            I => \N__31091\
        );

    \I__6153\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31088\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__31088\,
            I => \N__31085\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__31085\,
            I => n15670
        );

    \I__6150\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31076\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__31076\,
            I => \N__31070\
        );

    \I__6147\ : InMux
    port map (
            O => \N__31075\,
            I => \N__31065\
        );

    \I__6146\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31065\
        );

    \I__6145\ : InMux
    port map (
            O => \N__31073\,
            I => \N__31062\
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__31070\,
            I => n13475
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__31065\,
            I => n13475
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__31062\,
            I => n13475
        );

    \I__6141\ : InMux
    port map (
            O => \N__31055\,
            I => \N__31052\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__6139\ : Odrv4
    port map (
            O => \N__31049\,
            I => n15_adj_1203
        );

    \I__6138\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31043\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__6136\ : Span4Mux_v
    port map (
            O => \N__31040\,
            I => \N__31037\
        );

    \I__6135\ : Span4Mux_h
    port map (
            O => \N__31037\,
            I => \N__31033\
        );

    \I__6134\ : InMux
    port map (
            O => \N__31036\,
            I => \N__31030\
        );

    \I__6133\ : Odrv4
    port map (
            O => \N__31033\,
            I => tmp_buf_15
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__31030\,
            I => tmp_buf_15
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__31025\,
            I => \N__31022\
        );

    \I__6130\ : InMux
    port map (
            O => \N__31022\,
            I => \N__31019\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__31019\,
            I => \CLOCK_DDS.tmp_buf_0\
        );

    \I__6128\ : CascadeMux
    port map (
            O => \N__31016\,
            I => \N__31013\
        );

    \I__6127\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31010\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__31010\,
            I => \CLOCK_DDS.tmp_buf_1\
        );

    \I__6125\ : SRMux
    port map (
            O => \N__31007\,
            I => \N__31004\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__31004\,
            I => \N__31001\
        );

    \I__6123\ : Span4Mux_v
    port map (
            O => \N__31001\,
            I => \N__30997\
        );

    \I__6122\ : SRMux
    port map (
            O => \N__31000\,
            I => \N__30993\
        );

    \I__6121\ : Sp12to4
    port map (
            O => \N__30997\,
            I => \N__30990\
        );

    \I__6120\ : SRMux
    port map (
            O => \N__30996\,
            I => \N__30987\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30984\
        );

    \I__6118\ : Span12Mux_h
    port map (
            O => \N__30990\,
            I => \N__30979\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__30987\,
            I => \N__30979\
        );

    \I__6116\ : Span4Mux_h
    port map (
            O => \N__30984\,
            I => \N__30976\
        );

    \I__6115\ : Odrv12
    port map (
            O => \N__30979\,
            I => \comm_spi.data_tx_7__N_813\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__30976\,
            I => \comm_spi.data_tx_7__N_813\
        );

    \I__6113\ : InMux
    port map (
            O => \N__30971\,
            I => \N__30968\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30964\
        );

    \I__6111\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30961\
        );

    \I__6110\ : Span4Mux_v
    port map (
            O => \N__30964\,
            I => \N__30958\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30955\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__30958\,
            I => \N__30951\
        );

    \I__6107\ : Span4Mux_v
    port map (
            O => \N__30955\,
            I => \N__30948\
        );

    \I__6106\ : InMux
    port map (
            O => \N__30954\,
            I => \N__30945\
        );

    \I__6105\ : Sp12to4
    port map (
            O => \N__30951\,
            I => \N__30938\
        );

    \I__6104\ : Sp12to4
    port map (
            O => \N__30948\,
            I => \N__30938\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30938\
        );

    \I__6102\ : Span12Mux_h
    port map (
            O => \N__30938\,
            I => \N__30935\
        );

    \I__6101\ : Odrv12
    port map (
            O => \N__30935\,
            I => comm_tx_buf_3
        );

    \I__6100\ : SRMux
    port map (
            O => \N__30932\,
            I => \N__30929\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__30929\,
            I => \N__30926\
        );

    \I__6098\ : Span4Mux_v
    port map (
            O => \N__30926\,
            I => \N__30923\
        );

    \I__6097\ : Span4Mux_h
    port map (
            O => \N__30923\,
            I => \N__30920\
        );

    \I__6096\ : Odrv4
    port map (
            O => \N__30920\,
            I => \comm_spi.data_tx_7__N_825\
        );

    \I__6095\ : InMux
    port map (
            O => \N__30917\,
            I => \N__30914\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__30914\,
            I => \N__30911\
        );

    \I__6093\ : Span4Mux_v
    port map (
            O => \N__30911\,
            I => \N__30908\
        );

    \I__6092\ : Span4Mux_h
    port map (
            O => \N__30908\,
            I => \N__30905\
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__30905\,
            I => buf_data1_22
        );

    \I__6090\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30899\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__30899\,
            I => \N__30896\
        );

    \I__6088\ : Span12Mux_h
    port map (
            O => \N__30896\,
            I => \N__30893\
        );

    \I__6087\ : Odrv12
    port map (
            O => \N__30893\,
            I => n66
        );

    \I__6086\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30887\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__30887\,
            I => \N__30883\
        );

    \I__6084\ : InMux
    port map (
            O => \N__30886\,
            I => \N__30880\
        );

    \I__6083\ : Span4Mux_h
    port map (
            O => \N__30883\,
            I => \N__30877\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30874\
        );

    \I__6081\ : Span4Mux_h
    port map (
            O => \N__30877\,
            I => \N__30871\
        );

    \I__6080\ : Span12Mux_h
    port map (
            O => \N__30874\,
            I => \N__30868\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__30871\,
            I => \comm_spi.n10452\
        );

    \I__6078\ : Odrv12
    port map (
            O => \N__30868\,
            I => \comm_spi.n10452\
        );

    \I__6077\ : InMux
    port map (
            O => \N__30863\,
            I => \N__30860\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__30860\,
            I => \N__30857\
        );

    \I__6075\ : Span4Mux_v
    port map (
            O => \N__30857\,
            I => \N__30853\
        );

    \I__6074\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30850\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__30853\,
            I => \comm_spi.n10451\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__30850\,
            I => \comm_spi.n10451\
        );

    \I__6071\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30839\
        );

    \I__6070\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30836\
        );

    \I__6069\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30831\
        );

    \I__6068\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30828\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__30839\,
            I => \N__30825\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__30836\,
            I => \N__30822\
        );

    \I__6065\ : InMux
    port map (
            O => \N__30835\,
            I => \N__30819\
        );

    \I__6064\ : InMux
    port map (
            O => \N__30834\,
            I => \N__30816\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__30831\,
            I => \N__30813\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30810\
        );

    \I__6061\ : Span12Mux_v
    port map (
            O => \N__30825\,
            I => \N__30807\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__30822\,
            I => \N__30800\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__30819\,
            I => \N__30800\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__30816\,
            I => \N__30800\
        );

    \I__6057\ : Span4Mux_v
    port map (
            O => \N__30813\,
            I => \N__30795\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__30810\,
            I => \N__30795\
        );

    \I__6055\ : Odrv12
    port map (
            O => \N__30807\,
            I => \comm_spi.n10444\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__30800\,
            I => \comm_spi.n10444\
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__30795\,
            I => \comm_spi.n10444\
        );

    \I__6052\ : InMux
    port map (
            O => \N__30788\,
            I => \N__30785\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__30785\,
            I => \N__30782\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__30782\,
            I => \comm_spi.n10445\
        );

    \I__6049\ : SRMux
    port map (
            O => \N__30779\,
            I => \N__30775\
        );

    \I__6048\ : SRMux
    port map (
            O => \N__30778\,
            I => \N__30772\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__30775\,
            I => \N__30769\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__30772\,
            I => \N__30765\
        );

    \I__6045\ : Span4Mux_h
    port map (
            O => \N__30769\,
            I => \N__30762\
        );

    \I__6044\ : SRMux
    port map (
            O => \N__30768\,
            I => \N__30759\
        );

    \I__6043\ : Span4Mux_h
    port map (
            O => \N__30765\,
            I => \N__30756\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__30762\,
            I => \N__30751\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30751\
        );

    \I__6040\ : Span4Mux_h
    port map (
            O => \N__30756\,
            I => \N__30748\
        );

    \I__6039\ : Odrv4
    port map (
            O => \N__30751\,
            I => \comm_spi.data_tx_7__N_805\
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__30748\,
            I => \comm_spi.data_tx_7__N_805\
        );

    \I__6037\ : SRMux
    port map (
            O => \N__30743\,
            I => \N__30740\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__30740\,
            I => \N__30737\
        );

    \I__6035\ : Span4Mux_h
    port map (
            O => \N__30737\,
            I => \N__30733\
        );

    \I__6034\ : SRMux
    port map (
            O => \N__30736\,
            I => \N__30730\
        );

    \I__6033\ : Span4Mux_h
    port map (
            O => \N__30733\,
            I => \N__30727\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__30730\,
            I => \N__30724\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__30727\,
            I => \N__30721\
        );

    \I__6030\ : Span4Mux_h
    port map (
            O => \N__30724\,
            I => \N__30718\
        );

    \I__6029\ : Sp12to4
    port map (
            O => \N__30721\,
            I => \N__30715\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__30718\,
            I => \N__30712\
        );

    \I__6027\ : Odrv12
    port map (
            O => \N__30715\,
            I => n10640
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__30712\,
            I => n10640
        );

    \I__6025\ : SRMux
    port map (
            O => \N__30707\,
            I => \N__30704\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__30704\,
            I => \N__30700\
        );

    \I__6023\ : SRMux
    port map (
            O => \N__30703\,
            I => \N__30697\
        );

    \I__6022\ : Span4Mux_v
    port map (
            O => \N__30700\,
            I => \N__30692\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__30697\,
            I => \N__30692\
        );

    \I__6020\ : Sp12to4
    port map (
            O => \N__30692\,
            I => \N__30689\
        );

    \I__6019\ : Odrv12
    port map (
            O => \N__30689\,
            I => n10532
        );

    \I__6018\ : SRMux
    port map (
            O => \N__30686\,
            I => \N__30683\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__30680\,
            I => \N__30677\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__30677\,
            I => n15344
        );

    \I__6014\ : InMux
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__30671\,
            I => \N__30668\
        );

    \I__6012\ : Span12Mux_h
    port map (
            O => \N__30668\,
            I => \N__30665\
        );

    \I__6011\ : Odrv12
    port map (
            O => \N__30665\,
            I => n15171
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__30662\,
            I => \n15328_cascade_\
        );

    \I__6009\ : InMux
    port map (
            O => \N__30659\,
            I => \N__30649\
        );

    \I__6008\ : InMux
    port map (
            O => \N__30658\,
            I => \N__30649\
        );

    \I__6007\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30642\
        );

    \I__6006\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30642\
        );

    \I__6005\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30637\
        );

    \I__6004\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30637\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30633\
        );

    \I__6002\ : InMux
    port map (
            O => \N__30648\,
            I => \N__30630\
        );

    \I__6001\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30627\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__30642\,
            I => \N__30622\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__30637\,
            I => \N__30622\
        );

    \I__5998\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30619\
        );

    \I__5997\ : Span4Mux_h
    port map (
            O => \N__30633\,
            I => \N__30615\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__30630\,
            I => \N__30610\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30610\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__30622\,
            I => \N__30605\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__30619\,
            I => \N__30605\
        );

    \I__5992\ : InMux
    port map (
            O => \N__30618\,
            I => \N__30601\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__30615\,
            I => \N__30598\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__30610\,
            I => \N__30595\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__30605\,
            I => \N__30592\
        );

    \I__5988\ : InMux
    port map (
            O => \N__30604\,
            I => \N__30589\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__30601\,
            I => acadc_trig
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__30598\,
            I => acadc_trig
        );

    \I__5985\ : Odrv4
    port map (
            O => \N__30595\,
            I => acadc_trig
        );

    \I__5984\ : Odrv4
    port map (
            O => \N__30592\,
            I => acadc_trig
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__30589\,
            I => acadc_trig
        );

    \I__5982\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30573\
        );

    \I__5981\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30570\
        );

    \I__5980\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30567\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30560\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__30570\,
            I => \N__30560\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__30567\,
            I => \N__30560\
        );

    \I__5976\ : Span4Mux_v
    port map (
            O => \N__30560\,
            I => \N__30557\
        );

    \I__5975\ : Span4Mux_v
    port map (
            O => \N__30557\,
            I => \N__30554\
        );

    \I__5974\ : Odrv4
    port map (
            O => \N__30554\,
            I => data_index_6
        );

    \I__5973\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30548\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__30548\,
            I => \N__30545\
        );

    \I__5971\ : Odrv12
    port map (
            O => \N__30545\,
            I => n8_adj_1221
        );

    \I__5970\ : InMux
    port map (
            O => \N__30542\,
            I => \N__30538\
        );

    \I__5969\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30535\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__30538\,
            I => \N__30532\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__30535\,
            I => \N__30529\
        );

    \I__5966\ : Odrv12
    port map (
            O => \N__30532\,
            I => n7_adj_1220
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__30529\,
            I => n7_adj_1220
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__30524\,
            I => \N__30521\
        );

    \I__5963\ : CascadeBuf
    port map (
            O => \N__30521\,
            I => \N__30518\
        );

    \I__5962\ : CascadeMux
    port map (
            O => \N__30518\,
            I => \N__30515\
        );

    \I__5961\ : CascadeBuf
    port map (
            O => \N__30515\,
            I => \N__30512\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__30512\,
            I => \N__30509\
        );

    \I__5959\ : CascadeBuf
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__30506\,
            I => \N__30503\
        );

    \I__5957\ : CascadeBuf
    port map (
            O => \N__30503\,
            I => \N__30500\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__30500\,
            I => \N__30497\
        );

    \I__5955\ : CascadeBuf
    port map (
            O => \N__30497\,
            I => \N__30494\
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__30494\,
            I => \N__30491\
        );

    \I__5953\ : CascadeBuf
    port map (
            O => \N__30491\,
            I => \N__30488\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__30488\,
            I => \N__30485\
        );

    \I__5951\ : CascadeBuf
    port map (
            O => \N__30485\,
            I => \N__30482\
        );

    \I__5950\ : CascadeMux
    port map (
            O => \N__30482\,
            I => \N__30478\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__30481\,
            I => \N__30475\
        );

    \I__5948\ : CascadeBuf
    port map (
            O => \N__30478\,
            I => \N__30472\
        );

    \I__5947\ : CascadeBuf
    port map (
            O => \N__30475\,
            I => \N__30469\
        );

    \I__5946\ : CascadeMux
    port map (
            O => \N__30472\,
            I => \N__30466\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__30469\,
            I => \N__30463\
        );

    \I__5944\ : CascadeBuf
    port map (
            O => \N__30466\,
            I => \N__30460\
        );

    \I__5943\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30457\
        );

    \I__5942\ : CascadeMux
    port map (
            O => \N__30460\,
            I => \N__30454\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__30457\,
            I => \N__30451\
        );

    \I__5940\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30448\
        );

    \I__5939\ : Span12Mux_h
    port map (
            O => \N__30451\,
            I => \N__30445\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__30448\,
            I => \N__30442\
        );

    \I__5937\ : Span12Mux_v
    port map (
            O => \N__30445\,
            I => \N__30439\
        );

    \I__5936\ : Span4Mux_h
    port map (
            O => \N__30442\,
            I => \N__30436\
        );

    \I__5935\ : Odrv12
    port map (
            O => \N__30439\,
            I => \data_index_9_N_258_7\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__30436\,
            I => \data_index_9_N_258_7\
        );

    \I__5933\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30428\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__5931\ : Span4Mux_v
    port map (
            O => \N__30425\,
            I => \N__30421\
        );

    \I__5930\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30418\
        );

    \I__5929\ : Span4Mux_v
    port map (
            O => \N__30421\,
            I => \N__30413\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30413\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__30413\,
            I => n7_adj_1222
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__30410\,
            I => \N__30407\
        );

    \I__5925\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30404\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__30404\,
            I => \N__30401\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__30401\,
            I => \N__30398\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__30398\,
            I => \N__30394\
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__30397\,
            I => \N__30391\
        );

    \I__5920\ : Span4Mux_v
    port map (
            O => \N__30394\,
            I => \N__30388\
        );

    \I__5919\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30385\
        );

    \I__5918\ : Odrv4
    port map (
            O => \N__30388\,
            I => n8_adj_1223
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__30385\,
            I => n8_adj_1223
        );

    \I__5916\ : CascadeMux
    port map (
            O => \N__30380\,
            I => \N__30377\
        );

    \I__5915\ : CascadeBuf
    port map (
            O => \N__30377\,
            I => \N__30374\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__30374\,
            I => \N__30371\
        );

    \I__5913\ : CascadeBuf
    port map (
            O => \N__30371\,
            I => \N__30368\
        );

    \I__5912\ : CascadeMux
    port map (
            O => \N__30368\,
            I => \N__30365\
        );

    \I__5911\ : CascadeBuf
    port map (
            O => \N__30365\,
            I => \N__30362\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__30362\,
            I => \N__30359\
        );

    \I__5909\ : CascadeBuf
    port map (
            O => \N__30359\,
            I => \N__30356\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__30356\,
            I => \N__30353\
        );

    \I__5907\ : CascadeBuf
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__5906\ : CascadeMux
    port map (
            O => \N__30350\,
            I => \N__30347\
        );

    \I__5905\ : CascadeBuf
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__5903\ : CascadeBuf
    port map (
            O => \N__30341\,
            I => \N__30337\
        );

    \I__5902\ : CascadeMux
    port map (
            O => \N__30340\,
            I => \N__30334\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \N__30331\
        );

    \I__5900\ : CascadeBuf
    port map (
            O => \N__30334\,
            I => \N__30328\
        );

    \I__5899\ : CascadeBuf
    port map (
            O => \N__30331\,
            I => \N__30325\
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__30328\,
            I => \N__30322\
        );

    \I__5897\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30319\
        );

    \I__5896\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30316\
        );

    \I__5895\ : CascadeBuf
    port map (
            O => \N__30319\,
            I => \N__30313\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30310\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__30313\,
            I => \N__30307\
        );

    \I__5892\ : Span12Mux_s9_h
    port map (
            O => \N__30310\,
            I => \N__30304\
        );

    \I__5891\ : InMux
    port map (
            O => \N__30307\,
            I => \N__30301\
        );

    \I__5890\ : Span12Mux_v
    port map (
            O => \N__30304\,
            I => \N__30298\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__30301\,
            I => \N__30295\
        );

    \I__5888\ : Odrv12
    port map (
            O => \N__30298\,
            I => \data_index_9_N_258_6\
        );

    \I__5887\ : Odrv12
    port map (
            O => \N__30295\,
            I => \data_index_9_N_258_6\
        );

    \I__5886\ : IoInMux
    port map (
            O => \N__30290\,
            I => \N__30287\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__30287\,
            I => \N__30284\
        );

    \I__5884\ : Span4Mux_s3_h
    port map (
            O => \N__30284\,
            I => \N__30281\
        );

    \I__5883\ : Sp12to4
    port map (
            O => \N__30281\,
            I => \N__30278\
        );

    \I__5882\ : Span12Mux_s9_v
    port map (
            O => \N__30278\,
            I => \N__30275\
        );

    \I__5881\ : Odrv12
    port map (
            O => \N__30275\,
            I => \ICE_SPI_MISO\
        );

    \I__5880\ : InMux
    port map (
            O => \N__30272\,
            I => \N__30269\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__30269\,
            I => \comm_spi.n10446\
        );

    \I__5878\ : InMux
    port map (
            O => \N__30266\,
            I => n14035
        );

    \I__5877\ : InMux
    port map (
            O => \N__30263\,
            I => n14036
        );

    \I__5876\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30255\
        );

    \I__5875\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30252\
        );

    \I__5874\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30249\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__30255\,
            I => \N__30244\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__30252\,
            I => \N__30244\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__30249\,
            I => data_index_7
        );

    \I__5870\ : Odrv12
    port map (
            O => \N__30244\,
            I => data_index_7
        );

    \I__5869\ : InMux
    port map (
            O => \N__30239\,
            I => n14037
        );

    \I__5868\ : InMux
    port map (
            O => \N__30236\,
            I => \bfn_14_17_0_\
        );

    \I__5867\ : InMux
    port map (
            O => \N__30233\,
            I => \N__30228\
        );

    \I__5866\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30225\
        );

    \I__5865\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30222\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__30228\,
            I => data_index_3
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__30225\,
            I => data_index_3
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__30222\,
            I => data_index_3
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__30215\,
            I => \N__30209\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__30214\,
            I => \N__30206\
        );

    \I__5859\ : CascadeMux
    port map (
            O => \N__30213\,
            I => \N__30203\
        );

    \I__5858\ : InMux
    port map (
            O => \N__30212\,
            I => \N__30200\
        );

    \I__5857\ : InMux
    port map (
            O => \N__30209\,
            I => \N__30193\
        );

    \I__5856\ : InMux
    port map (
            O => \N__30206\,
            I => \N__30193\
        );

    \I__5855\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30193\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__30200\,
            I => \N__30190\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__30193\,
            I => \N__30187\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__30190\,
            I => \N__30182\
        );

    \I__5851\ : Span4Mux_v
    port map (
            O => \N__30187\,
            I => \N__30179\
        );

    \I__5850\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30174\
        );

    \I__5849\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30174\
        );

    \I__5848\ : Span4Mux_h
    port map (
            O => \N__30182\,
            I => \N__30171\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__30179\,
            I => \N__30168\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__30174\,
            I => \N__30165\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__30171\,
            I => \N__30162\
        );

    \I__5844\ : Span4Mux_h
    port map (
            O => \N__30168\,
            I => \N__30159\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__30165\,
            I => \N__30156\
        );

    \I__5842\ : Sp12to4
    port map (
            O => \N__30162\,
            I => \N__30151\
        );

    \I__5841\ : Sp12to4
    port map (
            O => \N__30159\,
            I => \N__30151\
        );

    \I__5840\ : Span4Mux_v
    port map (
            O => \N__30156\,
            I => \N__30148\
        );

    \I__5839\ : Odrv12
    port map (
            O => \N__30151\,
            I => \M_DRDY2\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__30148\,
            I => \M_DRDY2\
        );

    \I__5837\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30140\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30136\
        );

    \I__5835\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30133\
        );

    \I__5834\ : Span4Mux_v
    port map (
            O => \N__30136\,
            I => \N__30130\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__30133\,
            I => acadc_skipcnt_14
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__30130\,
            I => acadc_skipcnt_14
        );

    \I__5831\ : CascadeMux
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__5830\ : InMux
    port map (
            O => \N__30122\,
            I => \N__30118\
        );

    \I__5829\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30115\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30112\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__30115\,
            I => acadc_skipcnt_11
        );

    \I__5826\ : Odrv4
    port map (
            O => \N__30112\,
            I => acadc_skipcnt_11
        );

    \I__5825\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30102\
        );

    \I__5824\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30097\
        );

    \I__5823\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30097\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30094\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__30097\,
            I => \acadc_skipCount_11\
        );

    \I__5820\ : Odrv12
    port map (
            O => \N__30094\,
            I => \acadc_skipCount_11\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__30089\,
            I => \n23_adj_1199_cascade_\
        );

    \I__5818\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__30083\,
            I => n30
        );

    \I__5816\ : InMux
    port map (
            O => \N__30080\,
            I => \N__30077\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30073\
        );

    \I__5814\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30070\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__30073\,
            I => \N__30067\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__30070\,
            I => acadc_skipcnt_10
        );

    \I__5811\ : Odrv4
    port map (
            O => \N__30067\,
            I => acadc_skipcnt_10
        );

    \I__5810\ : InMux
    port map (
            O => \N__30062\,
            I => \N__30059\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__30059\,
            I => \N__30055\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__30058\,
            I => \N__30052\
        );

    \I__5807\ : Span4Mux_h
    port map (
            O => \N__30055\,
            I => \N__30049\
        );

    \I__5806\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30045\
        );

    \I__5805\ : Span4Mux_v
    port map (
            O => \N__30049\,
            I => \N__30042\
        );

    \I__5804\ : InMux
    port map (
            O => \N__30048\,
            I => \N__30039\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__30045\,
            I => \acadc_skipCount_12\
        );

    \I__5802\ : Odrv4
    port map (
            O => \N__30042\,
            I => \acadc_skipCount_12\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__30039\,
            I => \acadc_skipCount_12\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__5799\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30025\
        );

    \I__5798\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30022\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__30025\,
            I => \N__30019\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__30022\,
            I => acadc_skipcnt_12
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__30019\,
            I => acadc_skipcnt_12
        );

    \I__5794\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__30011\,
            I => n21
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \N__30005\
        );

    \I__5791\ : InMux
    port map (
            O => \N__30005\,
            I => \N__30000\
        );

    \I__5790\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29995\
        );

    \I__5789\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29995\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__30000\,
            I => \N__29992\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__29995\,
            I => data_index_0
        );

    \I__5786\ : Odrv4
    port map (
            O => \N__29992\,
            I => data_index_0
        );

    \I__5785\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__29981\,
            I => \data_index_9_N_647_0\
        );

    \I__5782\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29973\
        );

    \I__5781\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29970\
        );

    \I__5780\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29967\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__29973\,
            I => data_index_1
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__29970\,
            I => data_index_1
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__29967\,
            I => data_index_1
        );

    \I__5776\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29954\
        );

    \I__5775\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29954\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__29954\,
            I => n7_adj_1232
        );

    \I__5773\ : InMux
    port map (
            O => \N__29951\,
            I => n14031
        );

    \I__5772\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29943\
        );

    \I__5771\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29940\
        );

    \I__5770\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29937\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29932\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29932\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__29937\,
            I => data_index_2
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__29932\,
            I => data_index_2
        );

    \I__5765\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29921\
        );

    \I__5764\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29921\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__29921\,
            I => n7_adj_1230
        );

    \I__5762\ : InMux
    port map (
            O => \N__29918\,
            I => n14032
        );

    \I__5761\ : InMux
    port map (
            O => \N__29915\,
            I => n14033
        );

    \I__5760\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29908\
        );

    \I__5759\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29905\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__29908\,
            I => \N__29899\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__29905\,
            I => \N__29899\
        );

    \I__5756\ : InMux
    port map (
            O => \N__29904\,
            I => \N__29896\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__29899\,
            I => \N__29893\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__29896\,
            I => data_index_4
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__29893\,
            I => data_index_4
        );

    \I__5752\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29882\
        );

    \I__5751\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29882\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__29882\,
            I => \N__29879\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__29879\,
            I => n7_adj_1226
        );

    \I__5748\ : InMux
    port map (
            O => \N__29876\,
            I => n14034
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__29873\,
            I => \n7_adj_1177_cascade_\
        );

    \I__5746\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__29867\,
            I => n8_adj_1178
        );

    \I__5744\ : CascadeMux
    port map (
            O => \N__29864\,
            I => \N__29861\
        );

    \I__5743\ : CascadeBuf
    port map (
            O => \N__29861\,
            I => \N__29858\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__29858\,
            I => \N__29855\
        );

    \I__5741\ : CascadeBuf
    port map (
            O => \N__29855\,
            I => \N__29852\
        );

    \I__5740\ : CascadeMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__5739\ : CascadeBuf
    port map (
            O => \N__29849\,
            I => \N__29846\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__29846\,
            I => \N__29843\
        );

    \I__5737\ : CascadeBuf
    port map (
            O => \N__29843\,
            I => \N__29840\
        );

    \I__5736\ : CascadeMux
    port map (
            O => \N__29840\,
            I => \N__29837\
        );

    \I__5735\ : CascadeBuf
    port map (
            O => \N__29837\,
            I => \N__29834\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__29834\,
            I => \N__29831\
        );

    \I__5733\ : CascadeBuf
    port map (
            O => \N__29831\,
            I => \N__29828\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__5731\ : CascadeBuf
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__29822\,
            I => \N__29818\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__29821\,
            I => \N__29815\
        );

    \I__5728\ : CascadeBuf
    port map (
            O => \N__29818\,
            I => \N__29812\
        );

    \I__5727\ : CascadeBuf
    port map (
            O => \N__29815\,
            I => \N__29809\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__29812\,
            I => \N__29806\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__29809\,
            I => \N__29803\
        );

    \I__5724\ : CascadeBuf
    port map (
            O => \N__29806\,
            I => \N__29800\
        );

    \I__5723\ : InMux
    port map (
            O => \N__29803\,
            I => \N__29797\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__29800\,
            I => \N__29794\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__5720\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29788\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__29791\,
            I => \N__29785\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__29788\,
            I => \N__29782\
        );

    \I__5717\ : Span4Mux_v
    port map (
            O => \N__29785\,
            I => \N__29779\
        );

    \I__5716\ : Span4Mux_v
    port map (
            O => \N__29782\,
            I => \N__29776\
        );

    \I__5715\ : Span4Mux_h
    port map (
            O => \N__29779\,
            I => \N__29773\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__29776\,
            I => \N__29770\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__29773\,
            I => \N__29767\
        );

    \I__5712\ : Span4Mux_h
    port map (
            O => \N__29770\,
            I => \N__29764\
        );

    \I__5711\ : Odrv4
    port map (
            O => \N__29767\,
            I => \data_index_9_N_258_0\
        );

    \I__5710\ : Odrv4
    port map (
            O => \N__29764\,
            I => \data_index_9_N_258_0\
        );

    \I__5709\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29756\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__29756\,
            I => \N__29752\
        );

    \I__5707\ : InMux
    port map (
            O => \N__29755\,
            I => \N__29749\
        );

    \I__5706\ : Span4Mux_h
    port map (
            O => \N__29752\,
            I => \N__29746\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__29749\,
            I => acadc_skipcnt_0
        );

    \I__5704\ : Odrv4
    port map (
            O => \N__29746\,
            I => acadc_skipcnt_0
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__5702\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29734\
        );

    \I__5701\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29731\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__29734\,
            I => \N__29728\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__29731\,
            I => acadc_skipcnt_6
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__29728\,
            I => acadc_skipcnt_6
        );

    \I__5697\ : InMux
    port map (
            O => \N__29723\,
            I => \N__29720\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__29720\,
            I => \N__29717\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__29717\,
            I => n18_adj_1276
        );

    \I__5694\ : CascadeMux
    port map (
            O => \N__29714\,
            I => \n17_adj_1277_cascade_\
        );

    \I__5693\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29705\
        );

    \I__5692\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29705\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__29705\,
            I => n31
        );

    \I__5690\ : CascadeMux
    port map (
            O => \N__29702\,
            I => \n31_cascade_\
        );

    \I__5689\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29696\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__29696\,
            I => n15187
        );

    \I__5687\ : InMux
    port map (
            O => \N__29693\,
            I => \N__29687\
        );

    \I__5686\ : InMux
    port map (
            O => \N__29692\,
            I => \N__29687\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__29687\,
            I => n8_adj_1231
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__29684\,
            I => \N__29681\
        );

    \I__5683\ : CascadeBuf
    port map (
            O => \N__29681\,
            I => \N__29678\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__29678\,
            I => \N__29675\
        );

    \I__5681\ : CascadeBuf
    port map (
            O => \N__29675\,
            I => \N__29672\
        );

    \I__5680\ : CascadeMux
    port map (
            O => \N__29672\,
            I => \N__29669\
        );

    \I__5679\ : CascadeBuf
    port map (
            O => \N__29669\,
            I => \N__29666\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__29666\,
            I => \N__29663\
        );

    \I__5677\ : CascadeBuf
    port map (
            O => \N__29663\,
            I => \N__29660\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__29660\,
            I => \N__29657\
        );

    \I__5675\ : CascadeBuf
    port map (
            O => \N__29657\,
            I => \N__29654\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__29654\,
            I => \N__29651\
        );

    \I__5673\ : CascadeBuf
    port map (
            O => \N__29651\,
            I => \N__29648\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__29648\,
            I => \N__29645\
        );

    \I__5671\ : CascadeBuf
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__29642\,
            I => \N__29638\
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__29641\,
            I => \N__29635\
        );

    \I__5668\ : CascadeBuf
    port map (
            O => \N__29638\,
            I => \N__29632\
        );

    \I__5667\ : CascadeBuf
    port map (
            O => \N__29635\,
            I => \N__29629\
        );

    \I__5666\ : CascadeMux
    port map (
            O => \N__29632\,
            I => \N__29626\
        );

    \I__5665\ : CascadeMux
    port map (
            O => \N__29629\,
            I => \N__29623\
        );

    \I__5664\ : CascadeBuf
    port map (
            O => \N__29626\,
            I => \N__29620\
        );

    \I__5663\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29617\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__29620\,
            I => \N__29614\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__29617\,
            I => \N__29611\
        );

    \I__5660\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29608\
        );

    \I__5659\ : Span4Mux_h
    port map (
            O => \N__29611\,
            I => \N__29605\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29602\
        );

    \I__5657\ : Sp12to4
    port map (
            O => \N__29605\,
            I => \N__29599\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__29602\,
            I => \N__29596\
        );

    \I__5655\ : Span12Mux_v
    port map (
            O => \N__29599\,
            I => \N__29593\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__29596\,
            I => \N__29590\
        );

    \I__5653\ : Odrv12
    port map (
            O => \N__29593\,
            I => \data_index_9_N_258_2\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__29590\,
            I => \data_index_9_N_258_2\
        );

    \I__5651\ : IoInMux
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__29582\,
            I => \N__29578\
        );

    \I__5649\ : InMux
    port map (
            O => \N__29581\,
            I => \N__29575\
        );

    \I__5648\ : Span4Mux_s0_v
    port map (
            O => \N__29578\,
            I => \N__29572\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__29575\,
            I => \N__29569\
        );

    \I__5646\ : Span4Mux_v
    port map (
            O => \N__29572\,
            I => \N__29566\
        );

    \I__5645\ : Span4Mux_v
    port map (
            O => \N__29569\,
            I => \N__29562\
        );

    \I__5644\ : Span4Mux_v
    port map (
            O => \N__29566\,
            I => \N__29559\
        );

    \I__5643\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29556\
        );

    \I__5642\ : Span4Mux_h
    port map (
            O => \N__29562\,
            I => \N__29553\
        );

    \I__5641\ : Odrv4
    port map (
            O => \N__29559\,
            I => \M_FLT1\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__29556\,
            I => \M_FLT1\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__29553\,
            I => \M_FLT1\
        );

    \I__5638\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29541\
        );

    \I__5637\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29538\
        );

    \I__5636\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29535\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29532\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__29538\,
            I => \N__29529\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__29535\,
            I => buf_dds_14
        );

    \I__5632\ : Odrv12
    port map (
            O => \N__29532\,
            I => buf_dds_14
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__29529\,
            I => buf_dds_14
        );

    \I__5630\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__29516\,
            I => n4219
        );

    \I__5627\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29508\
        );

    \I__5626\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29505\
        );

    \I__5625\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29502\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__29508\,
            I => \N__29499\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29496\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__29502\,
            I => req_data_cnt_15
        );

    \I__5621\ : Odrv12
    port map (
            O => \N__29499\,
            I => req_data_cnt_15
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__29496\,
            I => req_data_cnt_15
        );

    \I__5619\ : InMux
    port map (
            O => \N__29489\,
            I => \N__29485\
        );

    \I__5618\ : InMux
    port map (
            O => \N__29488\,
            I => \N__29481\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__29485\,
            I => \N__29478\
        );

    \I__5616\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29475\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__29481\,
            I => req_data_cnt_9
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__29478\,
            I => req_data_cnt_9
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__29475\,
            I => req_data_cnt_9
        );

    \I__5612\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29465\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__29465\,
            I => n22
        );

    \I__5610\ : CascadeMux
    port map (
            O => \N__29462\,
            I => \n24_adj_1216_cascade_\
        );

    \I__5609\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29456\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__29456\,
            I => n30_adj_1278
        );

    \I__5607\ : CascadeMux
    port map (
            O => \N__29453\,
            I => \n6791_cascade_\
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__29450\,
            I => \n8_adj_1178_cascade_\
        );

    \I__5605\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29444\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__29444\,
            I => n7_adj_1177
        );

    \I__5603\ : IoInMux
    port map (
            O => \N__29441\,
            I => \N__29438\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__29438\,
            I => \N__29435\
        );

    \I__5601\ : Span4Mux_s2_v
    port map (
            O => \N__29435\,
            I => \N__29432\
        );

    \I__5600\ : Span4Mux_h
    port map (
            O => \N__29432\,
            I => \N__29429\
        );

    \I__5599\ : Sp12to4
    port map (
            O => \N__29429\,
            I => \N__29425\
        );

    \I__5598\ : InMux
    port map (
            O => \N__29428\,
            I => \N__29421\
        );

    \I__5597\ : Span12Mux_v
    port map (
            O => \N__29425\,
            I => \N__29418\
        );

    \I__5596\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29415\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__29421\,
            I => \N__29412\
        );

    \I__5594\ : Odrv12
    port map (
            O => \N__29418\,
            I => \M_OSR1\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__29415\,
            I => \M_OSR1\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__29412\,
            I => \M_OSR1\
        );

    \I__5591\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29402\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__29402\,
            I => \N__29399\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__29399\,
            I => n15479
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__29396\,
            I => \N__29393\
        );

    \I__5587\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29390\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29387\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__29387\,
            I => \N__29383\
        );

    \I__5584\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29380\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__29383\,
            I => cmd_rdadctmp_31_adj_1081
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__29380\,
            I => cmd_rdadctmp_31_adj_1081
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__29375\,
            I => \n8_adj_1221_cascade_\
        );

    \I__5580\ : CascadeMux
    port map (
            O => \N__29372\,
            I => \N__29369\
        );

    \I__5579\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29363\
        );

    \I__5577\ : Odrv4
    port map (
            O => \N__29363\,
            I => n4205
        );

    \I__5576\ : InMux
    port map (
            O => \N__29360\,
            I => \N__29357\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__29357\,
            I => \N__29353\
        );

    \I__5574\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29350\
        );

    \I__5573\ : Span4Mux_v
    port map (
            O => \N__29353\,
            I => \N__29347\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__29350\,
            I => buf_device_acadc_7
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__29347\,
            I => buf_device_acadc_7
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__29342\,
            I => \n4260_cascade_\
        );

    \I__5569\ : InMux
    port map (
            O => \N__29339\,
            I => \N__29336\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__29336\,
            I => \N__29333\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__29333\,
            I => \N__29330\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__29330\,
            I => n15402
        );

    \I__5565\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29324\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__29321\,
            I => \N__29318\
        );

    \I__5562\ : Span4Mux_v
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__5561\ : Span4Mux_v
    port map (
            O => \N__29315\,
            I => \N__29312\
        );

    \I__5560\ : Sp12to4
    port map (
            O => \N__29312\,
            I => \N__29309\
        );

    \I__5559\ : Span12Mux_h
    port map (
            O => \N__29309\,
            I => \N__29306\
        );

    \I__5558\ : Odrv12
    port map (
            O => \N__29306\,
            I => \ICE_CHKCABLE\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__29303\,
            I => \n90_adj_1154_cascade_\
        );

    \I__5556\ : InMux
    port map (
            O => \N__29300\,
            I => \N__29297\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__29297\,
            I => \N__29294\
        );

    \I__5554\ : Span4Mux_h
    port map (
            O => \N__29294\,
            I => \N__29291\
        );

    \I__5553\ : Span4Mux_h
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__29288\,
            I => n72
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__29285\,
            I => \N__29282\
        );

    \I__5550\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29279\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__29279\,
            I => \CLOCK_DDS.tmp_buf_10\
        );

    \I__5548\ : InMux
    port map (
            O => \N__29276\,
            I => \N__29273\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__29273\,
            I => \CLOCK_DDS.tmp_buf_11\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__29270\,
            I => \N__29267\
        );

    \I__5545\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29264\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29261\
        );

    \I__5543\ : Odrv4
    port map (
            O => \N__29261\,
            I => \CLOCK_DDS.tmp_buf_12\
        );

    \I__5542\ : CascadeMux
    port map (
            O => \N__29258\,
            I => \N__29255\
        );

    \I__5541\ : InMux
    port map (
            O => \N__29255\,
            I => \N__29252\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__29252\,
            I => \CLOCK_DDS.tmp_buf_13\
        );

    \I__5539\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29246\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__29246\,
            I => \CLOCK_DDS.tmp_buf_14\
        );

    \I__5537\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29240\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__29240\,
            I => \N__29236\
        );

    \I__5535\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29233\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__29236\,
            I => \N__29228\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29228\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__29228\,
            I => \N__29224\
        );

    \I__5531\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29221\
        );

    \I__5530\ : Sp12to4
    port map (
            O => \N__29224\,
            I => \N__29218\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__29221\,
            I => buf_dds_9
        );

    \I__5528\ : Odrv12
    port map (
            O => \N__29218\,
            I => buf_dds_9
        );

    \I__5527\ : CascadeMux
    port map (
            O => \N__29213\,
            I => \N__29210\
        );

    \I__5526\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29207\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__29207\,
            I => \CLOCK_DDS.tmp_buf_9\
        );

    \I__5524\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29201\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__29201\,
            I => \CLOCK_DDS.tmp_buf_8\
        );

    \I__5522\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29195\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29192\
        );

    \I__5520\ : Span4Mux_h
    port map (
            O => \N__29192\,
            I => \N__29189\
        );

    \I__5519\ : Span4Mux_v
    port map (
            O => \N__29189\,
            I => \N__29186\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__29186\,
            I => n15474
        );

    \I__5517\ : InMux
    port map (
            O => \N__29183\,
            I => \N__29180\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__29180\,
            I => \N__29177\
        );

    \I__5515\ : Span4Mux_h
    port map (
            O => \N__29177\,
            I => \N__29174\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__29174\,
            I => \N__29171\
        );

    \I__5513\ : Odrv4
    port map (
            O => \N__29171\,
            I => n15478
        );

    \I__5512\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29165\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__29165\,
            I => \N__29162\
        );

    \I__5510\ : Span4Mux_v
    port map (
            O => \N__29162\,
            I => \N__29159\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__29159\,
            I => n15680
        );

    \I__5508\ : InMux
    port map (
            O => \N__29156\,
            I => \N__29153\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29149\
        );

    \I__5506\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29146\
        );

    \I__5505\ : Span12Mux_v
    port map (
            O => \N__29149\,
            I => \N__29143\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29140\
        );

    \I__5503\ : Odrv12
    port map (
            O => \N__29143\,
            I => \comm_spi.n10449\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__29140\,
            I => \comm_spi.n10449\
        );

    \I__5501\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29132\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__29132\,
            I => \N__29129\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__29129\,
            I => \N__29125\
        );

    \I__5498\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29122\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__29125\,
            I => \comm_spi.n10448\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__29122\,
            I => \comm_spi.n10448\
        );

    \I__5495\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29114\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29111\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__29111\,
            I => \N__29108\
        );

    \I__5492\ : Span4Mux_h
    port map (
            O => \N__29108\,
            I => \N__29105\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__29105\,
            I => n15387
        );

    \I__5490\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29099\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__29099\,
            I => \N__29096\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__29096\,
            I => \N__29093\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__29093\,
            I => \N__29090\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__29090\,
            I => n15390
        );

    \I__5485\ : InMux
    port map (
            O => \N__29087\,
            I => \N__29084\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__29084\,
            I => \N__29081\
        );

    \I__5483\ : Odrv12
    port map (
            O => \N__29081\,
            I => buf_data2_22
        );

    \I__5482\ : InMux
    port map (
            O => \N__29078\,
            I => \N__29075\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29071\
        );

    \I__5480\ : CascadeMux
    port map (
            O => \N__29074\,
            I => \N__29068\
        );

    \I__5479\ : Span4Mux_h
    port map (
            O => \N__29071\,
            I => \N__29065\
        );

    \I__5478\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29062\
        );

    \I__5477\ : Span4Mux_h
    port map (
            O => \N__29065\,
            I => \N__29056\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__29062\,
            I => \N__29056\
        );

    \I__5475\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29053\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__29056\,
            I => \N__29050\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__29053\,
            I => buf_adcdata4_22
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__29050\,
            I => buf_adcdata4_22
        );

    \I__5471\ : InMux
    port map (
            O => \N__29045\,
            I => \N__29042\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__29042\,
            I => \N__29039\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__29036\,
            I => \N__29033\
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__29033\,
            I => n4102
        );

    \I__5466\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29025\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29022\
        );

    \I__5464\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29019\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__29025\,
            I => \comm_spi.n16902\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__29022\,
            I => \comm_spi.n16902\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__29019\,
            I => \comm_spi.n16902\
        );

    \I__5460\ : InMux
    port map (
            O => \N__29012\,
            I => \N__29009\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__29006\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__29006\,
            I => \N__29002\
        );

    \I__5457\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28999\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__29002\,
            I => \comm_spi.n10476\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__28999\,
            I => \comm_spi.n10476\
        );

    \I__5454\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28991\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28988\
        );

    \I__5452\ : Span4Mux_v
    port map (
            O => \N__28988\,
            I => \N__28985\
        );

    \I__5451\ : Span4Mux_h
    port map (
            O => \N__28985\,
            I => \N__28981\
        );

    \I__5450\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28978\
        );

    \I__5449\ : Odrv4
    port map (
            O => \N__28981\,
            I => \comm_spi.n10480\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__28978\,
            I => \comm_spi.n10480\
        );

    \I__5447\ : SRMux
    port map (
            O => \N__28973\,
            I => \N__28970\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__28970\,
            I => \comm_spi.data_tx_7__N_816\
        );

    \I__5445\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28964\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__28964\,
            I => \N__28960\
        );

    \I__5443\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28957\
        );

    \I__5442\ : Span4Mux_v
    port map (
            O => \N__28960\,
            I => \N__28954\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__28957\,
            I => \comm_spi.n10472\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__28954\,
            I => \comm_spi.n10472\
        );

    \I__5439\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28946\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__28946\,
            I => \N__28942\
        );

    \I__5437\ : InMux
    port map (
            O => \N__28945\,
            I => \N__28939\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__28942\,
            I => \comm_spi.n10471\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__28939\,
            I => \comm_spi.n10471\
        );

    \I__5434\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28931\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28928\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__28928\,
            I => \N__28924\
        );

    \I__5431\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28921\
        );

    \I__5430\ : Odrv4
    port map (
            O => \N__28924\,
            I => \comm_spi.n10475\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__28921\,
            I => \comm_spi.n10475\
        );

    \I__5428\ : SRMux
    port map (
            O => \N__28916\,
            I => \N__28913\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__28913\,
            I => \N__28910\
        );

    \I__5426\ : Odrv4
    port map (
            O => \N__28910\,
            I => \comm_spi.data_tx_7__N_807\
        );

    \I__5425\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28904\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__28904\,
            I => \N__28901\
        );

    \I__5423\ : Span4Mux_v
    port map (
            O => \N__28901\,
            I => \N__28898\
        );

    \I__5422\ : Span4Mux_h
    port map (
            O => \N__28898\,
            I => \N__28893\
        );

    \I__5421\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28890\
        );

    \I__5420\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28887\
        );

    \I__5419\ : Odrv4
    port map (
            O => \N__28893\,
            I => \comm_spi.n16896\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__28890\,
            I => \comm_spi.n16896\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__28887\,
            I => \comm_spi.n16896\
        );

    \I__5416\ : InMux
    port map (
            O => \N__28880\,
            I => n13972
        );

    \I__5415\ : InMux
    port map (
            O => \N__28877\,
            I => n13973
        );

    \I__5414\ : InMux
    port map (
            O => \N__28874\,
            I => \bfn_13_18_0_\
        );

    \I__5413\ : InMux
    port map (
            O => \N__28871\,
            I => n13975
        );

    \I__5412\ : InMux
    port map (
            O => \N__28868\,
            I => n13976
        );

    \I__5411\ : InMux
    port map (
            O => \N__28865\,
            I => n13977
        );

    \I__5410\ : InMux
    port map (
            O => \N__28862\,
            I => n13978
        );

    \I__5409\ : InMux
    port map (
            O => \N__28859\,
            I => n13979
        );

    \I__5408\ : InMux
    port map (
            O => \N__28856\,
            I => n13980
        );

    \I__5407\ : SRMux
    port map (
            O => \N__28853\,
            I => \N__28850\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__28850\,
            I => \N__28845\
        );

    \I__5405\ : SRMux
    port map (
            O => \N__28849\,
            I => \N__28842\
        );

    \I__5404\ : SRMux
    port map (
            O => \N__28848\,
            I => \N__28839\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__28845\,
            I => \N__28830\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__28842\,
            I => \N__28830\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__28839\,
            I => \N__28830\
        );

    \I__5400\ : SRMux
    port map (
            O => \N__28838\,
            I => \N__28827\
        );

    \I__5399\ : SRMux
    port map (
            O => \N__28837\,
            I => \N__28824\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__28830\,
            I => \N__28814\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__28827\,
            I => \N__28814\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28814\
        );

    \I__5395\ : SRMux
    port map (
            O => \N__28823\,
            I => \N__28811\
        );

    \I__5394\ : SRMux
    port map (
            O => \N__28822\,
            I => \N__28808\
        );

    \I__5393\ : SRMux
    port map (
            O => \N__28821\,
            I => \N__28803\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__28814\,
            I => \N__28795\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__28811\,
            I => \N__28795\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28795\
        );

    \I__5389\ : SRMux
    port map (
            O => \N__28807\,
            I => \N__28792\
        );

    \I__5388\ : SRMux
    port map (
            O => \N__28806\,
            I => \N__28789\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28786\
        );

    \I__5386\ : SRMux
    port map (
            O => \N__28802\,
            I => \N__28783\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__28795\,
            I => \N__28775\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28775\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28775\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__28786\,
            I => \N__28762\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__28783\,
            I => \N__28762\
        );

    \I__5380\ : IoInMux
    port map (
            O => \N__28782\,
            I => \N__28759\
        );

    \I__5379\ : Span4Mux_v
    port map (
            O => \N__28775\,
            I => \N__28756\
        );

    \I__5378\ : SRMux
    port map (
            O => \N__28774\,
            I => \N__28753\
        );

    \I__5377\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28744\
        );

    \I__5376\ : InMux
    port map (
            O => \N__28772\,
            I => \N__28744\
        );

    \I__5375\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28744\
        );

    \I__5374\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28735\
        );

    \I__5373\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28735\
        );

    \I__5372\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28735\
        );

    \I__5371\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28735\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__28762\,
            I => \N__28732\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__28759\,
            I => \N__28729\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__28756\,
            I => \N__28724\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__28753\,
            I => \N__28724\
        );

    \I__5366\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28721\
        );

    \I__5365\ : InMux
    port map (
            O => \N__28751\,
            I => \N__28718\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__28744\,
            I => \N__28713\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__28735\,
            I => \N__28713\
        );

    \I__5362\ : Span4Mux_h
    port map (
            O => \N__28732\,
            I => \N__28710\
        );

    \I__5361\ : Span4Mux_s2_v
    port map (
            O => \N__28729\,
            I => \N__28707\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__28724\,
            I => \N__28704\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__28721\,
            I => \N__28699\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__28718\,
            I => \N__28699\
        );

    \I__5357\ : Span12Mux_v
    port map (
            O => \N__28713\,
            I => \N__28696\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__28710\,
            I => \N__28691\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__28707\,
            I => \N__28691\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__28704\,
            I => \N__28686\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__28699\,
            I => \N__28686\
        );

    \I__5352\ : Odrv12
    port map (
            O => \N__28696\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__28691\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5350\ : Odrv4
    port map (
            O => \N__28686\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5349\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28675\
        );

    \I__5348\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28672\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__28675\,
            I => \N__28669\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__28672\,
            I => acadc_skipcnt_1
        );

    \I__5345\ : Odrv4
    port map (
            O => \N__28669\,
            I => acadc_skipcnt_1
        );

    \I__5344\ : InMux
    port map (
            O => \N__28664\,
            I => \bfn_13_17_0_\
        );

    \I__5343\ : InMux
    port map (
            O => \N__28661\,
            I => n13967
        );

    \I__5342\ : InMux
    port map (
            O => \N__28658\,
            I => n13968
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__28655\,
            I => \N__28652\
        );

    \I__5340\ : InMux
    port map (
            O => \N__28652\,
            I => \N__28648\
        );

    \I__5339\ : InMux
    port map (
            O => \N__28651\,
            I => \N__28645\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__28648\,
            I => \N__28642\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__28645\,
            I => acadc_skipcnt_4
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__28642\,
            I => acadc_skipcnt_4
        );

    \I__5335\ : InMux
    port map (
            O => \N__28637\,
            I => n13969
        );

    \I__5334\ : InMux
    port map (
            O => \N__28634\,
            I => n13970
        );

    \I__5333\ : InMux
    port map (
            O => \N__28631\,
            I => n13971
        );

    \I__5332\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28625\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__28625\,
            I => \N__28622\
        );

    \I__5330\ : Span12Mux_h
    port map (
            O => \N__28622\,
            I => \N__28619\
        );

    \I__5329\ : Odrv12
    port map (
            O => \N__28619\,
            I => buf_data2_13
        );

    \I__5328\ : InMux
    port map (
            O => \N__28616\,
            I => \N__28611\
        );

    \I__5327\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28608\
        );

    \I__5326\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28605\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__28611\,
            I => \N__28598\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28598\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__28605\,
            I => \N__28598\
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__28598\,
            I => buf_adcdata4_13
        );

    \I__5321\ : InMux
    port map (
            O => \N__28595\,
            I => \N__28592\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__28592\,
            I => \N__28589\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__5318\ : Span4Mux_h
    port map (
            O => \N__28586\,
            I => \N__28583\
        );

    \I__5317\ : Span4Mux_h
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__28580\,
            I => n4059
        );

    \I__5315\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28574\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__28574\,
            I => n8_adj_1233
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__28571\,
            I => \n8_adj_1233_cascade_\
        );

    \I__5312\ : IoInMux
    port map (
            O => \N__28568\,
            I => \N__28565\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__28565\,
            I => \N__28562\
        );

    \I__5310\ : Span4Mux_s3_v
    port map (
            O => \N__28562\,
            I => \N__28559\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__28559\,
            I => \N__28555\
        );

    \I__5308\ : CascadeMux
    port map (
            O => \N__28558\,
            I => \N__28551\
        );

    \I__5307\ : Span4Mux_v
    port map (
            O => \N__28555\,
            I => \N__28548\
        );

    \I__5306\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28545\
        );

    \I__5305\ : InMux
    port map (
            O => \N__28551\,
            I => \N__28542\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__28548\,
            I => \M_FLT0\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__28545\,
            I => \M_FLT0\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__28542\,
            I => \M_FLT0\
        );

    \I__5301\ : InMux
    port map (
            O => \N__28535\,
            I => \N__28532\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__28532\,
            I => \N__28529\
        );

    \I__5299\ : Odrv12
    port map (
            O => \N__28529\,
            I => n66_adj_1166
        );

    \I__5298\ : InMux
    port map (
            O => \N__28526\,
            I => \bfn_13_16_0_\
        );

    \I__5297\ : InMux
    port map (
            O => \N__28523\,
            I => \N__28519\
        );

    \I__5296\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28516\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__28519\,
            I => \eis_end_N_773\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__28516\,
            I => \eis_end_N_773\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__28511\,
            I => \eis_end_N_773_cascade_\
        );

    \I__5292\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28505\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__28505\,
            I => n15510
        );

    \I__5290\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28496\
        );

    \I__5289\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28496\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__28496\,
            I => n8_adj_1227
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__28493\,
            I => \N__28490\
        );

    \I__5286\ : InMux
    port map (
            O => \N__28490\,
            I => \N__28484\
        );

    \I__5285\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28484\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28480\
        );

    \I__5283\ : CascadeMux
    port map (
            O => \N__28483\,
            I => \N__28477\
        );

    \I__5282\ : Span4Mux_h
    port map (
            O => \N__28480\,
            I => \N__28474\
        );

    \I__5281\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28471\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__28474\,
            I => cmd_rdadctmp_24_adj_1088
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__28471\,
            I => cmd_rdadctmp_24_adj_1088
        );

    \I__5278\ : CascadeMux
    port map (
            O => \N__28466\,
            I => \N__28463\
        );

    \I__5277\ : CascadeBuf
    port map (
            O => \N__28463\,
            I => \N__28460\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__28460\,
            I => \N__28457\
        );

    \I__5275\ : CascadeBuf
    port map (
            O => \N__28457\,
            I => \N__28454\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__28454\,
            I => \N__28451\
        );

    \I__5273\ : CascadeBuf
    port map (
            O => \N__28451\,
            I => \N__28448\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__28448\,
            I => \N__28445\
        );

    \I__5271\ : CascadeBuf
    port map (
            O => \N__28445\,
            I => \N__28442\
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__28442\,
            I => \N__28439\
        );

    \I__5269\ : CascadeBuf
    port map (
            O => \N__28439\,
            I => \N__28436\
        );

    \I__5268\ : CascadeMux
    port map (
            O => \N__28436\,
            I => \N__28433\
        );

    \I__5267\ : CascadeBuf
    port map (
            O => \N__28433\,
            I => \N__28430\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__5265\ : CascadeBuf
    port map (
            O => \N__28427\,
            I => \N__28423\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__28426\,
            I => \N__28420\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__28423\,
            I => \N__28417\
        );

    \I__5262\ : CascadeBuf
    port map (
            O => \N__28420\,
            I => \N__28414\
        );

    \I__5261\ : CascadeBuf
    port map (
            O => \N__28417\,
            I => \N__28411\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__28414\,
            I => \N__28408\
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__28411\,
            I => \N__28405\
        );

    \I__5258\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28402\
        );

    \I__5257\ : CascadeBuf
    port map (
            O => \N__28405\,
            I => \N__28399\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__28402\,
            I => \N__28396\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__28399\,
            I => \N__28393\
        );

    \I__5254\ : Span4Mux_h
    port map (
            O => \N__28396\,
            I => \N__28390\
        );

    \I__5253\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28387\
        );

    \I__5252\ : Span4Mux_v
    port map (
            O => \N__28390\,
            I => \N__28384\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__28387\,
            I => \N__28381\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__5249\ : Span4Mux_v
    port map (
            O => \N__28381\,
            I => \N__28375\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__28378\,
            I => \N__28372\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__28375\,
            I => \N__28369\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__28372\,
            I => \data_index_9_N_258_1\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__28369\,
            I => \data_index_9_N_258_1\
        );

    \I__5244\ : SRMux
    port map (
            O => \N__28364\,
            I => \N__28360\
        );

    \I__5243\ : SRMux
    port map (
            O => \N__28363\,
            I => \N__28355\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__28360\,
            I => \N__28350\
        );

    \I__5241\ : SRMux
    port map (
            O => \N__28359\,
            I => \N__28347\
        );

    \I__5240\ : SRMux
    port map (
            O => \N__28358\,
            I => \N__28341\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__28355\,
            I => \N__28337\
        );

    \I__5238\ : SRMux
    port map (
            O => \N__28354\,
            I => \N__28334\
        );

    \I__5237\ : SRMux
    port map (
            O => \N__28353\,
            I => \N__28331\
        );

    \I__5236\ : Span4Mux_v
    port map (
            O => \N__28350\,
            I => \N__28326\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__28347\,
            I => \N__28326\
        );

    \I__5234\ : SRMux
    port map (
            O => \N__28346\,
            I => \N__28323\
        );

    \I__5233\ : SRMux
    port map (
            O => \N__28345\,
            I => \N__28319\
        );

    \I__5232\ : SRMux
    port map (
            O => \N__28344\,
            I => \N__28316\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28313\
        );

    \I__5230\ : SRMux
    port map (
            O => \N__28340\,
            I => \N__28310\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__28337\,
            I => \N__28305\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28305\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__28331\,
            I => \N__28302\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__28326\,
            I => \N__28297\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__28323\,
            I => \N__28297\
        );

    \I__5224\ : SRMux
    port map (
            O => \N__28322\,
            I => \N__28294\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__28319\,
            I => \N__28291\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__28316\,
            I => \N__28288\
        );

    \I__5221\ : Span4Mux_h
    port map (
            O => \N__28313\,
            I => \N__28285\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__28310\,
            I => \N__28282\
        );

    \I__5219\ : Span4Mux_v
    port map (
            O => \N__28305\,
            I => \N__28273\
        );

    \I__5218\ : Span4Mux_h
    port map (
            O => \N__28302\,
            I => \N__28273\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__28297\,
            I => \N__28273\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__28294\,
            I => \N__28273\
        );

    \I__5215\ : Span4Mux_v
    port map (
            O => \N__28291\,
            I => \N__28269\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__28288\,
            I => \N__28266\
        );

    \I__5213\ : Span4Mux_v
    port map (
            O => \N__28285\,
            I => \N__28261\
        );

    \I__5212\ : Span4Mux_h
    port map (
            O => \N__28282\,
            I => \N__28261\
        );

    \I__5211\ : Span4Mux_v
    port map (
            O => \N__28273\,
            I => \N__28258\
        );

    \I__5210\ : SRMux
    port map (
            O => \N__28272\,
            I => \N__28255\
        );

    \I__5209\ : Span4Mux_h
    port map (
            O => \N__28269\,
            I => \N__28252\
        );

    \I__5208\ : Span4Mux_v
    port map (
            O => \N__28266\,
            I => \N__28249\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__28261\,
            I => \N__28242\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__28258\,
            I => \N__28242\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__28255\,
            I => \N__28242\
        );

    \I__5204\ : Span4Mux_h
    port map (
            O => \N__28252\,
            I => \N__28239\
        );

    \I__5203\ : Span4Mux_h
    port map (
            O => \N__28249\,
            I => \N__28236\
        );

    \I__5202\ : Sp12to4
    port map (
            O => \N__28242\,
            I => \N__28233\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__28239\,
            I => \raw_buf1_N_775\
        );

    \I__5200\ : Odrv4
    port map (
            O => \N__28236\,
            I => \raw_buf1_N_775\
        );

    \I__5199\ : Odrv12
    port map (
            O => \N__28233\,
            I => \raw_buf1_N_775\
        );

    \I__5198\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28222\
        );

    \I__5197\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28219\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__28222\,
            I => \N__28214\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28214\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__28214\,
            I => \N__28211\
        );

    \I__5193\ : Odrv4
    port map (
            O => \N__28211\,
            I => n14087
        );

    \I__5192\ : CascadeMux
    port map (
            O => \N__28208\,
            I => \n15356_cascade_\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__28205\,
            I => \n15695_cascade_\
        );

    \I__5190\ : InMux
    port map (
            O => \N__28202\,
            I => \N__28199\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__28199\,
            I => n15696
        );

    \I__5188\ : CascadeMux
    port map (
            O => \N__28196\,
            I => \n15700_cascade_\
        );

    \I__5187\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28190\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__28190\,
            I => n3
        );

    \I__5185\ : CEMux
    port map (
            O => \N__28187\,
            I => \N__28184\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__28184\,
            I => n8459
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__28181\,
            I => \N__28178\
        );

    \I__5182\ : CascadeBuf
    port map (
            O => \N__28178\,
            I => \N__28175\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__28175\,
            I => \N__28172\
        );

    \I__5180\ : CascadeBuf
    port map (
            O => \N__28172\,
            I => \N__28169\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__28169\,
            I => \N__28166\
        );

    \I__5178\ : CascadeBuf
    port map (
            O => \N__28166\,
            I => \N__28163\
        );

    \I__5177\ : CascadeMux
    port map (
            O => \N__28163\,
            I => \N__28160\
        );

    \I__5176\ : CascadeBuf
    port map (
            O => \N__28160\,
            I => \N__28157\
        );

    \I__5175\ : CascadeMux
    port map (
            O => \N__28157\,
            I => \N__28154\
        );

    \I__5174\ : CascadeBuf
    port map (
            O => \N__28154\,
            I => \N__28151\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__28151\,
            I => \N__28148\
        );

    \I__5172\ : CascadeBuf
    port map (
            O => \N__28148\,
            I => \N__28145\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__28145\,
            I => \N__28142\
        );

    \I__5170\ : CascadeBuf
    port map (
            O => \N__28142\,
            I => \N__28138\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__28141\,
            I => \N__28135\
        );

    \I__5168\ : CascadeMux
    port map (
            O => \N__28138\,
            I => \N__28132\
        );

    \I__5167\ : CascadeBuf
    port map (
            O => \N__28135\,
            I => \N__28129\
        );

    \I__5166\ : CascadeBuf
    port map (
            O => \N__28132\,
            I => \N__28126\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__28129\,
            I => \N__28123\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__5163\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28117\
        );

    \I__5162\ : CascadeBuf
    port map (
            O => \N__28120\,
            I => \N__28114\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__28117\,
            I => \N__28111\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__28114\,
            I => \N__28108\
        );

    \I__5159\ : Span4Mux_v
    port map (
            O => \N__28111\,
            I => \N__28105\
        );

    \I__5158\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28102\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__28105\,
            I => \N__28099\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28096\
        );

    \I__5155\ : Span4Mux_h
    port map (
            O => \N__28099\,
            I => \N__28093\
        );

    \I__5154\ : Span12Mux_v
    port map (
            O => \N__28096\,
            I => \N__28090\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__28093\,
            I => \data_index_9_N_258_4\
        );

    \I__5152\ : Odrv12
    port map (
            O => \N__28090\,
            I => \data_index_9_N_258_4\
        );

    \I__5151\ : IoInMux
    port map (
            O => \N__28085\,
            I => \N__28082\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__28082\,
            I => \N__28079\
        );

    \I__5149\ : IoSpan4Mux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__5148\ : Span4Mux_s3_v
    port map (
            O => \N__28076\,
            I => \N__28073\
        );

    \I__5147\ : Sp12to4
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__5146\ : Span12Mux_s10_v
    port map (
            O => \N__28070\,
            I => \N__28067\
        );

    \I__5145\ : Span12Mux_h
    port map (
            O => \N__28067\,
            I => \N__28062\
        );

    \I__5144\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28057\
        );

    \I__5143\ : InMux
    port map (
            O => \N__28065\,
            I => \N__28057\
        );

    \I__5142\ : Odrv12
    port map (
            O => \N__28062\,
            I => \M_OSR0\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__28057\,
            I => \M_OSR0\
        );

    \I__5140\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28049\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__28049\,
            I => \N__28046\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__28046\,
            I => \N__28043\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__28043\,
            I => n15555
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__28040\,
            I => \n3_cascade_\
        );

    \I__5135\ : CascadeMux
    port map (
            O => \N__28037\,
            I => \n10_adj_1242_cascade_\
        );

    \I__5134\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28031\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__28031\,
            I => n8_adj_1212
        );

    \I__5132\ : InMux
    port map (
            O => \N__28028\,
            I => \N__28024\
        );

    \I__5131\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28021\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__28024\,
            I => eis_end
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__28021\,
            I => eis_end
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__28016\,
            I => \n15171_cascade_\
        );

    \I__5127\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28010\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__28007\,
            I => n15475
        );

    \I__5124\ : CascadeMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__5123\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27998\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__27998\,
            I => n15835
        );

    \I__5121\ : InMux
    port map (
            O => \N__27995\,
            I => \N__27992\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__27992\,
            I => \N__27989\
        );

    \I__5119\ : Span4Mux_h
    port map (
            O => \N__27989\,
            I => \N__27986\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__27986\,
            I => \N__27983\
        );

    \I__5117\ : Odrv4
    port map (
            O => \N__27983\,
            I => n15542
        );

    \I__5116\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27977\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__27977\,
            I => \N__27974\
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__27974\,
            I => n15679
        );

    \I__5113\ : InMux
    port map (
            O => \N__27971\,
            I => \N__27968\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27965\
        );

    \I__5111\ : Span4Mux_v
    port map (
            O => \N__27965\,
            I => \N__27962\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__27962\,
            I => n15543
        );

    \I__5109\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27956\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__27956\,
            I => \N__27951\
        );

    \I__5107\ : InMux
    port map (
            O => \N__27955\,
            I => \N__27948\
        );

    \I__5106\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27945\
        );

    \I__5105\ : Span12Mux_s11_h
    port map (
            O => \N__27951\,
            I => \N__27942\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__27948\,
            I => \N__27939\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__27945\,
            I => buf_adcdata3_17
        );

    \I__5102\ : Odrv12
    port map (
            O => \N__27942\,
            I => buf_adcdata3_17
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__27939\,
            I => buf_adcdata3_17
        );

    \I__5100\ : IoInMux
    port map (
            O => \N__27932\,
            I => \N__27929\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__27929\,
            I => \N__27926\
        );

    \I__5098\ : IoSpan4Mux
    port map (
            O => \N__27926\,
            I => \N__27922\
        );

    \I__5097\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27919\
        );

    \I__5096\ : Sp12to4
    port map (
            O => \N__27922\,
            I => \N__27916\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__27919\,
            I => \N__27912\
        );

    \I__5094\ : Span12Mux_v
    port map (
            O => \N__27916\,
            I => \N__27909\
        );

    \I__5093\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27906\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__27912\,
            I => \N__27903\
        );

    \I__5091\ : Odrv12
    port map (
            O => \N__27909\,
            I => \M_DCSEL\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__27906\,
            I => \M_DCSEL\
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__27903\,
            I => \M_DCSEL\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__27896\,
            I => \n90_adj_1023_cascade_\
        );

    \I__5087\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27890\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__27890\,
            I => n69_adj_1113
        );

    \I__5085\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27884\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27881\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__27881\,
            I => n96
        );

    \I__5082\ : InMux
    port map (
            O => \N__27878\,
            I => \N__27874\
        );

    \I__5081\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27871\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__27874\,
            I => buf_device_acadc_4
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__27871\,
            I => buf_device_acadc_4
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__27866\,
            I => \n4814_cascade_\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__27863\,
            I => \N__27857\
        );

    \I__5076\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27851\
        );

    \I__5075\ : InMux
    port map (
            O => \N__27861\,
            I => \N__27851\
        );

    \I__5074\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27848\
        );

    \I__5073\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27845\
        );

    \I__5072\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27842\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__27851\,
            I => n5_adj_1235
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__27848\,
            I => n5_adj_1235
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__27845\,
            I => n5_adj_1235
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__27842\,
            I => n5_adj_1235
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__27833\,
            I => \n13475_cascade_\
        );

    \I__5066\ : CascadeMux
    port map (
            O => \N__27830\,
            I => \n15802_cascade_\
        );

    \I__5065\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27824\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__27824\,
            I => \N__27821\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__27818\,
            I => \N__27815\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__27815\,
            I => n10_adj_1249
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__27812\,
            I => \n15657_cascade_\
        );

    \I__5059\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27806\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__5057\ : Span4Mux_h
    port map (
            O => \N__27803\,
            I => \N__27800\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__27800\,
            I => \N__27797\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__27797\,
            I => n13_adj_1042
        );

    \I__5054\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27791\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__27791\,
            I => \N__27788\
        );

    \I__5052\ : Span4Mux_h
    port map (
            O => \N__27788\,
            I => \N__27784\
        );

    \I__5051\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27781\
        );

    \I__5050\ : Span4Mux_h
    port map (
            O => \N__27784\,
            I => \N__27778\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27775\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__27778\,
            I => \comm_spi.n10479\
        );

    \I__5047\ : Odrv12
    port map (
            O => \N__27775\,
            I => \comm_spi.n10479\
        );

    \I__5046\ : SRMux
    port map (
            O => \N__27770\,
            I => \N__27767\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27764\
        );

    \I__5044\ : Span4Mux_v
    port map (
            O => \N__27764\,
            I => \N__27761\
        );

    \I__5043\ : Odrv4
    port map (
            O => \N__27761\,
            I => \comm_spi.data_tx_7__N_806\
        );

    \I__5042\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27752\
        );

    \I__5040\ : Odrv12
    port map (
            O => \N__27752\,
            I => n15576
        );

    \I__5039\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27746\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__27746\,
            I => \N__27743\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__27743\,
            I => \N__27740\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__27740\,
            I => n15691
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__27737\,
            I => \n15567_cascade_\
        );

    \I__5034\ : InMux
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__27731\,
            I => \N__27728\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__27728\,
            I => \N__27725\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__27725\,
            I => n7_adj_1255
        );

    \I__5030\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27719\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__27719\,
            I => n6
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__27716\,
            I => \n5_adj_1235_cascade_\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__27713\,
            I => \n15535_cascade_\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__27710\,
            I => \n15_cascade_\
        );

    \I__5025\ : CEMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27701\
        );

    \I__5023\ : Span4Mux_h
    port map (
            O => \N__27701\,
            I => \N__27698\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__27698\,
            I => n9021
        );

    \I__5021\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27692\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__27692\,
            I => n4814
        );

    \I__5019\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27680\
        );

    \I__5018\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27680\
        );

    \I__5017\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27680\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__27680\,
            I => \N__27677\
        );

    \I__5015\ : Span4Mux_h
    port map (
            O => \N__27677\,
            I => \N__27674\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__27674\,
            I => \N__27671\
        );

    \I__5013\ : Odrv4
    port map (
            O => \N__27671\,
            I => comm_tx_buf_6
        );

    \I__5012\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27665\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__27662\,
            I => \N__27659\
        );

    \I__5009\ : Span4Mux_h
    port map (
            O => \N__27659\,
            I => \N__27654\
        );

    \I__5008\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27651\
        );

    \I__5007\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27648\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__27654\,
            I => \comm_spi.n16884\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__27651\,
            I => \comm_spi.n16884\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__27648\,
            I => \comm_spi.n16884\
        );

    \I__5003\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27638\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__27638\,
            I => \N__27635\
        );

    \I__5001\ : Span4Mux_v
    port map (
            O => \N__27635\,
            I => \N__27632\
        );

    \I__5000\ : Span4Mux_h
    port map (
            O => \N__27632\,
            I => \N__27629\
        );

    \I__4999\ : Span4Mux_h
    port map (
            O => \N__27629\,
            I => \N__27626\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__27626\,
            I => buf_data1_23
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__27623\,
            I => \n18_cascade_\
        );

    \I__4996\ : CascadeMux
    port map (
            O => \N__27620\,
            I => \n15466_cascade_\
        );

    \I__4995\ : CascadeMux
    port map (
            O => \N__27617\,
            I => \N__27614\
        );

    \I__4994\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27611\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__4992\ : Span4Mux_h
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__27605\,
            I => \N__27602\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__27602\,
            I => n104
        );

    \I__4989\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27596\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__27596\,
            I => n56
        );

    \I__4987\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27590\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__27590\,
            I => \N__27587\
        );

    \I__4985\ : Span4Mux_h
    port map (
            O => \N__27587\,
            I => \N__27583\
        );

    \I__4984\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27580\
        );

    \I__4983\ : Span4Mux_h
    port map (
            O => \N__27583\,
            I => \N__27575\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__27580\,
            I => \N__27575\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__27575\,
            I => \N__27572\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__27572\,
            I => \N__27568\
        );

    \I__4979\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27565\
        );

    \I__4978\ : Span4Mux_h
    port map (
            O => \N__27568\,
            I => \N__27562\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__27565\,
            I => buf_adcdata3_1
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__27562\,
            I => buf_adcdata3_1
        );

    \I__4975\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27554\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__27554\,
            I => \N__27551\
        );

    \I__4973\ : Span12Mux_h
    port map (
            O => \N__27551\,
            I => \N__27548\
        );

    \I__4972\ : Odrv12
    port map (
            O => \N__27548\,
            I => buf_data1_1
        );

    \I__4971\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__27542\,
            I => \N__27539\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__27536\,
            I => \N__27533\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__27533\,
            I => n4151
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__27530\,
            I => \N__27521\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__27529\,
            I => \N__27518\
        );

    \I__4964\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27506\
        );

    \I__4963\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27506\
        );

    \I__4962\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27503\
        );

    \I__4961\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27490\
        );

    \I__4960\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27490\
        );

    \I__4959\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27490\
        );

    \I__4958\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27490\
        );

    \I__4957\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27490\
        );

    \I__4956\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27490\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__27515\,
            I => \N__27486\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__27514\,
            I => \N__27479\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__27513\,
            I => \N__27476\
        );

    \I__4952\ : CascadeMux
    port map (
            O => \N__27512\,
            I => \N__27473\
        );

    \I__4951\ : InMux
    port map (
            O => \N__27511\,
            I => \N__27461\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27454\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__27503\,
            I => \N__27454\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27444\
        );

    \I__4947\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27441\
        );

    \I__4946\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27438\
        );

    \I__4945\ : InMux
    port map (
            O => \N__27485\,
            I => \N__27429\
        );

    \I__4944\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27429\
        );

    \I__4943\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27429\
        );

    \I__4942\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27429\
        );

    \I__4941\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27416\
        );

    \I__4940\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27416\
        );

    \I__4939\ : InMux
    port map (
            O => \N__27473\,
            I => \N__27416\
        );

    \I__4938\ : InMux
    port map (
            O => \N__27472\,
            I => \N__27416\
        );

    \I__4937\ : InMux
    port map (
            O => \N__27471\,
            I => \N__27416\
        );

    \I__4936\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27416\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__27469\,
            I => \N__27412\
        );

    \I__4934\ : InMux
    port map (
            O => \N__27468\,
            I => \N__27407\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__27467\,
            I => \N__27404\
        );

    \I__4932\ : InMux
    port map (
            O => \N__27466\,
            I => \N__27400\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__27465\,
            I => \N__27395\
        );

    \I__4930\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27390\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27387\
        );

    \I__4928\ : InMux
    port map (
            O => \N__27460\,
            I => \N__27384\
        );

    \I__4927\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27381\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__27454\,
            I => \N__27369\
        );

    \I__4925\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27354\
        );

    \I__4924\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27354\
        );

    \I__4923\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27354\
        );

    \I__4922\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27354\
        );

    \I__4921\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27354\
        );

    \I__4920\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27354\
        );

    \I__4919\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27354\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__27444\,
            I => \N__27347\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__27441\,
            I => \N__27347\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__27438\,
            I => \N__27340\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__27429\,
            I => \N__27340\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__27416\,
            I => \N__27340\
        );

    \I__4913\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27337\
        );

    \I__4912\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27329\
        );

    \I__4911\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27329\
        );

    \I__4910\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27329\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__27407\,
            I => \N__27326\
        );

    \I__4908\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27323\
        );

    \I__4907\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27319\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27316\
        );

    \I__4905\ : InMux
    port map (
            O => \N__27399\,
            I => \N__27305\
        );

    \I__4904\ : InMux
    port map (
            O => \N__27398\,
            I => \N__27305\
        );

    \I__4903\ : InMux
    port map (
            O => \N__27395\,
            I => \N__27305\
        );

    \I__4902\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27305\
        );

    \I__4901\ : InMux
    port map (
            O => \N__27393\,
            I => \N__27305\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__27390\,
            I => \N__27302\
        );

    \I__4899\ : Span4Mux_v
    port map (
            O => \N__27387\,
            I => \N__27299\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__27384\,
            I => \N__27294\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__27381\,
            I => \N__27294\
        );

    \I__4896\ : InMux
    port map (
            O => \N__27380\,
            I => \N__27289\
        );

    \I__4895\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27289\
        );

    \I__4894\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27273\
        );

    \I__4893\ : InMux
    port map (
            O => \N__27377\,
            I => \N__27273\
        );

    \I__4892\ : InMux
    port map (
            O => \N__27376\,
            I => \N__27273\
        );

    \I__4891\ : InMux
    port map (
            O => \N__27375\,
            I => \N__27273\
        );

    \I__4890\ : InMux
    port map (
            O => \N__27374\,
            I => \N__27273\
        );

    \I__4889\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27273\
        );

    \I__4888\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27273\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__27369\,
            I => \N__27270\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__27354\,
            I => \N__27267\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27264\
        );

    \I__4884\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27261\
        );

    \I__4883\ : Span4Mux_h
    port map (
            O => \N__27347\,
            I => \N__27258\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__27340\,
            I => \N__27253\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__27337\,
            I => \N__27253\
        );

    \I__4880\ : InMux
    port map (
            O => \N__27336\,
            I => \N__27247\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__27329\,
            I => \N__27244\
        );

    \I__4878\ : Span4Mux_h
    port map (
            O => \N__27326\,
            I => \N__27239\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__27323\,
            I => \N__27239\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__27322\,
            I => \N__27231\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__27319\,
            I => \N__27222\
        );

    \I__4874\ : Span4Mux_h
    port map (
            O => \N__27316\,
            I => \N__27222\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__27305\,
            I => \N__27222\
        );

    \I__4872\ : Span4Mux_v
    port map (
            O => \N__27302\,
            I => \N__27215\
        );

    \I__4871\ : Span4Mux_v
    port map (
            O => \N__27299\,
            I => \N__27215\
        );

    \I__4870\ : Span4Mux_h
    port map (
            O => \N__27294\,
            I => \N__27215\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27212\
        );

    \I__4868\ : InMux
    port map (
            O => \N__27288\,
            I => \N__27209\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__27273\,
            I => \N__27202\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__27270\,
            I => \N__27202\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__27267\,
            I => \N__27202\
        );

    \I__4864\ : InMux
    port map (
            O => \N__27264\,
            I => \N__27199\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__27261\,
            I => \N__27194\
        );

    \I__4862\ : Sp12to4
    port map (
            O => \N__27258\,
            I => \N__27194\
        );

    \I__4861\ : Sp12to4
    port map (
            O => \N__27253\,
            I => \N__27191\
        );

    \I__4860\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27188\
        );

    \I__4859\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27183\
        );

    \I__4858\ : InMux
    port map (
            O => \N__27250\,
            I => \N__27183\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__27247\,
            I => \N__27180\
        );

    \I__4856\ : Span4Mux_v
    port map (
            O => \N__27244\,
            I => \N__27175\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__27239\,
            I => \N__27175\
        );

    \I__4854\ : InMux
    port map (
            O => \N__27238\,
            I => \N__27172\
        );

    \I__4853\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27161\
        );

    \I__4852\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27161\
        );

    \I__4851\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27161\
        );

    \I__4850\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27161\
        );

    \I__4849\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27161\
        );

    \I__4848\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27156\
        );

    \I__4847\ : InMux
    port map (
            O => \N__27229\,
            I => \N__27156\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__27222\,
            I => \N__27151\
        );

    \I__4845\ : Span4Mux_h
    port map (
            O => \N__27215\,
            I => \N__27151\
        );

    \I__4844\ : Span4Mux_h
    port map (
            O => \N__27212\,
            I => \N__27144\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__27209\,
            I => \N__27144\
        );

    \I__4842\ : Span4Mux_h
    port map (
            O => \N__27202\,
            I => \N__27144\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__27199\,
            I => \N__27137\
        );

    \I__4840\ : Span12Mux_v
    port map (
            O => \N__27194\,
            I => \N__27137\
        );

    \I__4839\ : Span12Mux_h
    port map (
            O => \N__27191\,
            I => \N__27137\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__27188\,
            I => adc_state_0_adj_1117
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__27183\,
            I => adc_state_0_adj_1117
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__27180\,
            I => adc_state_0_adj_1117
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__27175\,
            I => adc_state_0_adj_1117
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__27172\,
            I => adc_state_0_adj_1117
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__27161\,
            I => adc_state_0_adj_1117
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__27156\,
            I => adc_state_0_adj_1117
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__27151\,
            I => adc_state_0_adj_1117
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__27144\,
            I => adc_state_0_adj_1117
        );

    \I__4829\ : Odrv12
    port map (
            O => \N__27137\,
            I => adc_state_0_adj_1117
        );

    \I__4828\ : InMux
    port map (
            O => \N__27116\,
            I => \N__27106\
        );

    \I__4827\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27101\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \N__27098\
        );

    \I__4825\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27092\
        );

    \I__4824\ : InMux
    port map (
            O => \N__27112\,
            I => \N__27087\
        );

    \I__4823\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27087\
        );

    \I__4822\ : InMux
    port map (
            O => \N__27110\,
            I => \N__27082\
        );

    \I__4821\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27082\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__27106\,
            I => \N__27079\
        );

    \I__4819\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27076\
        );

    \I__4818\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27073\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__27101\,
            I => \N__27070\
        );

    \I__4816\ : InMux
    port map (
            O => \N__27098\,
            I => \N__27067\
        );

    \I__4815\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27060\
        );

    \I__4814\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27060\
        );

    \I__4813\ : InMux
    port map (
            O => \N__27095\,
            I => \N__27060\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__27092\,
            I => \N__27053\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__27087\,
            I => \N__27053\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27053\
        );

    \I__4809\ : Span4Mux_v
    port map (
            O => \N__27079\,
            I => \N__27048\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__27076\,
            I => \N__27048\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__27073\,
            I => \DTRIG_N_957_adj_1150\
        );

    \I__4806\ : Odrv12
    port map (
            O => \N__27070\,
            I => \DTRIG_N_957_adj_1150\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__27067\,
            I => \DTRIG_N_957_adj_1150\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__27060\,
            I => \DTRIG_N_957_adj_1150\
        );

    \I__4803\ : Odrv4
    port map (
            O => \N__27053\,
            I => \DTRIG_N_957_adj_1150\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__27048\,
            I => \DTRIG_N_957_adj_1150\
        );

    \I__4801\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27030\
        );

    \I__4800\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27027\
        );

    \I__4799\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27024\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__27030\,
            I => \N__27019\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27011\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27011\
        );

    \I__4795\ : InMux
    port map (
            O => \N__27023\,
            I => \N__27002\
        );

    \I__4794\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27002\
        );

    \I__4793\ : Span4Mux_v
    port map (
            O => \N__27019\,
            I => \N__26999\
        );

    \I__4792\ : InMux
    port map (
            O => \N__27018\,
            I => \N__26992\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27017\,
            I => \N__26992\
        );

    \I__4790\ : InMux
    port map (
            O => \N__27016\,
            I => \N__26992\
        );

    \I__4789\ : Span4Mux_h
    port map (
            O => \N__27011\,
            I => \N__26989\
        );

    \I__4788\ : InMux
    port map (
            O => \N__27010\,
            I => \N__26982\
        );

    \I__4787\ : InMux
    port map (
            O => \N__27009\,
            I => \N__26982\
        );

    \I__4786\ : InMux
    port map (
            O => \N__27008\,
            I => \N__26982\
        );

    \I__4785\ : InMux
    port map (
            O => \N__27007\,
            I => \N__26979\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__27002\,
            I => \N__26976\
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__26999\,
            I => adc_state_1_adj_1116
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__26992\,
            I => adc_state_1_adj_1116
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__26989\,
            I => adc_state_1_adj_1116
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__26982\,
            I => adc_state_1_adj_1116
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__26979\,
            I => adc_state_1_adj_1116
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__26976\,
            I => adc_state_1_adj_1116
        );

    \I__4777\ : CEMux
    port map (
            O => \N__26963\,
            I => \N__26959\
        );

    \I__4776\ : CEMux
    port map (
            O => \N__26962\,
            I => \N__26956\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__26959\,
            I => \N__26951\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__26956\,
            I => \N__26951\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__26951\,
            I => \ADC_VAC4.n12\
        );

    \I__4772\ : SRMux
    port map (
            O => \N__26948\,
            I => \N__26945\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__26945\,
            I => \N__26942\
        );

    \I__4770\ : Odrv12
    port map (
            O => \N__26942\,
            I => \ADC_VAC4.n14930\
        );

    \I__4769\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26935\
        );

    \I__4768\ : InMux
    port map (
            O => \N__26938\,
            I => \N__26932\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__26935\,
            I => \comm_spi.n10467\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__26932\,
            I => \comm_spi.n10467\
        );

    \I__4765\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__26924\,
            I => \N__26920\
        );

    \I__4763\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26917\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__26920\,
            I => \comm_spi.n10468\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__26917\,
            I => \comm_spi.n10468\
        );

    \I__4760\ : SRMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__26909\,
            I => \N__26906\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__26906\,
            I => \N__26903\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__26903\,
            I => \comm_spi.data_tx_7__N_822\
        );

    \I__4756\ : IoInMux
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__26897\,
            I => \N__26894\
        );

    \I__4754\ : IoSpan4Mux
    port map (
            O => \N__26894\,
            I => \N__26891\
        );

    \I__4753\ : Span4Mux_s0_v
    port map (
            O => \N__26891\,
            I => \N__26888\
        );

    \I__4752\ : Sp12to4
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__4751\ : Span12Mux_h
    port map (
            O => \N__26885\,
            I => \N__26882\
        );

    \I__4750\ : Odrv12
    port map (
            O => \N__26882\,
            I => \DDS_CS1\
        );

    \I__4749\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26870\
        );

    \I__4748\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26870\
        );

    \I__4747\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26870\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__26870\,
            I => \N__26867\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__26867\,
            I => \N__26864\
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__26864\,
            I => comm_tx_buf_7
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__26861\,
            I => \n15156_cascade_\
        );

    \I__4742\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26829\
        );

    \I__4741\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26820\
        );

    \I__4740\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26820\
        );

    \I__4739\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26820\
        );

    \I__4738\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26820\
        );

    \I__4737\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26813\
        );

    \I__4736\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26813\
        );

    \I__4735\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26813\
        );

    \I__4734\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26807\
        );

    \I__4733\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26804\
        );

    \I__4732\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26801\
        );

    \I__4731\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26798\
        );

    \I__4730\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26794\
        );

    \I__4729\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26791\
        );

    \I__4728\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26782\
        );

    \I__4727\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26782\
        );

    \I__4726\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26782\
        );

    \I__4725\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26782\
        );

    \I__4724\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26775\
        );

    \I__4723\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26775\
        );

    \I__4722\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26775\
        );

    \I__4721\ : InMux
    port map (
            O => \N__26837\,
            I => \N__26762\
        );

    \I__4720\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26762\
        );

    \I__4719\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26762\
        );

    \I__4718\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26762\
        );

    \I__4717\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26762\
        );

    \I__4716\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26762\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26757\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26757\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__26813\,
            I => \N__26754\
        );

    \I__4712\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26746\
        );

    \I__4711\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26746\
        );

    \I__4710\ : InMux
    port map (
            O => \N__26810\,
            I => \N__26746\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__26807\,
            I => \N__26743\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__26804\,
            I => \N__26736\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26736\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__26798\,
            I => \N__26736\
        );

    \I__4705\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26733\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__26794\,
            I => \N__26722\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__26791\,
            I => \N__26722\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__26782\,
            I => \N__26722\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__26775\,
            I => \N__26722\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__26762\,
            I => \N__26722\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__26757\,
            I => \N__26719\
        );

    \I__4698\ : Span4Mux_v
    port map (
            O => \N__26754\,
            I => \N__26716\
        );

    \I__4697\ : InMux
    port map (
            O => \N__26753\,
            I => \N__26713\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26710\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__26743\,
            I => \N__26705\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__26736\,
            I => \N__26705\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__26733\,
            I => \N__26700\
        );

    \I__4692\ : Span12Mux_v
    port map (
            O => \N__26722\,
            I => \N__26700\
        );

    \I__4691\ : Span4Mux_h
    port map (
            O => \N__26719\,
            I => \N__26695\
        );

    \I__4690\ : Span4Mux_v
    port map (
            O => \N__26716\,
            I => \N__26695\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__26713\,
            I => n9694
        );

    \I__4688\ : Odrv12
    port map (
            O => \N__26710\,
            I => n9694
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__26705\,
            I => n9694
        );

    \I__4686\ : Odrv12
    port map (
            O => \N__26700\,
            I => n9694
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__26695\,
            I => n9694
        );

    \I__4684\ : CascadeMux
    port map (
            O => \N__26684\,
            I => \ADC_VAC4.n15257_cascade_\
        );

    \I__4683\ : CEMux
    port map (
            O => \N__26681\,
            I => \N__26678\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__26678\,
            I => \ADC_VAC4.n15258\
        );

    \I__4681\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26672\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__26672\,
            I => \ADC_VAC4.n15278\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__26669\,
            I => \N__26666\
        );

    \I__4678\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26661\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__26665\,
            I => \N__26658\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__26664\,
            I => \N__26654\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__26661\,
            I => \N__26651\
        );

    \I__4674\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26648\
        );

    \I__4673\ : InMux
    port map (
            O => \N__26657\,
            I => \N__26643\
        );

    \I__4672\ : InMux
    port map (
            O => \N__26654\,
            I => \N__26643\
        );

    \I__4671\ : Span4Mux_h
    port map (
            O => \N__26651\,
            I => \N__26638\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__26648\,
            I => \N__26638\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__26643\,
            I => \N__26633\
        );

    \I__4668\ : Span4Mux_v
    port map (
            O => \N__26638\,
            I => \N__26630\
        );

    \I__4667\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26625\
        );

    \I__4666\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26625\
        );

    \I__4665\ : Span12Mux_v
    port map (
            O => \N__26633\,
            I => \N__26620\
        );

    \I__4664\ : Sp12to4
    port map (
            O => \N__26630\,
            I => \N__26620\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__26625\,
            I => \N__26617\
        );

    \I__4662\ : Span12Mux_h
    port map (
            O => \N__26620\,
            I => \N__26614\
        );

    \I__4661\ : Span12Mux_h
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__4660\ : Odrv12
    port map (
            O => \N__26614\,
            I => \M_DRDY4\
        );

    \I__4659\ : Odrv12
    port map (
            O => \N__26611\,
            I => \M_DRDY4\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__26606\,
            I => \n14_cascade_\
        );

    \I__4657\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__26597\,
            I => n15156
        );

    \I__4654\ : IoInMux
    port map (
            O => \N__26594\,
            I => \N__26591\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26588\
        );

    \I__4652\ : Span4Mux_s1_v
    port map (
            O => \N__26588\,
            I => \N__26585\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__26582\,
            I => \N__26578\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__26581\,
            I => \N__26575\
        );

    \I__4648\ : Sp12to4
    port map (
            O => \N__26578\,
            I => \N__26572\
        );

    \I__4647\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26569\
        );

    \I__4646\ : Odrv12
    port map (
            O => \N__26572\,
            I => \M_CS4\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__26569\,
            I => \M_CS4\
        );

    \I__4644\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__4642\ : Sp12to4
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__4641\ : Odrv12
    port map (
            O => \N__26555\,
            I => buf_data2_11
        );

    \I__4640\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26549\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26545\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__26548\,
            I => \N__26542\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__26545\,
            I => \N__26538\
        );

    \I__4636\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26535\
        );

    \I__4635\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26532\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__26538\,
            I => \N__26529\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__26535\,
            I => \N__26526\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26519\
        );

    \I__4631\ : Span4Mux_h
    port map (
            O => \N__26529\,
            I => \N__26519\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__26526\,
            I => \N__26519\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__26519\,
            I => buf_adcdata4_11
        );

    \I__4628\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26513\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__26513\,
            I => \N__26510\
        );

    \I__4626\ : Span4Mux_h
    port map (
            O => \N__26510\,
            I => \N__26507\
        );

    \I__4625\ : Span4Mux_v
    port map (
            O => \N__26507\,
            I => \N__26504\
        );

    \I__4624\ : Span4Mux_h
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__26501\,
            I => n4061
        );

    \I__4622\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__26495\,
            I => \ADC_VAC4.n17\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__26492\,
            I => \N__26489\
        );

    \I__4619\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26485\
        );

    \I__4618\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26482\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__26485\,
            I => \N__26478\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__26482\,
            I => \N__26475\
        );

    \I__4615\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26472\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__26478\,
            I => cmd_rdadctmp_26_adj_1086
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__26475\,
            I => cmd_rdadctmp_26_adj_1086
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__26472\,
            I => cmd_rdadctmp_26_adj_1086
        );

    \I__4611\ : InMux
    port map (
            O => \N__26465\,
            I => \N__26462\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__4609\ : Span4Mux_h
    port map (
            O => \N__26459\,
            I => \N__26455\
        );

    \I__4608\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26452\
        );

    \I__4607\ : Span4Mux_v
    port map (
            O => \N__26455\,
            I => \N__26448\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26445\
        );

    \I__4605\ : InMux
    port map (
            O => \N__26451\,
            I => \N__26442\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__26448\,
            I => \N__26437\
        );

    \I__4603\ : Span4Mux_v
    port map (
            O => \N__26445\,
            I => \N__26437\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__26442\,
            I => buf_adcdata3_18
        );

    \I__4601\ : Odrv4
    port map (
            O => \N__26437\,
            I => buf_adcdata3_18
        );

    \I__4600\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__4598\ : Span4Mux_h
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__26423\,
            I => n15811
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__4595\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26413\
        );

    \I__4594\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26410\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26405\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__26410\,
            I => \N__26405\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__26405\,
            I => \N__26401\
        );

    \I__4590\ : InMux
    port map (
            O => \N__26404\,
            I => \N__26398\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__26401\,
            I => cmd_rdadctmp_21_adj_1128
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__26398\,
            I => cmd_rdadctmp_21_adj_1128
        );

    \I__4587\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26389\
        );

    \I__4586\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26385\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__26389\,
            I => \N__26382\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__26388\,
            I => \N__26379\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__26385\,
            I => \N__26376\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__26382\,
            I => \N__26373\
        );

    \I__4581\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26370\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__26376\,
            I => cmd_rdadctmp_22_adj_1127
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__26373\,
            I => cmd_rdadctmp_22_adj_1127
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__26370\,
            I => cmd_rdadctmp_22_adj_1127
        );

    \I__4577\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26359\
        );

    \I__4576\ : InMux
    port map (
            O => \N__26362\,
            I => \N__26356\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26352\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__26356\,
            I => \N__26349\
        );

    \I__4573\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26346\
        );

    \I__4572\ : Span12Mux_h
    port map (
            O => \N__26352\,
            I => \N__26343\
        );

    \I__4571\ : Span4Mux_v
    port map (
            O => \N__26349\,
            I => \N__26340\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__26346\,
            I => buf_adcdata3_16
        );

    \I__4569\ : Odrv12
    port map (
            O => \N__26343\,
            I => buf_adcdata3_16
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__26340\,
            I => buf_adcdata3_16
        );

    \I__4567\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26330\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__26330\,
            I => n90
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__26327\,
            I => \N__26322\
        );

    \I__4564\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26319\
        );

    \I__4563\ : InMux
    port map (
            O => \N__26325\,
            I => \N__26314\
        );

    \I__4562\ : InMux
    port map (
            O => \N__26322\,
            I => \N__26314\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__26319\,
            I => cmd_rdadctmp_23_adj_1126
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__26314\,
            I => cmd_rdadctmp_23_adj_1126
        );

    \I__4559\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26304\
        );

    \I__4558\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26299\
        );

    \I__4557\ : InMux
    port map (
            O => \N__26307\,
            I => \N__26299\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__26304\,
            I => cmd_rdadctmp_24_adj_1125
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__26299\,
            I => cmd_rdadctmp_24_adj_1125
        );

    \I__4554\ : CascadeMux
    port map (
            O => \N__26294\,
            I => \N__26290\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__26293\,
            I => \N__26286\
        );

    \I__4552\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26281\
        );

    \I__4551\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26281\
        );

    \I__4550\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26278\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__26281\,
            I => \N__26275\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__26278\,
            I => \N__26272\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__26275\,
            I => cmd_rdadctmp_25_adj_1124
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__26272\,
            I => cmd_rdadctmp_25_adj_1124
        );

    \I__4545\ : IoInMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__4543\ : Span4Mux_s1_v
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__4542\ : Sp12to4
    port map (
            O => \N__26258\,
            I => \N__26254\
        );

    \I__4541\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26250\
        );

    \I__4540\ : Span12Mux_h
    port map (
            O => \N__26254\,
            I => \N__26247\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__26253\,
            I => \N__26244\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__26250\,
            I => \N__26241\
        );

    \I__4537\ : Span12Mux_v
    port map (
            O => \N__26247\,
            I => \N__26238\
        );

    \I__4536\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26235\
        );

    \I__4535\ : Span4Mux_h
    port map (
            O => \N__26241\,
            I => \N__26232\
        );

    \I__4534\ : Odrv12
    port map (
            O => \N__26238\,
            I => \M_POW\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__26235\,
            I => \M_POW\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__26232\,
            I => \M_POW\
        );

    \I__4531\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__26219\,
            I => \N__26216\
        );

    \I__4528\ : Span4Mux_h
    port map (
            O => \N__26216\,
            I => \N__26213\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__26213\,
            I => \N__26208\
        );

    \I__4526\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26205\
        );

    \I__4525\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26202\
        );

    \I__4524\ : Span4Mux_h
    port map (
            O => \N__26208\,
            I => \N__26199\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__26205\,
            I => buf_adcdata3_19
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__26202\,
            I => buf_adcdata3_19
        );

    \I__4521\ : Odrv4
    port map (
            O => \N__26199\,
            I => buf_adcdata3_19
        );

    \I__4520\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26189\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__26189\,
            I => n87
        );

    \I__4518\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26172\
        );

    \I__4517\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26172\
        );

    \I__4516\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26167\
        );

    \I__4515\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26167\
        );

    \I__4514\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26164\
        );

    \I__4513\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26154\
        );

    \I__4512\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26149\
        );

    \I__4511\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26149\
        );

    \I__4510\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26144\
        );

    \I__4509\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26144\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__26172\,
            I => \N__26139\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__26167\,
            I => \N__26139\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26136\
        );

    \I__4505\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26131\
        );

    \I__4504\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26131\
        );

    \I__4503\ : InMux
    port map (
            O => \N__26161\,
            I => \N__26128\
        );

    \I__4502\ : InMux
    port map (
            O => \N__26160\,
            I => \N__26117\
        );

    \I__4501\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26117\
        );

    \I__4500\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26117\
        );

    \I__4499\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26117\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26110\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__26149\,
            I => \N__26105\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__26144\,
            I => \N__26105\
        );

    \I__4495\ : Span4Mux_v
    port map (
            O => \N__26139\,
            I => \N__26096\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__26136\,
            I => \N__26096\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26096\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__26128\,
            I => \N__26096\
        );

    \I__4491\ : InMux
    port map (
            O => \N__26127\,
            I => \N__26093\
        );

    \I__4490\ : InMux
    port map (
            O => \N__26126\,
            I => \N__26090\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__26117\,
            I => \N__26085\
        );

    \I__4488\ : InMux
    port map (
            O => \N__26116\,
            I => \N__26076\
        );

    \I__4487\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26076\
        );

    \I__4486\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26076\
        );

    \I__4485\ : InMux
    port map (
            O => \N__26113\,
            I => \N__26076\
        );

    \I__4484\ : Span4Mux_h
    port map (
            O => \N__26110\,
            I => \N__26066\
        );

    \I__4483\ : Span4Mux_h
    port map (
            O => \N__26105\,
            I => \N__26063\
        );

    \I__4482\ : Span4Mux_h
    port map (
            O => \N__26096\,
            I => \N__26058\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26058\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__26090\,
            I => \N__26055\
        );

    \I__4479\ : InMux
    port map (
            O => \N__26089\,
            I => \N__26050\
        );

    \I__4478\ : InMux
    port map (
            O => \N__26088\,
            I => \N__26050\
        );

    \I__4477\ : Span4Mux_h
    port map (
            O => \N__26085\,
            I => \N__26045\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__26076\,
            I => \N__26045\
        );

    \I__4475\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26030\
        );

    \I__4474\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26030\
        );

    \I__4473\ : InMux
    port map (
            O => \N__26073\,
            I => \N__26030\
        );

    \I__4472\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26030\
        );

    \I__4471\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26030\
        );

    \I__4470\ : InMux
    port map (
            O => \N__26070\,
            I => \N__26030\
        );

    \I__4469\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26030\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__26066\,
            I => n8272
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__26063\,
            I => n8272
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__26058\,
            I => n8272
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__26055\,
            I => n8272
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__26050\,
            I => n8272
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__26045\,
            I => n8272
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__26030\,
            I => n8272
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__26015\,
            I => \n4_adj_1264_cascade_\
        );

    \I__4460\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__4458\ : Odrv12
    port map (
            O => \N__26006\,
            I => n8055
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__26003\,
            I => \N__25999\
        );

    \I__4456\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25996\
        );

    \I__4455\ : InMux
    port map (
            O => \N__25999\,
            I => \N__25992\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__25996\,
            I => \N__25989\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__25995\,
            I => \N__25986\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25983\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__25989\,
            I => \N__25980\
        );

    \I__4450\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25977\
        );

    \I__4449\ : Span12Mux_v
    port map (
            O => \N__25983\,
            I => \N__25972\
        );

    \I__4448\ : Sp12to4
    port map (
            O => \N__25980\,
            I => \N__25972\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__25977\,
            I => buf_adcdata4_15
        );

    \I__4446\ : Odrv12
    port map (
            O => \N__25972\,
            I => buf_adcdata4_15
        );

    \I__4445\ : CascadeMux
    port map (
            O => \N__25967\,
            I => \N__25963\
        );

    \I__4444\ : InMux
    port map (
            O => \N__25966\,
            I => \N__25957\
        );

    \I__4443\ : InMux
    port map (
            O => \N__25963\,
            I => \N__25952\
        );

    \I__4442\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25952\
        );

    \I__4441\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25949\
        );

    \I__4440\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25946\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25932\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__25952\,
            I => \N__25932\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__25949\,
            I => \N__25927\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__25946\,
            I => \N__25927\
        );

    \I__4435\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25917\
        );

    \I__4434\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25910\
        );

    \I__4433\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25910\
        );

    \I__4432\ : InMux
    port map (
            O => \N__25942\,
            I => \N__25910\
        );

    \I__4431\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25905\
        );

    \I__4430\ : InMux
    port map (
            O => \N__25940\,
            I => \N__25905\
        );

    \I__4429\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25898\
        );

    \I__4428\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25898\
        );

    \I__4427\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25898\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__25932\,
            I => \N__25894\
        );

    \I__4425\ : Span4Mux_h
    port map (
            O => \N__25927\,
            I => \N__25891\
        );

    \I__4424\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25884\
        );

    \I__4423\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25884\
        );

    \I__4422\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25884\
        );

    \I__4421\ : InMux
    port map (
            O => \N__25923\,
            I => \N__25875\
        );

    \I__4420\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25875\
        );

    \I__4419\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25875\
        );

    \I__4418\ : InMux
    port map (
            O => \N__25920\,
            I => \N__25872\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__25917\,
            I => \N__25869\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__25910\,
            I => \N__25866\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25861\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__25898\,
            I => \N__25861\
        );

    \I__4413\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25858\
        );

    \I__4412\ : Span4Mux_h
    port map (
            O => \N__25894\,
            I => \N__25853\
        );

    \I__4411\ : Span4Mux_v
    port map (
            O => \N__25891\,
            I => \N__25853\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__25884\,
            I => \N__25850\
        );

    \I__4409\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25847\
        );

    \I__4408\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25844\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__25875\,
            I => \N__25841\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__25872\,
            I => \N__25836\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__25869\,
            I => \N__25836\
        );

    \I__4404\ : Span4Mux_v
    port map (
            O => \N__25866\,
            I => \N__25833\
        );

    \I__4403\ : Span4Mux_v
    port map (
            O => \N__25861\,
            I => \N__25830\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25825\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__25853\,
            I => \N__25825\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__25850\,
            I => \N__25822\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__25847\,
            I => \N__25811\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__25844\,
            I => \N__25811\
        );

    \I__4397\ : Span4Mux_h
    port map (
            O => \N__25841\,
            I => \N__25811\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__25836\,
            I => \N__25811\
        );

    \I__4395\ : Span4Mux_v
    port map (
            O => \N__25833\,
            I => \N__25811\
        );

    \I__4394\ : Span4Mux_h
    port map (
            O => \N__25830\,
            I => \N__25806\
        );

    \I__4393\ : Span4Mux_v
    port map (
            O => \N__25825\,
            I => \N__25806\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__25822\,
            I => n15144
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__25811\,
            I => n15144
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__25806\,
            I => n15144
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__25799\,
            I => \N__25795\
        );

    \I__4388\ : InMux
    port map (
            O => \N__25798\,
            I => \N__25792\
        );

    \I__4387\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25789\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__25792\,
            I => \N__25786\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25783\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__25786\,
            I => \N__25780\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__25783\,
            I => \N__25776\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__25780\,
            I => \N__25773\
        );

    \I__4381\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25770\
        );

    \I__4380\ : Span4Mux_h
    port map (
            O => \N__25776\,
            I => \N__25767\
        );

    \I__4379\ : Span4Mux_h
    port map (
            O => \N__25773\,
            I => \N__25764\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__25770\,
            I => buf_adcdata4_17
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__25767\,
            I => buf_adcdata4_17
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__25764\,
            I => buf_adcdata4_17
        );

    \I__4375\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25754\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__25754\,
            I => n71
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__4372\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__25745\,
            I => \N__25742\
        );

    \I__4370\ : Span4Mux_v
    port map (
            O => \N__25742\,
            I => \N__25737\
        );

    \I__4369\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25734\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__25740\,
            I => \N__25731\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__25737\,
            I => \N__25728\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__25734\,
            I => \N__25725\
        );

    \I__4365\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25722\
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__25728\,
            I => cmd_rdadctmp_26_adj_1123
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__25725\,
            I => cmd_rdadctmp_26_adj_1123
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__25722\,
            I => cmd_rdadctmp_26_adj_1123
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__25715\,
            I => \N__25712\
        );

    \I__4360\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25709\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__25709\,
            I => \N__25704\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__25708\,
            I => \N__25701\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__25707\,
            I => \N__25698\
        );

    \I__4356\ : Span4Mux_v
    port map (
            O => \N__25704\,
            I => \N__25695\
        );

    \I__4355\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25690\
        );

    \I__4354\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25690\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__25695\,
            I => cmd_rdadctmp_27_adj_1085
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__25690\,
            I => cmd_rdadctmp_27_adj_1085
        );

    \I__4351\ : InMux
    port map (
            O => \N__25685\,
            I => \N__25682\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__25679\,
            I => \N__25676\
        );

    \I__4348\ : Sp12to4
    port map (
            O => \N__25676\,
            I => \N__25673\
        );

    \I__4347\ : Span12Mux_h
    port map (
            O => \N__25673\,
            I => \N__25670\
        );

    \I__4346\ : Span12Mux_v
    port map (
            O => \N__25670\,
            I => \N__25665\
        );

    \I__4345\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25660\
        );

    \I__4344\ : InMux
    port map (
            O => \N__25668\,
            I => \N__25660\
        );

    \I__4343\ : Odrv12
    port map (
            O => \N__25665\,
            I => buf_adcdata3_23
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__25660\,
            I => buf_adcdata3_23
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__25655\,
            I => \N__25652\
        );

    \I__4340\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25648\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__25651\,
            I => \N__25644\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__25648\,
            I => \N__25641\
        );

    \I__4337\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25638\
        );

    \I__4336\ : InMux
    port map (
            O => \N__25644\,
            I => \N__25635\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__25641\,
            I => \N__25632\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__25638\,
            I => cmd_rdadctmp_27_adj_1122
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__25635\,
            I => cmd_rdadctmp_27_adj_1122
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__25632\,
            I => cmd_rdadctmp_27_adj_1122
        );

    \I__4331\ : CascadeMux
    port map (
            O => \N__25625\,
            I => \N__25621\
        );

    \I__4330\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25618\
        );

    \I__4329\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25615\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__25618\,
            I => \N__25612\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__25615\,
            I => \N__25609\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__25612\,
            I => \N__25606\
        );

    \I__4325\ : Span4Mux_v
    port map (
            O => \N__25609\,
            I => \N__25602\
        );

    \I__4324\ : Span4Mux_v
    port map (
            O => \N__25606\,
            I => \N__25599\
        );

    \I__4323\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25596\
        );

    \I__4322\ : Span4Mux_v
    port map (
            O => \N__25602\,
            I => \N__25593\
        );

    \I__4321\ : Span4Mux_h
    port map (
            O => \N__25599\,
            I => \N__25588\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__25596\,
            I => \N__25588\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__25593\,
            I => cmd_rdadctmp_28_adj_1121
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__25588\,
            I => cmd_rdadctmp_28_adj_1121
        );

    \I__4317\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25576\
        );

    \I__4316\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25576\
        );

    \I__4315\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25573\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__25576\,
            I => \N__25568\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__25573\,
            I => \N__25565\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__25572\,
            I => \N__25562\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__25571\,
            I => \N__25559\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__25568\,
            I => \N__25555\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__25565\,
            I => \N__25552\
        );

    \I__4308\ : InMux
    port map (
            O => \N__25562\,
            I => \N__25545\
        );

    \I__4307\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25545\
        );

    \I__4306\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25545\
        );

    \I__4305\ : Span4Mux_h
    port map (
            O => \N__25555\,
            I => \N__25542\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__25552\,
            I => \N__25539\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__25545\,
            I => n15221
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__25542\,
            I => n15221
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__25539\,
            I => n15221
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__25532\,
            I => \n17_cascade_\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__25529\,
            I => \n8702_cascade_\
        );

    \I__4298\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25520\
        );

    \I__4297\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25520\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__25520\,
            I => bit_cnt_3
        );

    \I__4295\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25508\
        );

    \I__4294\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25508\
        );

    \I__4293\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25508\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__25508\,
            I => bit_cnt_2
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__25505\,
            I => \N__25501\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__25504\,
            I => \N__25496\
        );

    \I__4289\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25490\
        );

    \I__4288\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25490\
        );

    \I__4287\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25485\
        );

    \I__4286\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25485\
        );

    \I__4285\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25482\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__25490\,
            I => \N__25477\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__25485\,
            I => \N__25477\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__25482\,
            I => \N__25472\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__25477\,
            I => \N__25472\
        );

    \I__4280\ : Odrv4
    port map (
            O => \N__25472\,
            I => bit_cnt_0
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__25469\,
            I => \n16524_cascade_\
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__25466\,
            I => \n16527_cascade_\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__25463\,
            I => \n15565_cascade_\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__25460\,
            I => \n13_adj_1257_cascade_\
        );

    \I__4275\ : CEMux
    port map (
            O => \N__25457\,
            I => \N__25454\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__25454\,
            I => \N__25451\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__25451\,
            I => \N__25445\
        );

    \I__4272\ : CEMux
    port map (
            O => \N__25450\,
            I => \N__25442\
        );

    \I__4271\ : CEMux
    port map (
            O => \N__25449\,
            I => \N__25439\
        );

    \I__4270\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25436\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__25445\,
            I => \N__25427\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__25442\,
            I => \N__25427\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25427\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__25436\,
            I => \N__25427\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__25427\,
            I => \N__25424\
        );

    \I__4264\ : Odrv4
    port map (
            O => \N__25424\,
            I => n8823
        );

    \I__4263\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25418\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__25418\,
            I => \N__25414\
        );

    \I__4261\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25411\
        );

    \I__4260\ : Odrv4
    port map (
            O => \N__25414\,
            I => n41
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__25411\,
            I => n41
        );

    \I__4258\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25403\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__25403\,
            I => n13457
        );

    \I__4256\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25394\
        );

    \I__4255\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25394\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__25394\,
            I => n13458
        );

    \I__4253\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25388\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__25385\,
            I => \N__25382\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__25382\,
            I => \N__25379\
        );

    \I__4249\ : Span4Mux_h
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__4248\ : Span4Mux_v
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__25373\,
            I => buf_data4_13
        );

    \I__4246\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__25367\,
            I => \N__25364\
        );

    \I__4244\ : Span4Mux_h
    port map (
            O => \N__25364\,
            I => \N__25361\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__25361\,
            I => comm_buf_10_5
        );

    \I__4242\ : CEMux
    port map (
            O => \N__25358\,
            I => \N__25352\
        );

    \I__4241\ : CEMux
    port map (
            O => \N__25357\,
            I => \N__25349\
        );

    \I__4240\ : CEMux
    port map (
            O => \N__25356\,
            I => \N__25346\
        );

    \I__4239\ : CEMux
    port map (
            O => \N__25355\,
            I => \N__25343\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__25352\,
            I => \N__25340\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__25349\,
            I => \N__25337\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__25346\,
            I => \N__25334\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__25343\,
            I => \N__25331\
        );

    \I__4234\ : Span4Mux_v
    port map (
            O => \N__25340\,
            I => \N__25326\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__25337\,
            I => \N__25326\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__25334\,
            I => n9045
        );

    \I__4231\ : Odrv12
    port map (
            O => \N__25331\,
            I => n9045
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__25326\,
            I => n9045
        );

    \I__4229\ : SRMux
    port map (
            O => \N__25319\,
            I => \N__25314\
        );

    \I__4228\ : SRMux
    port map (
            O => \N__25318\,
            I => \N__25310\
        );

    \I__4227\ : SRMux
    port map (
            O => \N__25317\,
            I => \N__25307\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__25314\,
            I => \N__25304\
        );

    \I__4225\ : SRMux
    port map (
            O => \N__25313\,
            I => \N__25301\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__25310\,
            I => \N__25298\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__25307\,
            I => \N__25295\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__25304\,
            I => \N__25292\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25289\
        );

    \I__4220\ : Span4Mux_v
    port map (
            O => \N__25298\,
            I => \N__25284\
        );

    \I__4219\ : Span4Mux_v
    port map (
            O => \N__25295\,
            I => \N__25284\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__25292\,
            I => n10646
        );

    \I__4217\ : Odrv12
    port map (
            O => \N__25289\,
            I => n10646
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__25284\,
            I => n10646
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__25277\,
            I => \n11_adj_1279_cascade_\
        );

    \I__4214\ : CEMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25262\
        );

    \I__4212\ : CEMux
    port map (
            O => \N__25270\,
            I => \N__25259\
        );

    \I__4211\ : CEMux
    port map (
            O => \N__25269\,
            I => \N__25256\
        );

    \I__4210\ : CEMux
    port map (
            O => \N__25268\,
            I => \N__25253\
        );

    \I__4209\ : CEMux
    port map (
            O => \N__25267\,
            I => \N__25250\
        );

    \I__4208\ : CEMux
    port map (
            O => \N__25266\,
            I => \N__25247\
        );

    \I__4207\ : CEMux
    port map (
            O => \N__25265\,
            I => \N__25244\
        );

    \I__4206\ : Span4Mux_v
    port map (
            O => \N__25262\,
            I => \N__25239\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__25259\,
            I => \N__25239\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__25256\,
            I => \N__25234\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25234\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__25250\,
            I => \N__25231\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__25247\,
            I => \N__25228\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25225\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__25239\,
            I => \N__25221\
        );

    \I__4198\ : Span4Mux_v
    port map (
            O => \N__25234\,
            I => \N__25218\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__25231\,
            I => \N__25213\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__25228\,
            I => \N__25213\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__25225\,
            I => \N__25210\
        );

    \I__4194\ : InMux
    port map (
            O => \N__25224\,
            I => \N__25207\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__25221\,
            I => n8654
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__25218\,
            I => n8654
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__25213\,
            I => n8654
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__25210\,
            I => n8654
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__25207\,
            I => n8654
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__25196\,
            I => \N__25193\
        );

    \I__4187\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25189\
        );

    \I__4186\ : InMux
    port map (
            O => \N__25192\,
            I => \N__25186\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__25189\,
            I => \N__25183\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__25186\,
            I => \N__25180\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__25183\,
            I => n5
        );

    \I__4182\ : Odrv12
    port map (
            O => \N__25180\,
            I => n5
        );

    \I__4181\ : CEMux
    port map (
            O => \N__25175\,
            I => \N__25172\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__25172\,
            I => \N__25169\
        );

    \I__4179\ : Odrv12
    port map (
            O => \N__25169\,
            I => n8763
        );

    \I__4178\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25162\
        );

    \I__4177\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25159\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__25162\,
            I => n13470
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__25159\,
            I => n13470
        );

    \I__4174\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25151\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__25151\,
            I => n13497
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__25148\,
            I => \n13497_cascade_\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \n9045_cascade_\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__25142\,
            I => \N__25139\
        );

    \I__4169\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25136\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__25136\,
            I => \N__25133\
        );

    \I__4167\ : Span4Mux_h
    port map (
            O => \N__25133\,
            I => \N__25130\
        );

    \I__4166\ : Odrv4
    port map (
            O => \N__25130\,
            I => comm_buf_11_6
        );

    \I__4165\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__4163\ : Span4Mux_h
    port map (
            O => \N__25121\,
            I => \N__25118\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__25118\,
            I => n16488
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__4160\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__25109\,
            I => \N__25106\
        );

    \I__4158\ : Span4Mux_v
    port map (
            O => \N__25106\,
            I => \N__25103\
        );

    \I__4157\ : Span4Mux_h
    port map (
            O => \N__25103\,
            I => \N__25100\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__4155\ : Odrv4
    port map (
            O => \N__25097\,
            I => buf_data4_14
        );

    \I__4154\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25091\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__25091\,
            I => comm_buf_10_6
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__25088\,
            I => \n13457_cascade_\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__25085\,
            I => \n15161_cascade_\
        );

    \I__4150\ : CEMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__4147\ : Odrv4
    port map (
            O => \N__25073\,
            I => n8997
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__25070\,
            I => \n8997_cascade_\
        );

    \I__4145\ : SRMux
    port map (
            O => \N__25067\,
            I => \N__25064\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__25064\,
            I => n10632
        );

    \I__4143\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__25046\,
            I => buf_data4_16
        );

    \I__4137\ : InMux
    port map (
            O => \N__25043\,
            I => \N__25040\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__25040\,
            I => \N__25037\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__25037\,
            I => \N__25034\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__25034\,
            I => comm_buf_9_0
        );

    \I__4133\ : CEMux
    port map (
            O => \N__25031\,
            I => \N__25026\
        );

    \I__4132\ : CEMux
    port map (
            O => \N__25030\,
            I => \N__25023\
        );

    \I__4131\ : InMux
    port map (
            O => \N__25029\,
            I => \N__25020\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__25026\,
            I => n9027
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__25023\,
            I => n9027
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__25020\,
            I => n9027
        );

    \I__4127\ : SRMux
    port map (
            O => \N__25013\,
            I => \N__25009\
        );

    \I__4126\ : SRMux
    port map (
            O => \N__25012\,
            I => \N__25006\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24998\
        );

    \I__4123\ : Span4Mux_h
    port map (
            O => \N__25003\,
            I => \N__24998\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__24998\,
            I => n10639
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__4120\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__4118\ : Span4Mux_h
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__24983\,
            I => comm_buf_11_1
        );

    \I__4116\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24977\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__4114\ : Span4Mux_v
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__4113\ : Span4Mux_h
    port map (
            O => \N__24971\,
            I => \N__24968\
        );

    \I__4112\ : Odrv4
    port map (
            O => \N__24968\,
            I => n16422
        );

    \I__4111\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__4109\ : Span4Mux_h
    port map (
            O => \N__24959\,
            I => \N__24956\
        );

    \I__4108\ : Span4Mux_v
    port map (
            O => \N__24956\,
            I => \N__24953\
        );

    \I__4107\ : Span4Mux_v
    port map (
            O => \N__24953\,
            I => \N__24950\
        );

    \I__4106\ : Span4Mux_h
    port map (
            O => \N__24950\,
            I => \N__24947\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__24947\,
            I => \N__24944\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__24944\,
            I => buf_data4_9
        );

    \I__4103\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24938\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__24938\,
            I => comm_buf_10_1
        );

    \I__4101\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24929\
        );

    \I__4100\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24929\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__24929\,
            I => \N__24925\
        );

    \I__4098\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24922\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__24925\,
            I => \N__24919\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__24922\,
            I => \N__24916\
        );

    \I__4095\ : Span4Mux_v
    port map (
            O => \N__24919\,
            I => \N__24913\
        );

    \I__4094\ : Span12Mux_v
    port map (
            O => \N__24916\,
            I => \N__24910\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__24913\,
            I => comm_tx_buf_2
        );

    \I__4092\ : Odrv12
    port map (
            O => \N__24910\,
            I => comm_tx_buf_2
        );

    \I__4091\ : SRMux
    port map (
            O => \N__24905\,
            I => \N__24902\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__24902\,
            I => \N__24899\
        );

    \I__4089\ : Span4Mux_h
    port map (
            O => \N__24899\,
            I => \N__24896\
        );

    \I__4088\ : Sp12to4
    port map (
            O => \N__24896\,
            I => \N__24893\
        );

    \I__4087\ : Odrv12
    port map (
            O => \N__24893\,
            I => \comm_spi.data_tx_7__N_810\
        );

    \I__4086\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24886\
        );

    \I__4085\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24883\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__24886\,
            I => \comm_spi.n16905\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__24883\,
            I => \comm_spi.n16905\
        );

    \I__4082\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24875\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__4080\ : Span4Mux_v
    port map (
            O => \N__24872\,
            I => \N__24868\
        );

    \I__4079\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24865\
        );

    \I__4078\ : Span4Mux_h
    port map (
            O => \N__24868\,
            I => \N__24862\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24859\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__24862\,
            I => \comm_spi.n10463\
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__24859\,
            I => \comm_spi.n10463\
        );

    \I__4074\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24850\
        );

    \I__4073\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24847\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__24850\,
            I => \comm_spi.n10464\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__24847\,
            I => \comm_spi.n10464\
        );

    \I__4070\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24839\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__4067\ : Span4Mux_h
    port map (
            O => \N__24833\,
            I => \N__24830\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__24830\,
            I => \N__24827\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__24827\,
            I => buf_data4_21
        );

    \I__4064\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24821\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__24821\,
            I => \N__24818\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__24818\,
            I => \N__24815\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__24815\,
            I => comm_buf_9_5
        );

    \I__4060\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24806\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__24803\,
            I => \N__24800\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__24800\,
            I => \N__24797\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__24797\,
            I => buf_data4_22
        );

    \I__4054\ : CascadeMux
    port map (
            O => \N__24794\,
            I => \N__24791\
        );

    \I__4053\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__4051\ : Odrv12
    port map (
            O => \N__24785\,
            I => comm_buf_9_6
        );

    \I__4050\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24776\
        );

    \I__4048\ : Span4Mux_v
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__24767\,
            I => buf_data4_23
        );

    \I__4044\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24761\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24758\
        );

    \I__4042\ : Odrv12
    port map (
            O => \N__24758\,
            I => comm_buf_9_7
        );

    \I__4041\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24752\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__24752\,
            I => \N__24749\
        );

    \I__4039\ : Span4Mux_h
    port map (
            O => \N__24749\,
            I => \N__24746\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__24746\,
            I => \N__24743\
        );

    \I__4037\ : Span4Mux_h
    port map (
            O => \N__24743\,
            I => \N__24740\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__24740\,
            I => buf_data4_18
        );

    \I__4035\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24734\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__24734\,
            I => \N__24731\
        );

    \I__4033\ : Span4Mux_h
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__24728\,
            I => comm_buf_9_2
        );

    \I__4031\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24722\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__24722\,
            I => \N__24719\
        );

    \I__4029\ : Span4Mux_v
    port map (
            O => \N__24719\,
            I => \N__24716\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__24716\,
            I => \N__24713\
        );

    \I__4027\ : Span4Mux_h
    port map (
            O => \N__24713\,
            I => \N__24710\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__24710\,
            I => buf_data4_17
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__24707\,
            I => \N__24704\
        );

    \I__4024\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24701\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__24701\,
            I => \N__24698\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__24698\,
            I => \N__24695\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__24695\,
            I => comm_buf_9_1
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__24692\,
            I => \N__24688\
        );

    \I__4019\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24685\
        );

    \I__4018\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24682\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__24685\,
            I => \ADC_VAC4.bit_cnt_5\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__24682\,
            I => \ADC_VAC4.bit_cnt_5\
        );

    \I__4015\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24674\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__24674\,
            I => \ADC_VAC4.n15354\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__24671\,
            I => \ADC_VAC4.n15619_cascade_\
        );

    \I__4012\ : CEMux
    port map (
            O => \N__24668\,
            I => \N__24665\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__24665\,
            I => \ADC_VAC4.n9631\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__24662\,
            I => \ADC_VAC4.n9631_cascade_\
        );

    \I__4009\ : SRMux
    port map (
            O => \N__24659\,
            I => \N__24656\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__24656\,
            I => \ADC_VAC4.n10783\
        );

    \I__4007\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24649\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__24652\,
            I => \N__24646\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__24649\,
            I => \N__24643\
        );

    \I__4004\ : InMux
    port map (
            O => \N__24646\,
            I => \N__24640\
        );

    \I__4003\ : Span4Mux_v
    port map (
            O => \N__24643\,
            I => \N__24636\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24633\
        );

    \I__4001\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24630\
        );

    \I__4000\ : Sp12to4
    port map (
            O => \N__24636\,
            I => \N__24627\
        );

    \I__3999\ : Span4Mux_h
    port map (
            O => \N__24633\,
            I => \N__24624\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__24630\,
            I => buf_adcdata4_20
        );

    \I__3997\ : Odrv12
    port map (
            O => \N__24627\,
            I => buf_adcdata4_20
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__24624\,
            I => buf_adcdata4_20
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__24617\,
            I => \comm_spi.n16905_cascade_\
        );

    \I__3994\ : SRMux
    port map (
            O => \N__24614\,
            I => \N__24611\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__24611\,
            I => \N__24608\
        );

    \I__3992\ : Span4Mux_v
    port map (
            O => \N__24608\,
            I => \N__24605\
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__24605\,
            I => \comm_spi.data_tx_7__N_809\
        );

    \I__3990\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24599\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24596\
        );

    \I__3988\ : Span4Mux_v
    port map (
            O => \N__24596\,
            I => \N__24592\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__24595\,
            I => \N__24589\
        );

    \I__3986\ : Span4Mux_h
    port map (
            O => \N__24592\,
            I => \N__24586\
        );

    \I__3985\ : InMux
    port map (
            O => \N__24589\,
            I => \N__24583\
        );

    \I__3984\ : Span4Mux_h
    port map (
            O => \N__24586\,
            I => \N__24580\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__24583\,
            I => buf_adcdata1_9
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__24580\,
            I => buf_adcdata1_9
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \N__24570\
        );

    \I__3980\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24565\
        );

    \I__3979\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24565\
        );

    \I__3978\ : InMux
    port map (
            O => \N__24570\,
            I => \N__24562\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__24565\,
            I => cmd_rdadctmp_17
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__24562\,
            I => cmd_rdadctmp_17
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__24557\,
            I => \N__24553\
        );

    \I__3974\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24547\
        );

    \I__3973\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24547\
        );

    \I__3972\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24544\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__24547\,
            I => cmd_rdadctmp_19
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__24544\,
            I => cmd_rdadctmp_19
        );

    \I__3969\ : InMux
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__24533\,
            I => \N__24529\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__24532\,
            I => \N__24526\
        );

    \I__3965\ : Span4Mux_h
    port map (
            O => \N__24529\,
            I => \N__24523\
        );

    \I__3964\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24520\
        );

    \I__3963\ : Span4Mux_h
    port map (
            O => \N__24523\,
            I => \N__24517\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__24520\,
            I => buf_adcdata1_11
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__24517\,
            I => buf_adcdata1_11
        );

    \I__3960\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24508\
        );

    \I__3959\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24505\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__24505\,
            I => \N__24498\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__24502\,
            I => \N__24495\
        );

    \I__3955\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24492\
        );

    \I__3954\ : Span12Mux_s10_v
    port map (
            O => \N__24498\,
            I => \N__24489\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__24495\,
            I => \N__24486\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__24492\,
            I => buf_adcdata3_8
        );

    \I__3951\ : Odrv12
    port map (
            O => \N__24489\,
            I => buf_adcdata3_8
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__24486\,
            I => buf_adcdata3_8
        );

    \I__3949\ : InMux
    port map (
            O => \N__24479\,
            I => \N__24475\
        );

    \I__3948\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24472\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__24475\,
            I => \ADC_VAC4.bit_cnt_4\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__24472\,
            I => \ADC_VAC4.bit_cnt_4\
        );

    \I__3945\ : InMux
    port map (
            O => \N__24467\,
            I => \N__24463\
        );

    \I__3944\ : InMux
    port map (
            O => \N__24466\,
            I => \N__24460\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__24463\,
            I => \ADC_VAC4.bit_cnt_3\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__24460\,
            I => \ADC_VAC4.bit_cnt_3\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__24455\,
            I => \N__24451\
        );

    \I__3940\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24448\
        );

    \I__3939\ : InMux
    port map (
            O => \N__24451\,
            I => \N__24445\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__24448\,
            I => \ADC_VAC4.bit_cnt_1\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__24445\,
            I => \ADC_VAC4.bit_cnt_1\
        );

    \I__3936\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24436\
        );

    \I__3935\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24433\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__24436\,
            I => \ADC_VAC4.bit_cnt_2\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__24433\,
            I => \ADC_VAC4.bit_cnt_2\
        );

    \I__3932\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24424\
        );

    \I__3931\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24421\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__24424\,
            I => \N__24418\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__24421\,
            I => \ADC_VAC4.bit_cnt_6\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__24418\,
            I => \ADC_VAC4.bit_cnt_6\
        );

    \I__3927\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24409\
        );

    \I__3926\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24406\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__24409\,
            I => \ADC_VAC4.bit_cnt_0\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__24406\,
            I => \ADC_VAC4.bit_cnt_0\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__24401\,
            I => \ADC_VAC4.n15330_cascade_\
        );

    \I__3922\ : InMux
    port map (
            O => \N__24398\,
            I => \N__24394\
        );

    \I__3921\ : InMux
    port map (
            O => \N__24397\,
            I => \N__24391\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__24394\,
            I => \ADC_VAC4.bit_cnt_7\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__24391\,
            I => \ADC_VAC4.bit_cnt_7\
        );

    \I__3918\ : InMux
    port map (
            O => \N__24386\,
            I => \N__24383\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__24383\,
            I => \N__24380\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__24380\,
            I => n69
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__24377\,
            I => \N__24373\
        );

    \I__3914\ : CascadeMux
    port map (
            O => \N__24376\,
            I => \N__24370\
        );

    \I__3913\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24365\
        );

    \I__3912\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24365\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__24365\,
            I => buf_control_0
        );

    \I__3910\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__3908\ : Span12Mux_h
    port map (
            O => \N__24356\,
            I => \N__24353\
        );

    \I__3907\ : Odrv12
    port map (
            O => \N__24353\,
            I => buf_data2_8
        );

    \I__3906\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24347\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24343\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__24346\,
            I => \N__24340\
        );

    \I__3903\ : Span4Mux_h
    port map (
            O => \N__24343\,
            I => \N__24337\
        );

    \I__3902\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24333\
        );

    \I__3901\ : Span4Mux_h
    port map (
            O => \N__24337\,
            I => \N__24330\
        );

    \I__3900\ : CascadeMux
    port map (
            O => \N__24336\,
            I => \N__24327\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24324\
        );

    \I__3898\ : Sp12to4
    port map (
            O => \N__24330\,
            I => \N__24321\
        );

    \I__3897\ : InMux
    port map (
            O => \N__24327\,
            I => \N__24318\
        );

    \I__3896\ : Span4Mux_h
    port map (
            O => \N__24324\,
            I => \N__24315\
        );

    \I__3895\ : Span12Mux_v
    port map (
            O => \N__24321\,
            I => \N__24312\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__24318\,
            I => buf_adcdata4_8
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__24315\,
            I => buf_adcdata4_8
        );

    \I__3892\ : Odrv12
    port map (
            O => \N__24312\,
            I => buf_adcdata4_8
        );

    \I__3891\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24302\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24299\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__24299\,
            I => \N__24296\
        );

    \I__3888\ : Span4Mux_h
    port map (
            O => \N__24296\,
            I => \N__24293\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__24293\,
            I => n4064
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__24290\,
            I => \N__24287\
        );

    \I__3885\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24283\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__24286\,
            I => \N__24280\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24277\
        );

    \I__3882\ : InMux
    port map (
            O => \N__24280\,
            I => \N__24274\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__24277\,
            I => cmd_rdadctmp_5_adj_1107
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__24274\,
            I => cmd_rdadctmp_5_adj_1107
        );

    \I__3879\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24266\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__24263\,
            I => \N__24259\
        );

    \I__3876\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24256\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__24259\,
            I => cmd_rdadctmp_6_adj_1106
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__24256\,
            I => cmd_rdadctmp_6_adj_1106
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__3872\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24245\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__24245\,
            I => \N__24241\
        );

    \I__3870\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24238\
        );

    \I__3869\ : Span4Mux_h
    port map (
            O => \N__24241\,
            I => \N__24234\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__24238\,
            I => \N__24231\
        );

    \I__3867\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24228\
        );

    \I__3866\ : Odrv4
    port map (
            O => \N__24234\,
            I => cmd_rdadctmp_28_adj_1084
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__24231\,
            I => cmd_rdadctmp_28_adj_1084
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__24228\,
            I => cmd_rdadctmp_28_adj_1084
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__24221\,
            I => \n16503_cascade_\
        );

    \I__3862\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24215\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__24215\,
            I => n4_adj_1280
        );

    \I__3860\ : CascadeMux
    port map (
            O => \N__24212\,
            I => \n8047_cascade_\
        );

    \I__3859\ : SRMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__24206\,
            I => \N__24202\
        );

    \I__3857\ : SRMux
    port map (
            O => \N__24205\,
            I => \N__24199\
        );

    \I__3856\ : Span4Mux_h
    port map (
            O => \N__24202\,
            I => \N__24194\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__24199\,
            I => \N__24194\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__24194\,
            I => \N__24189\
        );

    \I__3853\ : SRMux
    port map (
            O => \N__24193\,
            I => \N__24183\
        );

    \I__3852\ : SRMux
    port map (
            O => \N__24192\,
            I => \N__24180\
        );

    \I__3851\ : Span4Mux_h
    port map (
            O => \N__24189\,
            I => \N__24177\
        );

    \I__3850\ : SRMux
    port map (
            O => \N__24188\,
            I => \N__24174\
        );

    \I__3849\ : SRMux
    port map (
            O => \N__24187\,
            I => \N__24171\
        );

    \I__3848\ : SRMux
    port map (
            O => \N__24186\,
            I => \N__24168\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__24183\,
            I => n10576
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__24180\,
            I => n10576
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__24177\,
            I => n10576
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__24174\,
            I => n10576
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__24171\,
            I => n10576
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__24168\,
            I => n10576
        );

    \I__3841\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24151\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__24154\,
            I => \N__24148\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__24151\,
            I => \N__24145\
        );

    \I__3838\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24141\
        );

    \I__3837\ : Span4Mux_h
    port map (
            O => \N__24145\,
            I => \N__24138\
        );

    \I__3836\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24135\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__24141\,
            I => cmd_rdadctmp_9
        );

    \I__3834\ : Odrv4
    port map (
            O => \N__24138\,
            I => cmd_rdadctmp_9
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__24135\,
            I => cmd_rdadctmp_9
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__24128\,
            I => \N__24124\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__24127\,
            I => \N__24121\
        );

    \I__3830\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24116\
        );

    \I__3829\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24116\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__24116\,
            I => buf_control_3
        );

    \I__3827\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24110\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__24110\,
            I => n69_adj_1029
        );

    \I__3825\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__24104\,
            I => \N__24100\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__24103\,
            I => \N__24097\
        );

    \I__3822\ : Span4Mux_v
    port map (
            O => \N__24100\,
            I => \N__24093\
        );

    \I__3821\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24090\
        );

    \I__3820\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24087\
        );

    \I__3819\ : Sp12to4
    port map (
            O => \N__24093\,
            I => \N__24084\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__24090\,
            I => \N__24081\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__24087\,
            I => buf_adcdata4_14
        );

    \I__3816\ : Odrv12
    port map (
            O => \N__24084\,
            I => buf_adcdata4_14
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__24081\,
            I => buf_adcdata4_14
        );

    \I__3814\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24070\
        );

    \I__3813\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24067\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24064\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__24067\,
            I => \N__24061\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__24064\,
            I => \N__24057\
        );

    \I__3809\ : Span12Mux_v
    port map (
            O => \N__24061\,
            I => \N__24054\
        );

    \I__3808\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24051\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__24057\,
            I => \N__24048\
        );

    \I__3806\ : Span12Mux_h
    port map (
            O => \N__24054\,
            I => \N__24045\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__24051\,
            I => buf_adcdata3_20
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__24048\,
            I => buf_adcdata3_20
        );

    \I__3803\ : Odrv12
    port map (
            O => \N__24045\,
            I => buf_adcdata3_20
        );

    \I__3802\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24035\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__24035\,
            I => \N__24032\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__24032\,
            I => \N__24029\
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__24029\,
            I => n61
        );

    \I__3798\ : CascadeMux
    port map (
            O => \N__24026\,
            I => \N__24022\
        );

    \I__3797\ : InMux
    port map (
            O => \N__24025\,
            I => \N__24017\
        );

    \I__3796\ : InMux
    port map (
            O => \N__24022\,
            I => \N__24017\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__24017\,
            I => buf_control_4
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__3793\ : InMux
    port map (
            O => \N__24011\,
            I => \N__24002\
        );

    \I__3792\ : InMux
    port map (
            O => \N__24010\,
            I => \N__24002\
        );

    \I__3791\ : InMux
    port map (
            O => \N__24009\,
            I => \N__24002\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__24002\,
            I => cmd_rdadctmp_25_adj_1087
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__23999\,
            I => \N__23996\
        );

    \I__3788\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23993\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__23993\,
            I => \N__23989\
        );

    \I__3786\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23986\
        );

    \I__3785\ : Odrv12
    port map (
            O => \N__23989\,
            I => cmd_rdadctmp_7_adj_1105
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__23986\,
            I => cmd_rdadctmp_7_adj_1105
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__23981\,
            I => \n16500_cascade_\
        );

    \I__3782\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23975\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__23975\,
            I => \N__23972\
        );

    \I__3780\ : Span4Mux_h
    port map (
            O => \N__23972\,
            I => \N__23969\
        );

    \I__3779\ : Sp12to4
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__3778\ : Span12Mux_v
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__3777\ : Odrv12
    port map (
            O => \N__23963\,
            I => buf_data4_12
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__23960\,
            I => \N__23957\
        );

    \I__3775\ : InMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__23954\,
            I => comm_buf_10_4
        );

    \I__3773\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23945\
        );

    \I__3771\ : Span4Mux_h
    port map (
            O => \N__23945\,
            I => \N__23942\
        );

    \I__3770\ : Span4Mux_h
    port map (
            O => \N__23942\,
            I => \N__23939\
        );

    \I__3769\ : Span4Mux_h
    port map (
            O => \N__23939\,
            I => \N__23936\
        );

    \I__3768\ : Span4Mux_h
    port map (
            O => \N__23936\,
            I => \N__23933\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__23933\,
            I => buf_data4_15
        );

    \I__3766\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23927\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__3764\ : Span4Mux_v
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__3763\ : Sp12to4
    port map (
            O => \N__23921\,
            I => \N__23918\
        );

    \I__3762\ : Odrv12
    port map (
            O => \N__23918\,
            I => comm_buf_10_7
        );

    \I__3761\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23912\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23909\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__23909\,
            I => \N__23906\
        );

    \I__3758\ : Sp12to4
    port map (
            O => \N__23906\,
            I => \N__23903\
        );

    \I__3757\ : Span12Mux_h
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__3756\ : Span12Mux_v
    port map (
            O => \N__23900\,
            I => \N__23897\
        );

    \I__3755\ : Odrv12
    port map (
            O => \N__23897\,
            I => buf_data4_8
        );

    \I__3754\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__23891\,
            I => \N__23888\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__23888\,
            I => \N__23885\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__23885\,
            I => comm_buf_10_0
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__23882\,
            I => \n16434_cascade_\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__23879\,
            I => \n16437_cascade_\
        );

    \I__3748\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23873\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__23873\,
            I => n109
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__23870\,
            I => \n8054_cascade_\
        );

    \I__3745\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__23864\,
            I => \N__23861\
        );

    \I__3743\ : Odrv12
    port map (
            O => \N__23861\,
            I => n59
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__23858\,
            I => \n8907_cascade_\
        );

    \I__3741\ : CEMux
    port map (
            O => \N__23855\,
            I => \N__23852\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__23852\,
            I => n8943
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__23849\,
            I => \n8943_cascade_\
        );

    \I__3738\ : SRMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23840\
        );

    \I__3736\ : Odrv12
    port map (
            O => \N__23840\,
            I => n10625
        );

    \I__3735\ : CEMux
    port map (
            O => \N__23837\,
            I => \N__23834\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23831\
        );

    \I__3733\ : Span4Mux_h
    port map (
            O => \N__23831\,
            I => \N__23828\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__23828\,
            I => n9123
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__23825\,
            I => \n9123_cascade_\
        );

    \I__3730\ : SRMux
    port map (
            O => \N__23822\,
            I => \N__23819\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__23819\,
            I => n10653
        );

    \I__3728\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23813\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__3726\ : Sp12to4
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__3725\ : Span12Mux_v
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__3724\ : Odrv12
    port map (
            O => \N__23804\,
            I => buf_data3_16
        );

    \I__3723\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__23798\,
            I => \N__23795\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__23792\,
            I => comm_buf_6_0
        );

    \I__3719\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23786\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__23786\,
            I => \N__23783\
        );

    \I__3717\ : Sp12to4
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__3716\ : Span12Mux_v
    port map (
            O => \N__23780\,
            I => \N__23777\
        );

    \I__3715\ : Odrv12
    port map (
            O => \N__23777\,
            I => buf_data3_17
        );

    \I__3714\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__3712\ : Span4Mux_h
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__23765\,
            I => comm_buf_6_1
        );

    \I__3710\ : CEMux
    port map (
            O => \N__23762\,
            I => \N__23758\
        );

    \I__3709\ : CEMux
    port map (
            O => \N__23761\,
            I => \N__23755\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__23758\,
            I => \N__23752\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__23755\,
            I => \N__23749\
        );

    \I__3706\ : Odrv12
    port map (
            O => \N__23752\,
            I => n8907
        );

    \I__3705\ : Odrv4
    port map (
            O => \N__23749\,
            I => n8907
        );

    \I__3704\ : SRMux
    port map (
            O => \N__23744\,
            I => \N__23740\
        );

    \I__3703\ : SRMux
    port map (
            O => \N__23743\,
            I => \N__23737\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__23740\,
            I => \N__23734\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__23737\,
            I => \N__23731\
        );

    \I__3700\ : Span4Mux_h
    port map (
            O => \N__23734\,
            I => \N__23728\
        );

    \I__3699\ : Odrv12
    port map (
            O => \N__23731\,
            I => n10618
        );

    \I__3698\ : Odrv4
    port map (
            O => \N__23728\,
            I => n10618
        );

    \I__3697\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23720\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__3694\ : Sp12to4
    port map (
            O => \N__23714\,
            I => \N__23711\
        );

    \I__3693\ : Span12Mux_v
    port map (
            O => \N__23711\,
            I => \N__23708\
        );

    \I__3692\ : Odrv12
    port map (
            O => \N__23708\,
            I => buf_data4_10
        );

    \I__3691\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23702\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__23702\,
            I => \N__23699\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__23699\,
            I => \N__23696\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__23696\,
            I => comm_buf_10_2
        );

    \I__3687\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__23687\,
            I => \N__23684\
        );

    \I__3684\ : Span4Mux_v
    port map (
            O => \N__23684\,
            I => \N__23681\
        );

    \I__3683\ : Span4Mux_h
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__23678\,
            I => \N__23675\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__23675\,
            I => buf_data4_11
        );

    \I__3680\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__23669\,
            I => \N__23666\
        );

    \I__3678\ : Span4Mux_h
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__23663\,
            I => comm_buf_10_3
        );

    \I__3676\ : InMux
    port map (
            O => \N__23660\,
            I => \N__23657\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23654\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__3673\ : Sp12to4
    port map (
            O => \N__23651\,
            I => \N__23648\
        );

    \I__3672\ : Odrv12
    port map (
            O => \N__23648\,
            I => buf_data3_1
        );

    \I__3671\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__23642\,
            I => \N__23639\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__23639\,
            I => \N__23636\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__23636\,
            I => comm_buf_8_1
        );

    \I__3667\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23630\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__23630\,
            I => \N__23627\
        );

    \I__3665\ : Span4Mux_v
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__3664\ : Span4Mux_h
    port map (
            O => \N__23624\,
            I => \N__23621\
        );

    \I__3663\ : Span4Mux_h
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__23618\,
            I => buf_data3_0
        );

    \I__3661\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23609\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__23606\,
            I => comm_buf_8_0
        );

    \I__3657\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23600\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__23600\,
            I => \N__23597\
        );

    \I__3655\ : Sp12to4
    port map (
            O => \N__23597\,
            I => \N__23594\
        );

    \I__3654\ : Span12Mux_v
    port map (
            O => \N__23594\,
            I => \N__23591\
        );

    \I__3653\ : Odrv12
    port map (
            O => \N__23591\,
            I => buf_data3_23
        );

    \I__3652\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23585\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__23585\,
            I => comm_buf_6_7
        );

    \I__3650\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23579\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__3648\ : Sp12to4
    port map (
            O => \N__23576\,
            I => \N__23573\
        );

    \I__3647\ : Span12Mux_v
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__3646\ : Odrv12
    port map (
            O => \N__23570\,
            I => buf_data3_22
        );

    \I__3645\ : InMux
    port map (
            O => \N__23567\,
            I => \N__23564\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__3642\ : Span4Mux_h
    port map (
            O => \N__23558\,
            I => \N__23555\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__23555\,
            I => comm_buf_6_6
        );

    \I__3640\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__3638\ : Span4Mux_v
    port map (
            O => \N__23546\,
            I => \N__23543\
        );

    \I__3637\ : Sp12to4
    port map (
            O => \N__23543\,
            I => \N__23540\
        );

    \I__3636\ : Odrv12
    port map (
            O => \N__23540\,
            I => buf_data3_21
        );

    \I__3635\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23531\
        );

    \I__3633\ : Span12Mux_h
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__3632\ : Odrv12
    port map (
            O => \N__23528\,
            I => comm_buf_6_5
        );

    \I__3631\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23522\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__23522\,
            I => \N__23519\
        );

    \I__3629\ : Sp12to4
    port map (
            O => \N__23519\,
            I => \N__23516\
        );

    \I__3628\ : Span12Mux_v
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__3627\ : Odrv12
    port map (
            O => \N__23513\,
            I => buf_data3_20
        );

    \I__3626\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23507\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__23504\,
            I => comm_buf_6_4
        );

    \I__3623\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23495\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__3620\ : Sp12to4
    port map (
            O => \N__23492\,
            I => \N__23489\
        );

    \I__3619\ : Odrv12
    port map (
            O => \N__23489\,
            I => buf_data3_19
        );

    \I__3618\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__23483\,
            I => \N__23480\
        );

    \I__3616\ : Span4Mux_h
    port map (
            O => \N__23480\,
            I => \N__23477\
        );

    \I__3615\ : Odrv4
    port map (
            O => \N__23477\,
            I => comm_buf_6_3
        );

    \I__3614\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23471\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23468\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__23468\,
            I => \N__23465\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__23465\,
            I => \N__23462\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__23462\,
            I => \N__23459\
        );

    \I__3609\ : Span4Mux_h
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__23456\,
            I => buf_data3_18
        );

    \I__3607\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__3605\ : Span4Mux_v
    port map (
            O => \N__23447\,
            I => \N__23444\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__23441\,
            I => comm_buf_6_2
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \N__23435\
        );

    \I__3601\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23431\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__23434\,
            I => \N__23427\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23424\
        );

    \I__3598\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23419\
        );

    \I__3597\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23419\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__23424\,
            I => cmd_rdadctmp_30_adj_1119
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__23419\,
            I => cmd_rdadctmp_30_adj_1119
        );

    \I__3594\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23408\
        );

    \I__3593\ : InMux
    port map (
            O => \N__23413\,
            I => \N__23408\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__23408\,
            I => cmd_rdadctmp_31_adj_1118
        );

    \I__3591\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23402\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__3589\ : Span4Mux_v
    port map (
            O => \N__23399\,
            I => \N__23396\
        );

    \I__3588\ : Sp12to4
    port map (
            O => \N__23396\,
            I => \N__23393\
        );

    \I__3587\ : Odrv12
    port map (
            O => \N__23393\,
            I => buf_data3_7
        );

    \I__3586\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23387\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__3584\ : Odrv4
    port map (
            O => \N__23384\,
            I => comm_buf_8_7
        );

    \I__3583\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23378\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__23372\,
            I => buf_data3_6
        );

    \I__3579\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__23360\,
            I => comm_buf_8_6
        );

    \I__3575\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23354\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23351\
        );

    \I__3573\ : Span4Mux_h
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__3571\ : Odrv4
    port map (
            O => \N__23345\,
            I => buf_data3_5
        );

    \I__3570\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__23339\,
            I => \N__23336\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__23336\,
            I => comm_buf_8_5
        );

    \I__3567\ : InMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23327\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__23327\,
            I => \N__23324\
        );

    \I__3564\ : Span4Mux_h
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__23321\,
            I => buf_data3_4
        );

    \I__3562\ : InMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__23312\,
            I => \N__23309\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__23309\,
            I => comm_buf_8_4
        );

    \I__3558\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23300\
        );

    \I__3556\ : Span4Mux_v
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__3555\ : Span4Mux_h
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__3554\ : Span4Mux_h
    port map (
            O => \N__23294\,
            I => \N__23291\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__23291\,
            I => buf_data3_3
        );

    \I__3552\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23285\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__23285\,
            I => \N__23282\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__23282\,
            I => \N__23279\
        );

    \I__3549\ : Span4Mux_h
    port map (
            O => \N__23279\,
            I => \N__23276\
        );

    \I__3548\ : Odrv4
    port map (
            O => \N__23276\,
            I => comm_buf_8_3
        );

    \I__3547\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23270\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__23270\,
            I => \N__23267\
        );

    \I__3545\ : Span12Mux_h
    port map (
            O => \N__23267\,
            I => \N__23264\
        );

    \I__3544\ : Odrv12
    port map (
            O => \N__23264\,
            I => buf_data3_2
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__3542\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23255\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__23255\,
            I => \N__23252\
        );

    \I__3540\ : Span4Mux_h
    port map (
            O => \N__23252\,
            I => \N__23249\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__23249\,
            I => comm_buf_8_2
        );

    \I__3538\ : InMux
    port map (
            O => \N__23246\,
            I => \ADC_VAC4.n14007\
        );

    \I__3537\ : InMux
    port map (
            O => \N__23243\,
            I => \ADC_VAC4.n14008\
        );

    \I__3536\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23237\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__23237\,
            I => \N__23232\
        );

    \I__3534\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23229\
        );

    \I__3533\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23226\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__23232\,
            I => \comm_spi.n16908\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__23229\,
            I => \comm_spi.n16908\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__23226\,
            I => \comm_spi.n16908\
        );

    \I__3529\ : InMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23212\
        );

    \I__3527\ : InMux
    port map (
            O => \N__23215\,
            I => \N__23209\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__23212\,
            I => \comm_spi.n10459\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__23209\,
            I => \comm_spi.n10459\
        );

    \I__3524\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23201\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__23201\,
            I => \N__23197\
        );

    \I__3522\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23194\
        );

    \I__3521\ : Span4Mux_h
    port map (
            O => \N__23197\,
            I => \N__23189\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__23194\,
            I => \N__23189\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__23189\,
            I => \comm_spi.n10460\
        );

    \I__3518\ : SRMux
    port map (
            O => \N__23186\,
            I => \N__23183\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__23183\,
            I => \N__23180\
        );

    \I__3516\ : Odrv12
    port map (
            O => \N__23180\,
            I => \comm_spi.data_tx_7__N_828\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__3514\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23170\
        );

    \I__3513\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23167\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__23170\,
            I => \N__23163\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__23167\,
            I => \N__23160\
        );

    \I__3510\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23157\
        );

    \I__3509\ : Span4Mux_h
    port map (
            O => \N__23163\,
            I => \N__23154\
        );

    \I__3508\ : Span12Mux_h
    port map (
            O => \N__23160\,
            I => \N__23151\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__23157\,
            I => buf_adcdata4_21
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__23154\,
            I => buf_adcdata4_21
        );

    \I__3505\ : Odrv12
    port map (
            O => \N__23151\,
            I => buf_adcdata4_21
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__23144\,
            I => \N__23141\
        );

    \I__3503\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23132\
        );

    \I__3502\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23132\
        );

    \I__3501\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23132\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__23132\,
            I => cmd_rdadctmp_29_adj_1120
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__23129\,
            I => \N__23125\
        );

    \I__3498\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23118\
        );

    \I__3497\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23118\
        );

    \I__3496\ : CascadeMux
    port map (
            O => \N__23124\,
            I => \N__23115\
        );

    \I__3495\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23112\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__23118\,
            I => \N__23108\
        );

    \I__3493\ : InMux
    port map (
            O => \N__23115\,
            I => \N__23105\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__23112\,
            I => \N__23102\
        );

    \I__3491\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23099\
        );

    \I__3490\ : Span4Mux_v
    port map (
            O => \N__23108\,
            I => \N__23094\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__23105\,
            I => \N__23094\
        );

    \I__3488\ : Span4Mux_v
    port map (
            O => \N__23102\,
            I => \N__23091\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__23099\,
            I => \N__23088\
        );

    \I__3486\ : Span4Mux_v
    port map (
            O => \N__23094\,
            I => \N__23085\
        );

    \I__3485\ : Span4Mux_v
    port map (
            O => \N__23091\,
            I => \N__23080\
        );

    \I__3484\ : Span4Mux_v
    port map (
            O => \N__23088\,
            I => \N__23080\
        );

    \I__3483\ : Sp12to4
    port map (
            O => \N__23085\,
            I => \N__23075\
        );

    \I__3482\ : Sp12to4
    port map (
            O => \N__23080\,
            I => \N__23075\
        );

    \I__3481\ : Span12Mux_h
    port map (
            O => \N__23075\,
            I => \N__23072\
        );

    \I__3480\ : Odrv12
    port map (
            O => \N__23072\,
            I => \M_DRDY3\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__23069\,
            I => \N__23063\
        );

    \I__3478\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23059\
        );

    \I__3477\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23050\
        );

    \I__3476\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23050\
        );

    \I__3475\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23050\
        );

    \I__3474\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23046\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__23059\,
            I => \N__23043\
        );

    \I__3472\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23036\
        );

    \I__3471\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23033\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__23050\,
            I => \N__23030\
        );

    \I__3469\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23027\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__23046\,
            I => \N__23024\
        );

    \I__3467\ : Span4Mux_h
    port map (
            O => \N__23043\,
            I => \N__23021\
        );

    \I__3466\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23018\
        );

    \I__3465\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23011\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23011\
        );

    \I__3463\ : InMux
    port map (
            O => \N__23039\,
            I => \N__23011\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__23036\,
            I => \N__23004\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__23033\,
            I => \N__23004\
        );

    \I__3460\ : Span4Mux_h
    port map (
            O => \N__23030\,
            I => \N__23004\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__23027\,
            I => adc_state_1_adj_1079
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__23024\,
            I => adc_state_1_adj_1079
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__23021\,
            I => adc_state_1_adj_1079
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__23018\,
            I => adc_state_1_adj_1079
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__23011\,
            I => adc_state_1_adj_1079
        );

    \I__3454\ : Odrv4
    port map (
            O => \N__23004\,
            I => adc_state_1_adj_1079
        );

    \I__3453\ : CEMux
    port map (
            O => \N__22991\,
            I => \N__22988\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__22988\,
            I => \ADC_VAC3.n9514\
        );

    \I__3451\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22973\
        );

    \I__3450\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22973\
        );

    \I__3449\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22966\
        );

    \I__3448\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22966\
        );

    \I__3447\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22966\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__22980\,
            I => \N__22963\
        );

    \I__3445\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22960\
        );

    \I__3444\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22957\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22948\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22948\
        );

    \I__3441\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22945\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22940\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__22957\,
            I => \N__22940\
        );

    \I__3438\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22937\
        );

    \I__3437\ : InMux
    port map (
            O => \N__22955\,
            I => \N__22930\
        );

    \I__3436\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22930\
        );

    \I__3435\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22930\
        );

    \I__3434\ : Span4Mux_v
    port map (
            O => \N__22948\,
            I => \N__22927\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__22945\,
            I => \DTRIG_N_957_adj_1114\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__22940\,
            I => \DTRIG_N_957_adj_1114\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__22937\,
            I => \DTRIG_N_957_adj_1114\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__22930\,
            I => \DTRIG_N_957_adj_1114\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__22927\,
            I => \DTRIG_N_957_adj_1114\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__22916\,
            I => \ADC_VAC3.n9514_cascade_\
        );

    \I__3427\ : SRMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__22910\,
            I => \N__22907\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__22907\,
            I => \N__22904\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__22904\,
            I => \ADC_VAC3.n10744\
        );

    \I__3423\ : InMux
    port map (
            O => \N__22901\,
            I => \bfn_10_17_0_\
        );

    \I__3422\ : InMux
    port map (
            O => \N__22898\,
            I => \ADC_VAC4.n14002\
        );

    \I__3421\ : InMux
    port map (
            O => \N__22895\,
            I => \ADC_VAC4.n14003\
        );

    \I__3420\ : InMux
    port map (
            O => \N__22892\,
            I => \ADC_VAC4.n14004\
        );

    \I__3419\ : InMux
    port map (
            O => \N__22889\,
            I => \ADC_VAC4.n14005\
        );

    \I__3418\ : InMux
    port map (
            O => \N__22886\,
            I => \ADC_VAC4.n14006\
        );

    \I__3417\ : InMux
    port map (
            O => \N__22883\,
            I => \N__22879\
        );

    \I__3416\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22876\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__22879\,
            I => \ADC_VAC3.bit_cnt_0\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__22876\,
            I => \ADC_VAC3.bit_cnt_0\
        );

    \I__3413\ : InMux
    port map (
            O => \N__22871\,
            I => \bfn_10_15_0_\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__22868\,
            I => \N__22864\
        );

    \I__3411\ : InMux
    port map (
            O => \N__22867\,
            I => \N__22861\
        );

    \I__3410\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22858\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__22861\,
            I => \ADC_VAC3.bit_cnt_1\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__22858\,
            I => \ADC_VAC3.bit_cnt_1\
        );

    \I__3407\ : InMux
    port map (
            O => \N__22853\,
            I => \ADC_VAC3.n13995\
        );

    \I__3406\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22846\
        );

    \I__3405\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22843\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__22846\,
            I => \ADC_VAC3.bit_cnt_2\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__22843\,
            I => \ADC_VAC3.bit_cnt_2\
        );

    \I__3402\ : InMux
    port map (
            O => \N__22838\,
            I => \ADC_VAC3.n13996\
        );

    \I__3401\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22831\
        );

    \I__3400\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22828\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__22831\,
            I => \ADC_VAC3.bit_cnt_3\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__22828\,
            I => \ADC_VAC3.bit_cnt_3\
        );

    \I__3397\ : InMux
    port map (
            O => \N__22823\,
            I => \ADC_VAC3.n13997\
        );

    \I__3396\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22816\
        );

    \I__3395\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22813\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__22816\,
            I => \ADC_VAC3.bit_cnt_4\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__22813\,
            I => \ADC_VAC3.bit_cnt_4\
        );

    \I__3392\ : InMux
    port map (
            O => \N__22808\,
            I => \ADC_VAC3.n13998\
        );

    \I__3391\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22801\
        );

    \I__3390\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22798\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__22801\,
            I => \ADC_VAC3.bit_cnt_5\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__22798\,
            I => \ADC_VAC3.bit_cnt_5\
        );

    \I__3387\ : InMux
    port map (
            O => \N__22793\,
            I => \ADC_VAC3.n13999\
        );

    \I__3386\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22786\
        );

    \I__3385\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22783\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__22786\,
            I => \ADC_VAC3.bit_cnt_6\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__22783\,
            I => \ADC_VAC3.bit_cnt_6\
        );

    \I__3382\ : InMux
    port map (
            O => \N__22778\,
            I => \ADC_VAC3.n14000\
        );

    \I__3381\ : InMux
    port map (
            O => \N__22775\,
            I => \ADC_VAC3.n14001\
        );

    \I__3380\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22768\
        );

    \I__3379\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22765\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__22768\,
            I => \ADC_VAC3.bit_cnt_7\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__22765\,
            I => \ADC_VAC3.bit_cnt_7\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__22760\,
            I => \N__22757\
        );

    \I__3375\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__22754\,
            I => \N__22750\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__22753\,
            I => \N__22747\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__22750\,
            I => \N__22744\
        );

    \I__3371\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22741\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__22744\,
            I => cmd_rdadctmp_31
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__22741\,
            I => cmd_rdadctmp_31
        );

    \I__3368\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22733\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__22733\,
            I => \N__22730\
        );

    \I__3366\ : Span12Mux_h
    port map (
            O => \N__22730\,
            I => \N__22726\
        );

    \I__3365\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22723\
        );

    \I__3364\ : Span12Mux_v
    port map (
            O => \N__22726\,
            I => \N__22720\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__22723\,
            I => buf_adcdata1_23
        );

    \I__3362\ : Odrv12
    port map (
            O => \N__22720\,
            I => buf_adcdata1_23
        );

    \I__3361\ : InMux
    port map (
            O => \N__22715\,
            I => \N__22712\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__22712\,
            I => \N__22707\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__22711\,
            I => \N__22704\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__22710\,
            I => \N__22701\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__22707\,
            I => \N__22698\
        );

    \I__3356\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22693\
        );

    \I__3355\ : InMux
    port map (
            O => \N__22701\,
            I => \N__22693\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__22698\,
            I => cmd_rdadctmp_23
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__22693\,
            I => cmd_rdadctmp_23
        );

    \I__3352\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22685\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22681\
        );

    \I__3350\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22678\
        );

    \I__3349\ : Span12Mux_s7_h
    port map (
            O => \N__22681\,
            I => \N__22675\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__22678\,
            I => buf_adcdata1_15
        );

    \I__3347\ : Odrv12
    port map (
            O => \N__22675\,
            I => buf_adcdata1_15
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__3345\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22663\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__22666\,
            I => \N__22660\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__22663\,
            I => \N__22657\
        );

    \I__3342\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22653\
        );

    \I__3341\ : Span4Mux_h
    port map (
            O => \N__22657\,
            I => \N__22650\
        );

    \I__3340\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22647\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__22653\,
            I => cmd_rdadctmp_20_adj_1129
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__22650\,
            I => cmd_rdadctmp_20_adj_1129
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__22647\,
            I => cmd_rdadctmp_20_adj_1129
        );

    \I__3336\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22636\
        );

    \I__3335\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22633\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__22636\,
            I => \ADC_VAC2.bit_cnt_4\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__22633\,
            I => \ADC_VAC2.bit_cnt_4\
        );

    \I__3332\ : InMux
    port map (
            O => \N__22628\,
            I => \N__22624\
        );

    \I__3331\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22621\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__22624\,
            I => \ADC_VAC2.bit_cnt_3\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__22621\,
            I => \ADC_VAC2.bit_cnt_3\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \N__22612\
        );

    \I__3327\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22609\
        );

    \I__3326\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22606\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__22609\,
            I => \ADC_VAC2.bit_cnt_5\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__22606\,
            I => \ADC_VAC2.bit_cnt_5\
        );

    \I__3323\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22597\
        );

    \I__3322\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22594\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__22597\,
            I => \ADC_VAC2.bit_cnt_2\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__22594\,
            I => \ADC_VAC2.bit_cnt_2\
        );

    \I__3319\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__22586\,
            I => \ADC_VAC2.n15596\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__22583\,
            I => \ADC_VAC3.n15334_cascade_\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__22580\,
            I => \ADC_VAC3.n15358_cascade_\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__22577\,
            I => \ADC_VAC3.n15602_cascade_\
        );

    \I__3314\ : CEMux
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__3312\ : Span4Mux_v
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__22562\,
            I => \ADC_VAC3.n15260\
        );

    \I__3309\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__22556\,
            I => \ADC_VAC3.n15259\
        );

    \I__3307\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__22544\,
            I => \ADC_VAC3.n17\
        );

    \I__3303\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__22535\,
            I => n8089
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__3299\ : InMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__22526\,
            I => \N__22523\
        );

    \I__3297\ : Odrv4
    port map (
            O => \N__22523\,
            I => n96_adj_1159
        );

    \I__3296\ : CascadeMux
    port map (
            O => \N__22520\,
            I => \n130_adj_1156_cascade_\
        );

    \I__3295\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22514\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__22514\,
            I => n15587
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__22511\,
            I => \n8051_cascade_\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__22508\,
            I => \N__22505\
        );

    \I__3291\ : InMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__22502\,
            I => \N__22497\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__22501\,
            I => \N__22494\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__22500\,
            I => \N__22491\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__22497\,
            I => \N__22488\
        );

    \I__3286\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22483\
        );

    \I__3285\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22483\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__22488\,
            I => cmd_rdadctmp_19_adj_1130
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__22483\,
            I => cmd_rdadctmp_19_adj_1130
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__22478\,
            I => \N__22473\
        );

    \I__3281\ : CascadeMux
    port map (
            O => \N__22477\,
            I => \N__22470\
        );

    \I__3280\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22467\
        );

    \I__3279\ : InMux
    port map (
            O => \N__22473\,
            I => \N__22464\
        );

    \I__3278\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22461\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__22467\,
            I => \N__22456\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__22464\,
            I => \N__22456\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__22461\,
            I => cmd_rdadctmp_8
        );

    \I__3274\ : Odrv12
    port map (
            O => \N__22456\,
            I => cmd_rdadctmp_8
        );

    \I__3273\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__3271\ : Sp12to4
    port map (
            O => \N__22445\,
            I => \N__22441\
        );

    \I__3270\ : InMux
    port map (
            O => \N__22444\,
            I => \N__22438\
        );

    \I__3269\ : Span12Mux_v
    port map (
            O => \N__22441\,
            I => \N__22435\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__22438\,
            I => buf_adcdata1_0
        );

    \I__3267\ : Odrv12
    port map (
            O => \N__22435\,
            I => buf_adcdata1_0
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__22430\,
            I => \n76_cascade_\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__22427\,
            I => \n4_adj_1195_cascade_\
        );

    \I__3264\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22421\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__22421\,
            I => n15632
        );

    \I__3262\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22415\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__22415\,
            I => n15589
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__22412\,
            I => \n87_adj_1165_cascade_\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__22409\,
            I => \n69_adj_1161_cascade_\
        );

    \I__3258\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__22403\,
            I => n130
        );

    \I__3256\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__22397\,
            I => n8050
        );

    \I__3254\ : SRMux
    port map (
            O => \N__22394\,
            I => \N__22389\
        );

    \I__3253\ : SRMux
    port map (
            O => \N__22393\,
            I => \N__22386\
        );

    \I__3252\ : SRMux
    port map (
            O => \N__22392\,
            I => \N__22380\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__22389\,
            I => \N__22377\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22374\
        );

    \I__3249\ : SRMux
    port map (
            O => \N__22385\,
            I => \N__22371\
        );

    \I__3248\ : SRMux
    port map (
            O => \N__22384\,
            I => \N__22367\
        );

    \I__3247\ : SRMux
    port map (
            O => \N__22383\,
            I => \N__22364\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__22380\,
            I => \N__22361\
        );

    \I__3245\ : Span4Mux_h
    port map (
            O => \N__22377\,
            I => \N__22358\
        );

    \I__3244\ : Span4Mux_h
    port map (
            O => \N__22374\,
            I => \N__22355\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__22371\,
            I => \N__22352\
        );

    \I__3242\ : SRMux
    port map (
            O => \N__22370\,
            I => \N__22349\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22343\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__22364\,
            I => \N__22343\
        );

    \I__3239\ : Span4Mux_h
    port map (
            O => \N__22361\,
            I => \N__22340\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__22358\,
            I => \N__22331\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__22355\,
            I => \N__22331\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__22352\,
            I => \N__22331\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22331\
        );

    \I__3234\ : SRMux
    port map (
            O => \N__22348\,
            I => \N__22328\
        );

    \I__3233\ : Span4Mux_h
    port map (
            O => \N__22343\,
            I => \N__22325\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__22340\,
            I => \N__22322\
        );

    \I__3231\ : Span4Mux_v
    port map (
            O => \N__22331\,
            I => \N__22319\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__22328\,
            I => \N__22316\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__22325\,
            I => n10660
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__22322\,
            I => n10660
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__22319\,
            I => n10660
        );

    \I__3226\ : Odrv12
    port map (
            O => \N__22316\,
            I => n10660
        );

    \I__3225\ : InMux
    port map (
            O => \N__22307\,
            I => \N__22304\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__22304\,
            I => comm_buf_7_4
        );

    \I__3223\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__22298\,
            I => \N__22295\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__22295\,
            I => comm_buf_11_4
        );

    \I__3220\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__22289\,
            I => comm_buf_9_4
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__22286\,
            I => \n16452_cascade_\
        );

    \I__3217\ : InMux
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__22280\,
            I => n16455
        );

    \I__3215\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22274\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__3213\ : Span4Mux_v
    port map (
            O => \N__22271\,
            I => \N__22268\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__22268\,
            I => \N__22265\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__22265\,
            I => comm_buf_5_4
        );

    \I__3210\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__22259\,
            I => \N__22256\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__22256\,
            I => comm_buf_4_4
        );

    \I__3207\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__22250\,
            I => n15400
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__22247\,
            I => \n15399_cascade_\
        );

    \I__3204\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22241\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__22241\,
            I => n16476
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__22238\,
            I => \n15633_cascade_\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__22235\,
            I => \n16458_cascade_\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__22232\,
            I => \n16461_cascade_\
        );

    \I__3199\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22226\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__22226\,
            I => \N__22223\
        );

    \I__3197\ : Span12Mux_h
    port map (
            O => \N__22223\,
            I => \N__22220\
        );

    \I__3196\ : Odrv12
    port map (
            O => \N__22220\,
            I => comm_buf_7_6
        );

    \I__3195\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22214\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__22214\,
            I => \N__22211\
        );

    \I__3193\ : Span12Mux_h
    port map (
            O => \N__22211\,
            I => \N__22208\
        );

    \I__3192\ : Odrv12
    port map (
            O => \N__22208\,
            I => buf_data3_13
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__22205\,
            I => \N__22202\
        );

    \I__3190\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22199\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__22199\,
            I => \N__22196\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__22193\,
            I => comm_buf_7_5
        );

    \I__3186\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__3184\ : Span4Mux_h
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__3183\ : Span4Mux_v
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__3181\ : Span4Mux_h
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__22172\,
            I => buf_data3_12
        );

    \I__3179\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__3176\ : Sp12to4
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__3175\ : Span12Mux_v
    port map (
            O => \N__22157\,
            I => \N__22154\
        );

    \I__3174\ : Odrv12
    port map (
            O => \N__22154\,
            I => buf_data3_11
        );

    \I__3173\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22148\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__22148\,
            I => \N__22145\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__22145\,
            I => comm_buf_7_3
        );

    \I__3170\ : InMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__22139\,
            I => \N__22136\
        );

    \I__3168\ : Span4Mux_v
    port map (
            O => \N__22136\,
            I => \N__22133\
        );

    \I__3167\ : Sp12to4
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__3166\ : Span12Mux_h
    port map (
            O => \N__22130\,
            I => \N__22127\
        );

    \I__3165\ : Span12Mux_v
    port map (
            O => \N__22127\,
            I => \N__22124\
        );

    \I__3164\ : Odrv12
    port map (
            O => \N__22124\,
            I => buf_data3_10
        );

    \I__3163\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__3161\ : Odrv12
    port map (
            O => \N__22115\,
            I => comm_buf_7_2
        );

    \I__3160\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__3158\ : Span4Mux_h
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__3157\ : Sp12to4
    port map (
            O => \N__22103\,
            I => \N__22100\
        );

    \I__3156\ : Span12Mux_v
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__3155\ : Span12Mux_h
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__3154\ : Odrv12
    port map (
            O => \N__22094\,
            I => buf_data3_9
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__3152\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__3150\ : Span4Mux_h
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__22079\,
            I => comm_buf_7_1
        );

    \I__3148\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__3146\ : Span4Mux_v
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__3145\ : Span4Mux_h
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__3144\ : Odrv4
    port map (
            O => \N__22064\,
            I => comm_buf_3_4
        );

    \I__3143\ : InMux
    port map (
            O => \N__22061\,
            I => \N__22058\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__3141\ : Span4Mux_v
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__22052\,
            I => comm_buf_2_4
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__22049\,
            I => \n15403_cascade_\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__22046\,
            I => \n16479_cascade_\
        );

    \I__3137\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__22040\,
            I => \N__22037\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__3134\ : Span4Mux_h
    port map (
            O => \N__22034\,
            I => \N__22031\
        );

    \I__3133\ : Sp12to4
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__3132\ : Odrv12
    port map (
            O => \N__22028\,
            I => buf_data4_3
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__3130\ : InMux
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__3128\ : Span4Mux_h
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__22013\,
            I => comm_buf_11_3
        );

    \I__3126\ : InMux
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__3124\ : Span4Mux_h
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__21998\,
            I => buf_data4_4
        );

    \I__3121\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21992\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__21989\,
            I => \N__21986\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__21986\,
            I => buf_data4_5
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__3116\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__21977\,
            I => comm_buf_11_5
        );

    \I__3114\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__3112\ : Span4Mux_h
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__3111\ : Span4Mux_h
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__21962\,
            I => buf_data4_6
        );

    \I__3109\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__21956\,
            I => \N__21953\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__21953\,
            I => \N__21950\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__21947\,
            I => buf_data4_7
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__3103\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__3101\ : Odrv4
    port map (
            O => \N__21935\,
            I => comm_buf_11_7
        );

    \I__3100\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__3097\ : Span4Mux_h
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__3096\ : Sp12to4
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__3095\ : Odrv12
    port map (
            O => \N__21917\,
            I => buf_data4_0
        );

    \I__3094\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__21911\,
            I => comm_buf_11_0
        );

    \I__3092\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__21896\,
            I => \N__21893\
        );

    \I__3087\ : Span4Mux_v
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__21890\,
            I => buf_data3_15
        );

    \I__3085\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__21881\,
            I => comm_buf_7_7
        );

    \I__3082\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__3080\ : Sp12to4
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__3079\ : Span12Mux_h
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__3078\ : Span12Mux_v
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__3077\ : Odrv12
    port map (
            O => \N__21863\,
            I => buf_data3_8
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__3075\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__21851\,
            I => comm_buf_7_0
        );

    \I__3072\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__3069\ : Span4Mux_v
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__3068\ : Span4Mux_h
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__3067\ : Span4Mux_h
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__21830\,
            I => buf_data3_14
        );

    \I__3065\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__21821\,
            I => comm_buf_3_7
        );

    \I__3062\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__3060\ : Span12Mux_h
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__3059\ : Odrv12
    port map (
            O => \N__21809\,
            I => comm_buf_2_7
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__21806\,
            I => \n15382_cascade_\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__21803\,
            I => \n16383_cascade_\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__21800\,
            I => \n16494_cascade_\
        );

    \I__3055\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__21794\,
            I => n16497
        );

    \I__3053\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__21788\,
            I => n15450
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__21785\,
            I => \n15451_cascade_\
        );

    \I__3050\ : InMux
    port map (
            O => \N__21782\,
            I => \N__21779\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__21779\,
            I => n16380
        );

    \I__3048\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__3046\ : Span12Mux_h
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__3045\ : Odrv12
    port map (
            O => \N__21767\,
            I => buf_data4_1
        );

    \I__3044\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21758\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__3041\ : Span4Mux_h
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__21749\,
            I => buf_data4_2
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__3037\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21740\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__21740\,
            I => \N__21737\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__21737\,
            I => comm_buf_11_2
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__3033\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__21728\,
            I => \N__21724\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__21727\,
            I => \N__21720\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__21724\,
            I => \N__21717\
        );

    \I__3029\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21712\
        );

    \I__3028\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21712\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__21717\,
            I => cmd_rdadctmp_14
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__21712\,
            I => cmd_rdadctmp_14
        );

    \I__3025\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21704\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__3022\ : Span4Mux_v
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__21695\,
            I => \N__21691\
        );

    \I__3020\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21688\
        );

    \I__3019\ : Span4Mux_h
    port map (
            O => \N__21691\,
            I => \N__21685\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__21688\,
            I => buf_adcdata1_6
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__21685\,
            I => buf_adcdata1_6
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__3015\ : InMux
    port map (
            O => \N__21677\,
            I => \N__21673\
        );

    \I__3014\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21670\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21667\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21664\
        );

    \I__3011\ : Span4Mux_h
    port map (
            O => \N__21667\,
            I => \N__21658\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__21664\,
            I => \N__21658\
        );

    \I__3009\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21655\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__21658\,
            I => cmd_rdadctmp_15_adj_1097
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__21655\,
            I => cmd_rdadctmp_15_adj_1097
        );

    \I__3006\ : IoInMux
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__3004\ : IoSpan4Mux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__3003\ : Span4Mux_s2_v
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__3002\ : Span4Mux_h
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__3001\ : Sp12to4
    port map (
            O => \N__21635\,
            I => \N__21631\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__21634\,
            I => \N__21628\
        );

    \I__2999\ : Span12Mux_s9_v
    port map (
            O => \N__21631\,
            I => \N__21625\
        );

    \I__2998\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21622\
        );

    \I__2997\ : Odrv12
    port map (
            O => \N__21625\,
            I => \M_SCLK4\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__21622\,
            I => \M_SCLK4\
        );

    \I__2995\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__21611\,
            I => \N__21607\
        );

    \I__2992\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21604\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__21607\,
            I => \comm_spi.n10434\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__21604\,
            I => \comm_spi.n10434\
        );

    \I__2989\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21594\
        );

    \I__2988\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21589\
        );

    \I__2987\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21589\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__21594\,
            I => \N__21586\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__21589\,
            I => comm_tx_buf_0
        );

    \I__2984\ : Odrv12
    port map (
            O => \N__21586\,
            I => comm_tx_buf_0
        );

    \I__2983\ : SRMux
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__21578\,
            I => \N__21575\
        );

    \I__2981\ : Odrv12
    port map (
            O => \N__21575\,
            I => \comm_spi.data_tx_7__N_834\
        );

    \I__2980\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21569\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__21569\,
            I => n16428
        );

    \I__2978\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__2976\ : Span12Mux_v
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__2975\ : Odrv12
    port map (
            O => \N__21557\,
            I => buf_data2_20
        );

    \I__2974\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21551\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__2972\ : Span4Mux_v
    port map (
            O => \N__21548\,
            I => \N__21545\
        );

    \I__2971\ : Odrv4
    port map (
            O => \N__21545\,
            I => n4104
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__21542\,
            I => \ADC_VAC2.n17_cascade_\
        );

    \I__2969\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21535\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__21538\,
            I => \N__21532\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__21535\,
            I => \N__21529\
        );

    \I__2966\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21526\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__21529\,
            I => cmd_rdadctmp_2_adj_1110
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__21526\,
            I => cmd_rdadctmp_2_adj_1110
        );

    \I__2963\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21517\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__21520\,
            I => \N__21514\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__21517\,
            I => \N__21511\
        );

    \I__2960\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21508\
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__21511\,
            I => cmd_rdadctmp_3_adj_1109
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__21508\,
            I => cmd_rdadctmp_3_adj_1109
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__21503\,
            I => \N__21499\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__21502\,
            I => \N__21496\
        );

    \I__2955\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21493\
        );

    \I__2954\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21490\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21487\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__21490\,
            I => acadc_dtrig2
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__21487\,
            I => acadc_dtrig2
        );

    \I__2950\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21478\
        );

    \I__2949\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21475\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__21478\,
            I => acadc_dtrig1
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__21475\,
            I => acadc_dtrig1
        );

    \I__2946\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21464\
        );

    \I__2945\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21464\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__21464\,
            I => acadc_dtrig4
        );

    \I__2943\ : InMux
    port map (
            O => \N__21461\,
            I => \N__21455\
        );

    \I__2942\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21455\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__21455\,
            I => acadc_dtrig3
        );

    \I__2940\ : InMux
    port map (
            O => \N__21452\,
            I => \ADC_VAC2.n13991\
        );

    \I__2939\ : InMux
    port map (
            O => \N__21449\,
            I => \ADC_VAC2.n13992\
        );

    \I__2938\ : InMux
    port map (
            O => \N__21446\,
            I => \ADC_VAC2.n13993\
        );

    \I__2937\ : InMux
    port map (
            O => \N__21443\,
            I => \ADC_VAC2.n13994\
        );

    \I__2936\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21436\
        );

    \I__2935\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21433\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__21436\,
            I => \ADC_VAC2.bit_cnt_1\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__21433\,
            I => \ADC_VAC2.bit_cnt_1\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__21428\,
            I => \N__21424\
        );

    \I__2931\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21421\
        );

    \I__2930\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21418\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__21421\,
            I => \ADC_VAC2.bit_cnt_7\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__21418\,
            I => \ADC_VAC2.bit_cnt_7\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__21413\,
            I => \ADC_VAC2.n15261_cascade_\
        );

    \I__2926\ : InMux
    port map (
            O => \N__21410\,
            I => \N__21407\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__21407\,
            I => \ADC_VAC2.n15595\
        );

    \I__2924\ : CEMux
    port map (
            O => \N__21404\,
            I => \N__21401\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__21401\,
            I => \ADC_VAC2.n15262\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__21398\,
            I => \N__21394\
        );

    \I__2921\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21391\
        );

    \I__2920\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21388\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__21391\,
            I => \ADC_VAC2.bit_cnt_6\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__21388\,
            I => \ADC_VAC2.bit_cnt_6\
        );

    \I__2917\ : InMux
    port map (
            O => \N__21383\,
            I => \N__21379\
        );

    \I__2916\ : InMux
    port map (
            O => \N__21382\,
            I => \N__21376\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__21379\,
            I => \ADC_VAC2.bit_cnt_0\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__21376\,
            I => \ADC_VAC2.bit_cnt_0\
        );

    \I__2913\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21368\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__21368\,
            I => \ADC_VAC2.n16\
        );

    \I__2911\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21362\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__21362\,
            I => \N__21359\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__21359\,
            I => \N__21356\
        );

    \I__2908\ : Sp12to4
    port map (
            O => \N__21356\,
            I => \N__21352\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__21355\,
            I => \N__21349\
        );

    \I__2906\ : Span12Mux_h
    port map (
            O => \N__21352\,
            I => \N__21346\
        );

    \I__2905\ : InMux
    port map (
            O => \N__21349\,
            I => \N__21343\
        );

    \I__2904\ : Span12Mux_v
    port map (
            O => \N__21346\,
            I => \N__21340\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__21343\,
            I => buf_adcdata1_22
        );

    \I__2902\ : Odrv12
    port map (
            O => \N__21340\,
            I => buf_adcdata1_22
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__21335\,
            I => \N__21332\
        );

    \I__2900\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21328\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__21331\,
            I => \N__21324\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21321\
        );

    \I__2897\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21318\
        );

    \I__2896\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21315\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__21321\,
            I => cmd_rdadctmp_24_adj_1052
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__21318\,
            I => cmd_rdadctmp_24_adj_1052
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__21315\,
            I => cmd_rdadctmp_24_adj_1052
        );

    \I__2892\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21305\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21301\
        );

    \I__2890\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__2889\ : Span12Mux_h
    port map (
            O => \N__21301\,
            I => \N__21295\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__21298\,
            I => buf_adcdata2_16
        );

    \I__2887\ : Odrv12
    port map (
            O => \N__21295\,
            I => buf_adcdata2_16
        );

    \I__2886\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21283\
        );

    \I__2885\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21283\
        );

    \I__2884\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21280\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__21283\,
            I => cmd_rdadctmp_29
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__21280\,
            I => cmd_rdadctmp_29
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__21275\,
            I => \N__21270\
        );

    \I__2880\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21263\
        );

    \I__2879\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21263\
        );

    \I__2878\ : InMux
    port map (
            O => \N__21270\,
            I => \N__21263\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__21263\,
            I => cmd_rdadctmp_30
        );

    \I__2876\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__2873\ : Sp12to4
    port map (
            O => \N__21251\,
            I => \N__21247\
        );

    \I__2872\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21244\
        );

    \I__2871\ : Span12Mux_v
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__21244\,
            I => buf_adcdata1_1
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__21241\,
            I => buf_adcdata1_1
        );

    \I__2868\ : InMux
    port map (
            O => \N__21236\,
            I => \bfn_9_13_0_\
        );

    \I__2867\ : InMux
    port map (
            O => \N__21233\,
            I => \ADC_VAC2.n13988\
        );

    \I__2866\ : InMux
    port map (
            O => \N__21230\,
            I => \ADC_VAC2.n13989\
        );

    \I__2865\ : InMux
    port map (
            O => \N__21227\,
            I => \ADC_VAC2.n13990\
        );

    \I__2864\ : IoInMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__2862\ : Span12Mux_s3_v
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__2861\ : Span12Mux_v
    port map (
            O => \N__21215\,
            I => \N__21211\
        );

    \I__2860\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21208\
        );

    \I__2859\ : Odrv12
    port map (
            O => \N__21211\,
            I => \DDS_MOSI1\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__21208\,
            I => \DDS_MOSI1\
        );

    \I__2857\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__21200\,
            I => n15522
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__2854\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__21191\,
            I => n15523
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__21188\,
            I => \n16398_cascade_\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__21185\,
            I => \n16401_cascade_\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__21182\,
            I => \n109_adj_1155_cascade_\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__21179\,
            I => \n8048_cascade_\
        );

    \I__2848\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__21170\,
            I => n15578
        );

    \I__2845\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__2843\ : Sp12to4
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__2842\ : Span12Mux_v
    port map (
            O => \N__21158\,
            I => \N__21154\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__21157\,
            I => \N__21151\
        );

    \I__2840\ : Span12Mux_v
    port map (
            O => \N__21154\,
            I => \N__21148\
        );

    \I__2839\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21145\
        );

    \I__2838\ : Span12Mux_h
    port map (
            O => \N__21148\,
            I => \N__21142\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__21145\,
            I => buf_adcdata1_21
        );

    \I__2836\ : Odrv12
    port map (
            O => \N__21142\,
            I => buf_adcdata1_21
        );

    \I__2835\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__21134\,
            I => \N__21131\
        );

    \I__2833\ : Span4Mux_v
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__21128\,
            I => \comm_buf_3_7_N_501_2\
        );

    \I__2831\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__2829\ : Odrv4
    port map (
            O => \N__21119\,
            I => comm_buf_3_2
        );

    \I__2828\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__21110\,
            I => \N__21107\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__21107\,
            I => comm_buf_3_3
        );

    \I__2824\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__2822\ : Span12Mux_h
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__2821\ : Odrv12
    port map (
            O => \N__21095\,
            I => buf_data4_19
        );

    \I__2820\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__2817\ : Sp12to4
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__2816\ : Odrv12
    port map (
            O => \N__21080\,
            I => comm_buf_9_3
        );

    \I__2815\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__21074\,
            I => \N__21071\
        );

    \I__2813\ : Span12Mux_v
    port map (
            O => \N__21071\,
            I => \N__21068\
        );

    \I__2812\ : Span12Mux_h
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__2811\ : Odrv12
    port map (
            O => \N__21065\,
            I => buf_data4_20
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__21062\,
            I => \n66_adj_1153_cascade_\
        );

    \I__2809\ : IoInMux
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__21053\
        );

    \I__2807\ : IoSpan4Mux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__2806\ : IoSpan4Mux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__2805\ : Sp12to4
    port map (
            O => \N__21047\,
            I => \N__21043\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__21046\,
            I => \N__21040\
        );

    \I__2803\ : Span12Mux_s7_v
    port map (
            O => \N__21043\,
            I => \N__21037\
        );

    \I__2802\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21034\
        );

    \I__2801\ : Odrv12
    port map (
            O => \N__21037\,
            I => \DDS_SCK1\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__21034\,
            I => \DDS_SCK1\
        );

    \I__2799\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21023\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__21023\,
            I => \N__21020\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__21020\,
            I => n16431
        );

    \I__2795\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21014\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__21008\,
            I => comm_buf_4_0
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__21005\,
            I => \n16506_cascade_\
        );

    \I__2790\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20999\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20996\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__20993\,
            I => comm_buf_5_0
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__2785\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__20984\,
            I => n16509
        );

    \I__2783\ : InMux
    port map (
            O => \N__20981\,
            I => \N__20978\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__20972\,
            I => n15424
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__2778\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20963\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__20963\,
            I => n15412
        );

    \I__2776\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20957\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__20957\,
            I => \N__20954\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__20954\,
            I => comm_buf_5_7
        );

    \I__2773\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__20948\,
            I => \N__20945\
        );

    \I__2771\ : Span4Mux_h
    port map (
            O => \N__20945\,
            I => \N__20942\
        );

    \I__2770\ : Odrv4
    port map (
            O => \N__20942\,
            I => comm_buf_4_7
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__20939\,
            I => \n16482_cascade_\
        );

    \I__2768\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20933\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__20933\,
            I => \N__20930\
        );

    \I__2766\ : Span4Mux_h
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__20927\,
            I => n16485
        );

    \I__2764\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20920\
        );

    \I__2763\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20917\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__20920\,
            I => \comm_spi.n16911\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__20917\,
            I => \comm_spi.n16911\
        );

    \I__2760\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20908\
        );

    \I__2759\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20905\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__20908\,
            I => \comm_spi.n10433\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__20905\,
            I => \comm_spi.n10433\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__20900\,
            I => \comm_spi.n16911_cascade_\
        );

    \I__2755\ : SRMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__2753\ : Span4Mux_v
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__20888\,
            I => \comm_spi.data_tx_7__N_811\
        );

    \I__2751\ : SRMux
    port map (
            O => \N__20885\,
            I => \N__20882\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__2749\ : Odrv12
    port map (
            O => \N__20879\,
            I => \comm_spi.data_tx_7__N_831\
        );

    \I__2748\ : SRMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__20873\,
            I => \comm_spi.data_tx_7__N_812\
        );

    \I__2746\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20861\
        );

    \I__2745\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20861\
        );

    \I__2744\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20861\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__2742\ : Span4Mux_v
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__20855\,
            I => comm_tx_buf_1
        );

    \I__2740\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20849\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__20849\,
            I => n15411
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__20846\,
            I => \n16446_cascade_\
        );

    \I__2737\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20840\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__20840\,
            I => n15391
        );

    \I__2735\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__20834\,
            I => n16449
        );

    \I__2733\ : InMux
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__2731\ : Span12Mux_h
    port map (
            O => \N__20825\,
            I => \N__20822\
        );

    \I__2730\ : Odrv12
    port map (
            O => \N__20822\,
            I => buf_data2_3
        );

    \I__2729\ : InMux
    port map (
            O => \N__20819\,
            I => \N__20815\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__20818\,
            I => \N__20812\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__20815\,
            I => \N__20808\
        );

    \I__2726\ : InMux
    port map (
            O => \N__20812\,
            I => \N__20805\
        );

    \I__2725\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20802\
        );

    \I__2724\ : Span12Mux_h
    port map (
            O => \N__20808\,
            I => \N__20797\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__20805\,
            I => \N__20797\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__20802\,
            I => buf_adcdata4_3
        );

    \I__2721\ : Odrv12
    port map (
            O => \N__20797\,
            I => buf_adcdata4_3
        );

    \I__2720\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20789\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__20789\,
            I => \N__20786\
        );

    \I__2718\ : Span4Mux_h
    port map (
            O => \N__20786\,
            I => \N__20783\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__20783\,
            I => n4305
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__2715\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__2713\ : Span4Mux_v
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__2712\ : Sp12to4
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__2711\ : Span12Mux_h
    port map (
            O => \N__20765\,
            I => \N__20762\
        );

    \I__2710\ : Odrv12
    port map (
            O => \N__20762\,
            I => \M_MISO3\
        );

    \I__2709\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20753\
        );

    \I__2708\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20753\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__20753\,
            I => cmd_rdadctmp_0_adj_1112
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__20750\,
            I => \N__20746\
        );

    \I__2705\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20743\
        );

    \I__2704\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20740\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__20743\,
            I => cmd_rdadctmp_1_adj_1111
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__20740\,
            I => cmd_rdadctmp_1_adj_1111
        );

    \I__2701\ : CEMux
    port map (
            O => \N__20735\,
            I => \N__20732\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__20729\,
            I => \N__20726\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__20726\,
            I => \ADC_VAC3.n12\
        );

    \I__2697\ : InMux
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__20717\,
            I => n15162
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__20714\,
            I => \n15162_cascade_\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__20711\,
            I => \n14_adj_1031_cascade_\
        );

    \I__2692\ : IoInMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__2690\ : Span4Mux_s0_v
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__2689\ : Sp12to4
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__2688\ : Span12Mux_s11_h
    port map (
            O => \N__20696\,
            I => \N__20692\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__20695\,
            I => \N__20689\
        );

    \I__2686\ : Span12Mux_v
    port map (
            O => \N__20692\,
            I => \N__20686\
        );

    \I__2685\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20683\
        );

    \I__2684\ : Odrv12
    port map (
            O => \N__20686\,
            I => \M_CS3\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__20683\,
            I => \M_CS3\
        );

    \I__2682\ : IoInMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__20675\,
            I => \N__20671\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__20674\,
            I => \N__20668\
        );

    \I__2679\ : Span12Mux_s11_v
    port map (
            O => \N__20671\,
            I => \N__20665\
        );

    \I__2678\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20662\
        );

    \I__2677\ : Odrv12
    port map (
            O => \N__20665\,
            I => \M_SCLK3\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__20662\,
            I => \M_SCLK3\
        );

    \I__2675\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20651\
        );

    \I__2674\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20651\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__20651\,
            I => cmd_rdadctmp_4_adj_1108
        );

    \I__2672\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__20645\,
            I => \N__20639\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__20644\,
            I => \N__20633\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__20643\,
            I => \N__20628\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__20642\,
            I => \N__20624\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__20639\,
            I => \N__20619\
        );

    \I__2666\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20612\
        );

    \I__2665\ : InMux
    port map (
            O => \N__20637\,
            I => \N__20612\
        );

    \I__2664\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20612\
        );

    \I__2663\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20605\
        );

    \I__2662\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20605\
        );

    \I__2661\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20605\
        );

    \I__2660\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20594\
        );

    \I__2659\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20594\
        );

    \I__2658\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20594\
        );

    \I__2657\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20594\
        );

    \I__2656\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20594\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__20619\,
            I => \DTRIG_N_957\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__20612\,
            I => \DTRIG_N_957\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__20605\,
            I => \DTRIG_N_957\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__20594\,
            I => \DTRIG_N_957\
        );

    \I__2651\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20582\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__20582\,
            I => \N__20577\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__20581\,
            I => \N__20570\
        );

    \I__2648\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20562\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__20577\,
            I => \N__20559\
        );

    \I__2646\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20552\
        );

    \I__2645\ : InMux
    port map (
            O => \N__20575\,
            I => \N__20552\
        );

    \I__2644\ : InMux
    port map (
            O => \N__20574\,
            I => \N__20552\
        );

    \I__2643\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20547\
        );

    \I__2642\ : InMux
    port map (
            O => \N__20570\,
            I => \N__20547\
        );

    \I__2641\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20536\
        );

    \I__2640\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20536\
        );

    \I__2639\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20536\
        );

    \I__2638\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20536\
        );

    \I__2637\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20536\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__20562\,
            I => adc_state_1
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__20559\,
            I => adc_state_1
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__20552\,
            I => adc_state_1
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__20547\,
            I => adc_state_1
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__20536\,
            I => adc_state_1
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__20525\,
            I => \N__20522\
        );

    \I__2630\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20519\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20515\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__20518\,
            I => \N__20511\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__20515\,
            I => \N__20508\
        );

    \I__2626\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20505\
        );

    \I__2625\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20502\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__20508\,
            I => cmd_rdadctmp_11
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__20505\,
            I => cmd_rdadctmp_11
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__20502\,
            I => cmd_rdadctmp_11
        );

    \I__2621\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20492\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20488\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__20491\,
            I => \N__20485\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__20488\,
            I => \N__20482\
        );

    \I__2617\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20478\
        );

    \I__2616\ : Sp12to4
    port map (
            O => \N__20482\,
            I => \N__20475\
        );

    \I__2615\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20472\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__20478\,
            I => \N__20469\
        );

    \I__2613\ : Span12Mux_h
    port map (
            O => \N__20475\,
            I => \N__20466\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__20472\,
            I => buf_adcdata4_12
        );

    \I__2611\ : Odrv12
    port map (
            O => \N__20469\,
            I => buf_adcdata4_12
        );

    \I__2610\ : Odrv12
    port map (
            O => \N__20466\,
            I => buf_adcdata4_12
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__20459\,
            I => \N__20455\
        );

    \I__2608\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__2607\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20446\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__20449\,
            I => \N__20442\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__20446\,
            I => \N__20439\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__20445\,
            I => \N__20436\
        );

    \I__2602\ : Span4Mux_h
    port map (
            O => \N__20442\,
            I => \N__20433\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__20439\,
            I => \N__20430\
        );

    \I__2600\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20427\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__20433\,
            I => cmd_rdadctmp_16_adj_1060
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__20430\,
            I => cmd_rdadctmp_16_adj_1060
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__20427\,
            I => cmd_rdadctmp_16_adj_1060
        );

    \I__2596\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__2593\ : Sp12to4
    port map (
            O => \N__20411\,
            I => \N__20407\
        );

    \I__2592\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20404\
        );

    \I__2591\ : Span12Mux_h
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__20404\,
            I => buf_adcdata2_8
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__20401\,
            I => buf_adcdata2_8
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20393\
        );

    \I__2587\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20388\
        );

    \I__2586\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20385\
        );

    \I__2585\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20382\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__20388\,
            I => cmd_rdadctmp_9_adj_1103
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__20385\,
            I => cmd_rdadctmp_9_adj_1103
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__20382\,
            I => cmd_rdadctmp_9_adj_1103
        );

    \I__2581\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20371\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__20374\,
            I => \N__20367\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__20371\,
            I => \N__20364\
        );

    \I__2578\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20359\
        );

    \I__2577\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20359\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__20364\,
            I => cmd_rdadctmp_28
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__20359\,
            I => cmd_rdadctmp_28
        );

    \I__2574\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__2572\ : Span4Mux_v
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__2571\ : Span4Mux_h
    port map (
            O => \N__20345\,
            I => \N__20341\
        );

    \I__2570\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20338\
        );

    \I__2569\ : Sp12to4
    port map (
            O => \N__20341\,
            I => \N__20335\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__20338\,
            I => buf_adcdata2_17
        );

    \I__2567\ : Odrv12
    port map (
            O => \N__20335\,
            I => buf_adcdata2_17
        );

    \I__2566\ : InMux
    port map (
            O => \N__20330\,
            I => \N__20327\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20323\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__20326\,
            I => \N__20319\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__20323\,
            I => \N__20316\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__20322\,
            I => \N__20313\
        );

    \I__2561\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20310\
        );

    \I__2560\ : Span4Mux_h
    port map (
            O => \N__20316\,
            I => \N__20307\
        );

    \I__2559\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20304\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__20310\,
            I => cmd_rdadctmp_13_adj_1099
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__20307\,
            I => cmd_rdadctmp_13_adj_1099
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__20304\,
            I => cmd_rdadctmp_13_adj_1099
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__20297\,
            I => \N__20293\
        );

    \I__2554\ : CascadeMux
    port map (
            O => \N__20296\,
            I => \N__20289\
        );

    \I__2553\ : InMux
    port map (
            O => \N__20293\,
            I => \N__20286\
        );

    \I__2552\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20281\
        );

    \I__2551\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20281\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__20286\,
            I => cmd_rdadctmp_14_adj_1098
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__20281\,
            I => cmd_rdadctmp_14_adj_1098
        );

    \I__2548\ : InMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__2546\ : Sp12to4
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__2545\ : Span12Mux_v
    port map (
            O => \N__20267\,
            I => \N__20264\
        );

    \I__2544\ : Span12Mux_h
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__2543\ : Odrv12
    port map (
            O => \N__20261\,
            I => buf_data2_14
        );

    \I__2542\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20255\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__20255\,
            I => \N__20252\
        );

    \I__2540\ : Odrv12
    port map (
            O => \N__20252\,
            I => n4058
        );

    \I__2539\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20240\
        );

    \I__2538\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20240\
        );

    \I__2537\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20240\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__20240\,
            I => cmd_rdadctmp_27
        );

    \I__2535\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__20234\,
            I => \N__20231\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__20228\,
            I => \N__20224\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__20227\,
            I => \N__20221\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__20224\,
            I => \N__20218\
        );

    \I__2529\ : InMux
    port map (
            O => \N__20221\,
            I => \N__20215\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__20218\,
            I => \N__20212\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__20215\,
            I => buf_adcdata1_19
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__20212\,
            I => buf_adcdata1_19
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__20207\,
            I => \N__20203\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__20206\,
            I => \N__20199\
        );

    \I__2523\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20192\
        );

    \I__2522\ : InMux
    port map (
            O => \N__20202\,
            I => \N__20192\
        );

    \I__2521\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20192\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__20192\,
            I => cmd_rdadctmp_25
        );

    \I__2519\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__2517\ : Span12Mux_v
    port map (
            O => \N__20183\,
            I => \N__20179\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__20182\,
            I => \N__20176\
        );

    \I__2515\ : Span12Mux_h
    port map (
            O => \N__20179\,
            I => \N__20173\
        );

    \I__2514\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20170\
        );

    \I__2513\ : Span12Mux_v
    port map (
            O => \N__20173\,
            I => \N__20167\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__20170\,
            I => buf_adcdata1_20
        );

    \I__2511\ : Odrv12
    port map (
            O => \N__20167\,
            I => buf_adcdata1_20
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__20162\,
            I => \n84_cascade_\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__20159\,
            I => \n15593_cascade_\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__20156\,
            I => \n8045_cascade_\
        );

    \I__2507\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__20150\,
            I => n15573
        );

    \I__2505\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20144\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__20141\,
            I => \N__20138\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__20138\,
            I => comm_buf_4_5
        );

    \I__2501\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__2499\ : Odrv12
    port map (
            O => \N__20129\,
            I => comm_buf_4_6
        );

    \I__2498\ : InMux
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__20123\,
            I => \N__20120\
        );

    \I__2496\ : Span4Mux_h
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__20111\,
            I => \N__20108\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__20108\,
            I => buf_data2_15
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__20105\,
            I => \n4057_cascade_\
        );

    \I__2490\ : SRMux
    port map (
            O => \N__20102\,
            I => \N__20099\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__20096\,
            I => \N__20092\
        );

    \I__2487\ : SRMux
    port map (
            O => \N__20095\,
            I => \N__20089\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__20092\,
            I => \N__20083\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__20089\,
            I => \N__20083\
        );

    \I__2484\ : SRMux
    port map (
            O => \N__20088\,
            I => \N__20080\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__20083\,
            I => \N__20077\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__20080\,
            I => \N__20074\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__20077\,
            I => n10604
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__20074\,
            I => n10604
        );

    \I__2479\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__20063\,
            I => \N__20060\
        );

    \I__2476\ : Span4Mux_h
    port map (
            O => \N__20060\,
            I => \N__20057\
        );

    \I__2475\ : Span4Mux_h
    port map (
            O => \N__20057\,
            I => \N__20053\
        );

    \I__2474\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20050\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__20053\,
            I => \N__20047\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__20050\,
            I => buf_adcdata1_17
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__20047\,
            I => buf_adcdata1_17
        );

    \I__2470\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20038\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__20041\,
            I => \N__20035\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__20038\,
            I => \N__20032\
        );

    \I__2467\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20029\
        );

    \I__2466\ : Span12Mux_h
    port map (
            O => \N__20032\,
            I => \N__20026\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20029\,
            I => buf_adcdata1_18
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__20026\,
            I => buf_adcdata1_18
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__20021\,
            I => \N__20016\
        );

    \I__2462\ : InMux
    port map (
            O => \N__20020\,
            I => \N__20009\
        );

    \I__2461\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20009\
        );

    \I__2460\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20009\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__20009\,
            I => cmd_rdadctmp_26
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__20006\,
            I => \n16407_cascade_\
        );

    \I__2457\ : InMux
    port map (
            O => \N__20003\,
            I => \N__20000\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__20000\,
            I => \N__19997\
        );

    \I__2455\ : Span4Mux_v
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__19994\,
            I => comm_buf_5_1
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__2452\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__19985\,
            I => \N__19982\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__19979\,
            I => comm_buf_4_1
        );

    \I__2448\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__19973\,
            I => n16515
        );

    \I__2446\ : InMux
    port map (
            O => \N__19970\,
            I => \N__19967\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__19967\,
            I => n16512
        );

    \I__2444\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__19961\,
            I => n7_adj_1240
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \n16425_cascade_\
        );

    \I__2441\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19949\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__2437\ : Span4Mux_h
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__2436\ : Sp12to4
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__2435\ : Odrv12
    port map (
            O => \N__19937\,
            I => buf_data2_12
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__19934\,
            I => \n4060_cascade_\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__19931\,
            I => \n16413_cascade_\
        );

    \I__2432\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19925\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__19922\,
            I => comm_buf_5_6
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__19919\,
            I => \n16518_cascade_\
        );

    \I__2428\ : InMux
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__19913\,
            I => n13493
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \n16521_cascade_\
        );

    \I__2425\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__19898\,
            I => comm_buf_2_6
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__19895\,
            I => \N__19892\
        );

    \I__2420\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__19889\,
            I => comm_buf_3_6
        );

    \I__2418\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__19883\,
            I => n16410
        );

    \I__2416\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19877\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__19877\,
            I => n16491
        );

    \I__2414\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19871\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19868\
        );

    \I__2412\ : Span4Mux_h
    port map (
            O => \N__19868\,
            I => \N__19865\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__19865\,
            I => comm_buf_2_1
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__19862\,
            I => \N__19859\
        );

    \I__2409\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__2407\ : Odrv12
    port map (
            O => \N__19853\,
            I => comm_buf_3_1
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__19850\,
            I => \n16404_cascade_\
        );

    \I__2405\ : InMux
    port map (
            O => \N__19847\,
            I => \N__19843\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__19846\,
            I => \N__19840\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19837\
        );

    \I__2402\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19834\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__19837\,
            I => cmd_rdadctmp_1_adj_1148
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__19834\,
            I => cmd_rdadctmp_1_adj_1148
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__2398\ : InMux
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__2395\ : Sp12to4
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__2394\ : Span12Mux_h
    port map (
            O => \N__19814\,
            I => \N__19811\
        );

    \I__2393\ : Span12Mux_h
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__2392\ : Odrv12
    port map (
            O => \N__19808\,
            I => \M_MISO4\
        );

    \I__2391\ : InMux
    port map (
            O => \N__19805\,
            I => \N__19801\
        );

    \I__2390\ : InMux
    port map (
            O => \N__19804\,
            I => \N__19798\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__19801\,
            I => cmd_rdadctmp_0_adj_1149
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__19798\,
            I => cmd_rdadctmp_0_adj_1149
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__2386\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__19784\,
            I => \N__19779\
        );

    \I__2383\ : InMux
    port map (
            O => \N__19783\,
            I => \N__19776\
        );

    \I__2382\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19773\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__19779\,
            I => cmd_rdadctmp_15
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__19776\,
            I => cmd_rdadctmp_15
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__19773\,
            I => cmd_rdadctmp_15
        );

    \I__2378\ : IoInMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__2376\ : IoSpan4Mux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__2375\ : Span4Mux_s1_v
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__19751\,
            I => \M_START\
        );

    \I__2372\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__19742\,
            I => comm_buf_3_0
        );

    \I__2369\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__19730\,
            I => comm_buf_2_0
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__19727\,
            I => \N__19723\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__19726\,
            I => \N__19719\
        );

    \I__2363\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19712\
        );

    \I__2362\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19712\
        );

    \I__2361\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19712\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__19712\,
            I => cmd_rdadctmp_18_adj_1131
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__19709\,
            I => \N__19705\
        );

    \I__2358\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19702\
        );

    \I__2357\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19699\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__19702\,
            I => \N__19696\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__19699\,
            I => \N__19692\
        );

    \I__2354\ : Span12Mux_v
    port map (
            O => \N__19696\,
            I => \N__19689\
        );

    \I__2353\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19686\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__19692\,
            I => \N__19683\
        );

    \I__2351\ : Span12Mux_h
    port map (
            O => \N__19689\,
            I => \N__19680\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__19686\,
            I => buf_adcdata4_10
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__19683\,
            I => buf_adcdata4_10
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__19680\,
            I => buf_adcdata4_10
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__19673\,
            I => \ADC_VAC1.n15263_cascade_\
        );

    \I__2346\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__19667\,
            I => \ADC_VAC1.n15553\
        );

    \I__2344\ : CEMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__19661\,
            I => \ADC_VAC1.n15264\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__19658\,
            I => \N__19654\
        );

    \I__2341\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19649\
        );

    \I__2340\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19649\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__19649\,
            I => \N__19644\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__19648\,
            I => \N__19641\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__19647\,
            I => \N__19637\
        );

    \I__2336\ : Span4Mux_v
    port map (
            O => \N__19644\,
            I => \N__19634\
        );

    \I__2335\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19631\
        );

    \I__2334\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19628\
        );

    \I__2333\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19625\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__19634\,
            I => \N__19622\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__19631\,
            I => \N__19615\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__19628\,
            I => \N__19615\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19615\
        );

    \I__2328\ : Sp12to4
    port map (
            O => \N__19622\,
            I => \N__19610\
        );

    \I__2327\ : Span12Mux_v
    port map (
            O => \N__19615\,
            I => \N__19610\
        );

    \I__2326\ : Odrv12
    port map (
            O => \N__19610\,
            I => \M_DRDY1\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__19607\,
            I => \ADC_VAC1.n17_cascade_\
        );

    \I__2324\ : CEMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__19598\,
            I => \ADC_VAC1.n12\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__19595\,
            I => \N__19592\
        );

    \I__2320\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19587\
        );

    \I__2319\ : InMux
    port map (
            O => \N__19591\,
            I => \N__19584\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__19590\,
            I => \N__19581\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19578\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__19584\,
            I => \N__19575\
        );

    \I__2315\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19572\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__19578\,
            I => cmd_rdadctmp_13
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__19575\,
            I => cmd_rdadctmp_13
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__19572\,
            I => cmd_rdadctmp_13
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__19565\,
            I => \N__19561\
        );

    \I__2310\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19558\
        );

    \I__2309\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19555\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__19558\,
            I => \N__19552\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__19555\,
            I => \N__19548\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__19552\,
            I => \N__19545\
        );

    \I__2305\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19542\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__19548\,
            I => \N__19539\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__19545\,
            I => \N__19536\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__19542\,
            I => buf_adcdata3_5
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__19539\,
            I => buf_adcdata3_5
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__19536\,
            I => buf_adcdata3_5
        );

    \I__2299\ : InMux
    port map (
            O => \N__19529\,
            I => \N__19525\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__19528\,
            I => \N__19522\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__19525\,
            I => \N__19519\
        );

    \I__2296\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19516\
        );

    \I__2295\ : Span4Mux_h
    port map (
            O => \N__19519\,
            I => \N__19512\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19509\
        );

    \I__2293\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19506\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19503\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__19509\,
            I => \N__19500\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__19506\,
            I => buf_adcdata3_6
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__19503\,
            I => buf_adcdata3_6
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__19500\,
            I => buf_adcdata3_6
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__19493\,
            I => \N__19489\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__19492\,
            I => \N__19485\
        );

    \I__2285\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19480\
        );

    \I__2284\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19480\
        );

    \I__2283\ : InMux
    port map (
            O => \N__19485\,
            I => \N__19477\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__19480\,
            I => cmd_rdadctmp_12
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__19477\,
            I => cmd_rdadctmp_12
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__19472\,
            I => \N__19467\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__19471\,
            I => \N__19464\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__19470\,
            I => \N__19461\
        );

    \I__2277\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19456\
        );

    \I__2276\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19456\
        );

    \I__2275\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19453\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__19456\,
            I => cmd_rdadctmp_10_adj_1102
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__19453\,
            I => cmd_rdadctmp_10_adj_1102
        );

    \I__2272\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19442\
        );

    \I__2271\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19442\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19438\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__2267\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__19432\,
            I => cmd_rdadctmp_16_adj_1133
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__19429\,
            I => cmd_rdadctmp_16_adj_1133
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__19424\,
            I => \N__19419\
        );

    \I__2263\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19412\
        );

    \I__2262\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19412\
        );

    \I__2261\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19412\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__19412\,
            I => cmd_rdadctmp_17_adj_1132
        );

    \I__2259\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__19406\,
            I => comm_buf_4_3
        );

    \I__2257\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__19394\,
            I => comm_buf_5_3
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__19391\,
            I => \n16440_cascade_\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__2251\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19382\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__19382\,
            I => n15423
        );

    \I__2249\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__19376\,
            I => n15397
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__19373\,
            I => \n16392_cascade_\
        );

    \I__2246\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19367\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__19367\,
            I => n16443
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__19364\,
            I => \n16395_cascade_\
        );

    \I__2243\ : IoInMux
    port map (
            O => \N__19361\,
            I => \N__19358\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__2241\ : IoSpan4Mux
    port map (
            O => \N__19355\,
            I => \N__19352\
        );

    \I__2240\ : Span4Mux_s2_h
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__2239\ : Sp12to4
    port map (
            O => \N__19349\,
            I => \N__19345\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__19348\,
            I => \N__19342\
        );

    \I__2237\ : Span12Mux_v
    port map (
            O => \N__19345\,
            I => \N__19339\
        );

    \I__2236\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19336\
        );

    \I__2235\ : Odrv12
    port map (
            O => \N__19339\,
            I => \M_SCLK2\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__19336\,
            I => \M_SCLK2\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__19331\,
            I => \n15388_cascade_\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__19328\,
            I => \n16389_cascade_\
        );

    \I__2231\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__19322\,
            I => comm_buf_4_2
        );

    \I__2229\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19316\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19313\
        );

    \I__2227\ : Odrv12
    port map (
            O => \N__19313\,
            I => comm_buf_5_2
        );

    \I__2226\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19307\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__19307\,
            I => n15448
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__19304\,
            I => \n15447_cascade_\
        );

    \I__2223\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19298\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__19298\,
            I => n16386
        );

    \I__2221\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__19292\,
            I => \N__19289\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__19289\,
            I => \N__19286\
        );

    \I__2218\ : Span4Mux_h
    port map (
            O => \N__19286\,
            I => \N__19282\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__19285\,
            I => \N__19279\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__19282\,
            I => \N__19275\
        );

    \I__2215\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19272\
        );

    \I__2214\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19269\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__19275\,
            I => \N__19264\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__19272\,
            I => \N__19264\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__19269\,
            I => buf_adcdata4_18
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__19264\,
            I => buf_adcdata4_18
        );

    \I__2209\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19256\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__19250\,
            I => comm_buf_2_3
        );

    \I__2205\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19244\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__19244\,
            I => \N__19241\
        );

    \I__2203\ : Span4Mux_h
    port map (
            O => \N__19241\,
            I => \N__19238\
        );

    \I__2202\ : Span4Mux_v
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__19229\,
            I => buf_data2_17
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__19226\,
            I => \n4107_cascade_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__19217\,
            I => \N__19214\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__19211\,
            I => \N__19208\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__19205\,
            I => buf_data2_18
        );

    \I__2190\ : CEMux
    port map (
            O => \N__19202\,
            I => \N__19198\
        );

    \I__2189\ : CEMux
    port map (
            O => \N__19201\,
            I => \N__19195\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__19198\,
            I => \N__19192\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__19195\,
            I => \N__19189\
        );

    \I__2186\ : Span4Mux_v
    port map (
            O => \N__19192\,
            I => \N__19186\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__19189\,
            I => \N__19183\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__19186\,
            I => n8787
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__19183\,
            I => n8787
        );

    \I__2182\ : SRMux
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__19175\,
            I => \N__19171\
        );

    \I__2180\ : SRMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__19171\,
            I => \N__19165\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__19168\,
            I => \N__19162\
        );

    \I__2177\ : Span4Mux_h
    port map (
            O => \N__19165\,
            I => \N__19157\
        );

    \I__2176\ : Span4Mux_v
    port map (
            O => \N__19162\,
            I => \N__19157\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__19157\,
            I => n10599
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__2173\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__19148\,
            I => comm_buf_2_2
        );

    \I__2171\ : InMux
    port map (
            O => \N__19145\,
            I => \ADC_VAC1.n13987\
        );

    \I__2170\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19138\
        );

    \I__2169\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19135\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__19138\,
            I => \ADC_VAC1.bit_cnt_7\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__19135\,
            I => \ADC_VAC1.bit_cnt_7\
        );

    \I__2166\ : CEMux
    port map (
            O => \N__19130\,
            I => \N__19127\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__19124\,
            I => \ADC_VAC1.n9312\
        );

    \I__2163\ : SRMux
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__19118\,
            I => \ADC_VAC1.n10667\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__19115\,
            I => \n16470_cascade_\
        );

    \I__2160\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__19109\,
            I => \N__19106\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__19103\,
            I => comm_buf_5_5
        );

    \I__2156\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19097\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__19097\,
            I => \N__19094\
        );

    \I__2154\ : Span4Mux_h
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__19091\,
            I => comm_buf_2_5
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \n16416_cascade_\
        );

    \I__2151\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19082\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__19082\,
            I => n16473
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__19079\,
            I => \n16419_cascade_\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \n7_adj_1238_cascade_\
        );

    \I__2147\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__2145\ : Span4Mux_v
    port map (
            O => \N__19067\,
            I => \N__19064\
        );

    \I__2144\ : Sp12to4
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__2143\ : Span12Mux_h
    port map (
            O => \N__19061\,
            I => \N__19058\
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__19058\,
            I => buf_data2_21
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__19055\,
            I => \n4103_cascade_\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__19052\,
            I => \N__19049\
        );

    \I__2139\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__19046\,
            I => comm_buf_3_5
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__19043\,
            I => \ADC_VAC1.n15360_cascade_\
        );

    \I__2136\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19036\
        );

    \I__2135\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19033\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__19036\,
            I => \ADC_VAC1.bit_cnt_0\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__19033\,
            I => \ADC_VAC1.bit_cnt_0\
        );

    \I__2132\ : InMux
    port map (
            O => \N__19028\,
            I => \bfn_6_16_0_\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__19025\,
            I => \N__19021\
        );

    \I__2130\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19018\
        );

    \I__2129\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19015\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__19018\,
            I => \ADC_VAC1.bit_cnt_1\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__19015\,
            I => \ADC_VAC1.bit_cnt_1\
        );

    \I__2126\ : InMux
    port map (
            O => \N__19010\,
            I => \ADC_VAC1.n13981\
        );

    \I__2125\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19003\
        );

    \I__2124\ : InMux
    port map (
            O => \N__19006\,
            I => \N__19000\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__19003\,
            I => \ADC_VAC1.bit_cnt_2\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__19000\,
            I => \ADC_VAC1.bit_cnt_2\
        );

    \I__2121\ : InMux
    port map (
            O => \N__18995\,
            I => \ADC_VAC1.n13982\
        );

    \I__2120\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18988\
        );

    \I__2119\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__18988\,
            I => \ADC_VAC1.bit_cnt_3\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__18985\,
            I => \ADC_VAC1.bit_cnt_3\
        );

    \I__2116\ : InMux
    port map (
            O => \N__18980\,
            I => \ADC_VAC1.n13983\
        );

    \I__2115\ : InMux
    port map (
            O => \N__18977\,
            I => \N__18973\
        );

    \I__2114\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18970\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__18973\,
            I => \ADC_VAC1.bit_cnt_4\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__18970\,
            I => \ADC_VAC1.bit_cnt_4\
        );

    \I__2111\ : InMux
    port map (
            O => \N__18965\,
            I => \ADC_VAC1.n13984\
        );

    \I__2110\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18958\
        );

    \I__2109\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18955\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__18958\,
            I => \N__18952\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__18955\,
            I => \ADC_VAC1.bit_cnt_5\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__18952\,
            I => \ADC_VAC1.bit_cnt_5\
        );

    \I__2105\ : InMux
    port map (
            O => \N__18947\,
            I => \ADC_VAC1.n13985\
        );

    \I__2104\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18940\
        );

    \I__2103\ : InMux
    port map (
            O => \N__18943\,
            I => \N__18937\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__18940\,
            I => \ADC_VAC1.bit_cnt_6\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__18937\,
            I => \ADC_VAC1.bit_cnt_6\
        );

    \I__2100\ : InMux
    port map (
            O => \N__18932\,
            I => \ADC_VAC1.n13986\
        );

    \I__2099\ : InMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__18926\,
            I => n15168
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__18923\,
            I => \n15168_cascade_\
        );

    \I__2096\ : IoInMux
    port map (
            O => \N__18920\,
            I => \N__18917\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__18917\,
            I => \N__18914\
        );

    \I__2094\ : IoSpan4Mux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__2093\ : Span4Mux_s3_h
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__2092\ : Span4Mux_h
    port map (
            O => \N__18908\,
            I => \N__18904\
        );

    \I__2091\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__18904\,
            I => \M_CS1\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__18901\,
            I => \M_CS1\
        );

    \I__2088\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__18893\,
            I => n14_adj_1039
        );

    \I__2086\ : IoInMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__2084\ : IoSpan4Mux
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__2083\ : Span4Mux_s3_h
    port map (
            O => \N__18881\,
            I => \N__18877\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__18880\,
            I => \N__18874\
        );

    \I__2081\ : Span4Mux_h
    port map (
            O => \N__18877\,
            I => \N__18871\
        );

    \I__2080\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18868\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__18871\,
            I => \M_SCLK1\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__18868\,
            I => \M_SCLK1\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__18863\,
            I => \ADC_VAC1.n9312_cascade_\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__18860\,
            I => \ADC_VAC1.n15338_cascade_\
        );

    \I__2075\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18853\
        );

    \I__2074\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__18853\,
            I => cmd_rdadctmp_2
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__18850\,
            I => cmd_rdadctmp_2
        );

    \I__2071\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18839\
        );

    \I__2070\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18839\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__18839\,
            I => cmd_rdadctmp_7
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__2067\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18827\
        );

    \I__2066\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18827\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__18827\,
            I => cmd_rdadctmp_6
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__2063\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18815\
        );

    \I__2062\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18815\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__18815\,
            I => cmd_rdadctmp_5
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \N__18808\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__18811\,
            I => \N__18805\
        );

    \I__2058\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18800\
        );

    \I__2057\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18800\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__18800\,
            I => cmd_rdadctmp_3
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__2054\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18788\
        );

    \I__2053\ : InMux
    port map (
            O => \N__18793\,
            I => \N__18788\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__18788\,
            I => cmd_rdadctmp_4
        );

    \I__2051\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__2049\ : Span12Mux_s10_h
    port map (
            O => \N__18779\,
            I => \N__18775\
        );

    \I__2048\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__2047\ : Span12Mux_h
    port map (
            O => \N__18775\,
            I => \N__18769\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__18772\,
            I => buf_adcdata1_3
        );

    \I__2045\ : Odrv12
    port map (
            O => \N__18769\,
            I => buf_adcdata1_3
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__18764\,
            I => \N__18761\
        );

    \I__2043\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18757\
        );

    \I__2042\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18754\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__18757\,
            I => \N__18750\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__18754\,
            I => \N__18747\
        );

    \I__2039\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18744\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__18750\,
            I => \N__18739\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__18747\,
            I => \N__18739\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__18744\,
            I => buf_adcdata3_4
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__18739\,
            I => buf_adcdata3_4
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__18734\,
            I => \N__18730\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__18733\,
            I => \N__18727\
        );

    \I__2032\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18722\
        );

    \I__2031\ : InMux
    port map (
            O => \N__18727\,
            I => \N__18722\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__18722\,
            I => cmd_rdadctmp_1
        );

    \I__2029\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18716\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__18716\,
            I => \N__18712\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__18715\,
            I => \N__18709\
        );

    \I__2026\ : Span4Mux_h
    port map (
            O => \N__18712\,
            I => \N__18705\
        );

    \I__2025\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18702\
        );

    \I__2024\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18699\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__18705\,
            I => \N__18696\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__18702\,
            I => \N__18693\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__18699\,
            I => buf_adcdata3_7
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__18696\,
            I => buf_adcdata3_7
        );

    \I__2019\ : Odrv12
    port map (
            O => \N__18693\,
            I => buf_adcdata3_7
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__2017\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18680\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__2014\ : Span4Mux_h
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__18671\,
            I => \N__18668\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__18668\,
            I => \M_MISO1\
        );

    \I__2011\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18659\
        );

    \I__2010\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18659\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__18659\,
            I => cmd_rdadctmp_0
        );

    \I__2008\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18652\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18649\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__18652\,
            I => \N__18645\
        );

    \I__2005\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18640\
        );

    \I__2004\ : InMux
    port map (
            O => \N__18648\,
            I => \N__18640\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__18645\,
            I => cmd_rdadctmp_12_adj_1100
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__18640\,
            I => cmd_rdadctmp_12_adj_1100
        );

    \I__2001\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__18629\,
            I => \N__18625\
        );

    \I__1998\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18622\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__18625\,
            I => \N__18619\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__18622\,
            I => buf_adcdata1_4
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__18619\,
            I => buf_adcdata1_4
        );

    \I__1994\ : SRMux
    port map (
            O => \N__18614\,
            I => \N__18609\
        );

    \I__1993\ : SRMux
    port map (
            O => \N__18613\,
            I => \N__18606\
        );

    \I__1992\ : SRMux
    port map (
            O => \N__18612\,
            I => \N__18603\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__18609\,
            I => \N__18600\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18597\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__18603\,
            I => \N__18594\
        );

    \I__1988\ : Span4Mux_h
    port map (
            O => \N__18600\,
            I => \N__18591\
        );

    \I__1987\ : Odrv12
    port map (
            O => \N__18597\,
            I => n10590
        );

    \I__1986\ : Odrv12
    port map (
            O => \N__18594\,
            I => n10590
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__18591\,
            I => n10590
        );

    \I__1984\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18580\
        );

    \I__1983\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18577\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__18580\,
            I => \N__18574\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__18577\,
            I => secclk_cnt_21
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__18574\,
            I => secclk_cnt_21
        );

    \I__1979\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18565\
        );

    \I__1978\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18562\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__18565\,
            I => \N__18559\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__18562\,
            I => secclk_cnt_19
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__18559\,
            I => secclk_cnt_19
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__1973\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__18548\,
            I => \N__18544\
        );

    \I__1971\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18541\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__18544\,
            I => \N__18538\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__18541\,
            I => secclk_cnt_12
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__18538\,
            I => secclk_cnt_12
        );

    \I__1967\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18529\
        );

    \I__1966\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18526\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__18529\,
            I => \N__18523\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__18526\,
            I => secclk_cnt_22
        );

    \I__1963\ : Odrv12
    port map (
            O => \N__18523\,
            I => secclk_cnt_22
        );

    \I__1962\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__1960\ : Span12Mux_v
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__18509\,
            I => n14_adj_1163
        );

    \I__1958\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__1954\ : Sp12to4
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__1953\ : Span12Mux_v
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__1952\ : Odrv12
    port map (
            O => \N__18488\,
            I => buf_data2_10
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__18485\,
            I => \n4062_cascade_\
        );

    \I__1950\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__1948\ : Span4Mux_v
    port map (
            O => \N__18476\,
            I => \N__18472\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__18475\,
            I => \N__18469\
        );

    \I__1946\ : Span4Mux_h
    port map (
            O => \N__18472\,
            I => \N__18466\
        );

    \I__1945\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18463\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__18466\,
            I => \N__18460\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__18463\,
            I => \N__18454\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__1941\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18451\
        );

    \I__1940\ : Span4Mux_h
    port map (
            O => \N__18454\,
            I => \N__18448\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__18451\,
            I => buf_adcdata3_2
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__18448\,
            I => buf_adcdata3_2
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__18443\,
            I => \N__18439\
        );

    \I__1936\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18431\
        );

    \I__1935\ : InMux
    port map (
            O => \N__18439\,
            I => \N__18431\
        );

    \I__1934\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18431\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__18431\,
            I => cmd_rdadctmp_11_adj_1101
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__18428\,
            I => \n8787_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__1929\ : Span4Mux_v
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__1928\ : Sp12to4
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__1927\ : Span12Mux_h
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__1926\ : Odrv12
    port map (
            O => \N__18410\,
            I => buf_data1_2
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \n4150_cascade_\
        );

    \I__1924\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__1922\ : Odrv12
    port map (
            O => \N__18398\,
            I => buf_data1_4
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__18395\,
            I => \n4148_cascade_\
        );

    \I__1920\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__1918\ : Span4Mux_h
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__18383\,
            I => buf_data1_5
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__18380\,
            I => \n4147_cascade_\
        );

    \I__1915\ : CEMux
    port map (
            O => \N__18377\,
            I => \N__18372\
        );

    \I__1914\ : CEMux
    port map (
            O => \N__18376\,
            I => \N__18369\
        );

    \I__1913\ : CEMux
    port map (
            O => \N__18375\,
            I => \N__18366\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__18372\,
            I => n8738
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__18369\,
            I => n8738
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__18366\,
            I => n8738
        );

    \I__1909\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18356\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__18353\,
            I => buf_data1_7
        );

    \I__1906\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__18344\,
            I => n4145
        );

    \I__1903\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18338\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__18338\,
            I => n4152
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \n15131_cascade_\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__18332\,
            I => \n8738_cascade_\
        );

    \I__1899\ : CEMux
    port map (
            O => \N__18329\,
            I => \N__18326\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__18326\,
            I => \N__18322\
        );

    \I__1897\ : CEMux
    port map (
            O => \N__18325\,
            I => \N__18319\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__18322\,
            I => \N__18316\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18313\
        );

    \I__1894\ : Span4Mux_h
    port map (
            O => \N__18316\,
            I => \N__18310\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__18313\,
            I => \N__18307\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__18310\,
            I => n8847
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__18307\,
            I => n8847
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \n8847_cascade_\
        );

    \I__1889\ : SRMux
    port map (
            O => \N__18299\,
            I => \N__18295\
        );

    \I__1888\ : SRMux
    port map (
            O => \N__18298\,
            I => \N__18292\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__18295\,
            I => n10611
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__18292\,
            I => n10611
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__1884\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18278\
        );

    \I__1883\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18278\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__18278\,
            I => cmd_rdadctmp_7_adj_1142
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__18275\,
            I => \N__18271\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__1879\ : InMux
    port map (
            O => \N__18271\,
            I => \N__18262\
        );

    \I__1878\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__1877\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18259\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__18262\,
            I => cmd_rdadctmp_8_adj_1141
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__18259\,
            I => cmd_rdadctmp_8_adj_1141
        );

    \I__1874\ : InMux
    port map (
            O => \N__18254\,
            I => \N__18250\
        );

    \I__1873\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18247\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__18250\,
            I => cmd_rdadctmp_5_adj_1144
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__18247\,
            I => cmd_rdadctmp_5_adj_1144
        );

    \I__1870\ : InMux
    port map (
            O => \N__18242\,
            I => \N__18236\
        );

    \I__1869\ : InMux
    port map (
            O => \N__18241\,
            I => \N__18236\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__18236\,
            I => cmd_rdadctmp_6_adj_1143
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__18233\,
            I => \N__18230\
        );

    \I__1866\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18227\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18224\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__18224\,
            I => \N__18221\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__18221\,
            I => \N__18216\
        );

    \I__1862\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18213\
        );

    \I__1861\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18210\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__18216\,
            I => cmd_rdadctmp_11_adj_1138
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__18213\,
            I => cmd_rdadctmp_11_adj_1138
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__18210\,
            I => cmd_rdadctmp_11_adj_1138
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__18203\,
            I => \N__18199\
        );

    \I__1856\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18196\
        );

    \I__1855\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18193\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__18196\,
            I => cmd_rdadctmp_4_adj_1145
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__18193\,
            I => cmd_rdadctmp_4_adj_1145
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__18188\,
            I => \N__18184\
        );

    \I__1851\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18179\
        );

    \I__1850\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18179\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__18179\,
            I => cmd_rdadctmp_3_adj_1146
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__18176\,
            I => \N__18172\
        );

    \I__1847\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18169\
        );

    \I__1846\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18166\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__18169\,
            I => cmd_rdadctmp_2_adj_1147
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__18166\,
            I => cmd_rdadctmp_2_adj_1147
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__1842\ : InMux
    port map (
            O => \N__18158\,
            I => \N__18155\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__18152\,
            I => \N__18147\
        );

    \I__1839\ : InMux
    port map (
            O => \N__18151\,
            I => \N__18144\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__18150\,
            I => \N__18141\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__18147\,
            I => \N__18138\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18135\
        );

    \I__1835\ : InMux
    port map (
            O => \N__18141\,
            I => \N__18132\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__18138\,
            I => cmd_rdadctmp_12_adj_1137
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__18135\,
            I => cmd_rdadctmp_12_adj_1137
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__18132\,
            I => cmd_rdadctmp_12_adj_1137
        );

    \I__1831\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18117\
        );

    \I__1829\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18114\
        );

    \I__1828\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18111\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__18117\,
            I => \N__18108\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__18114\,
            I => buf_adcdata4_4
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__18111\,
            I => buf_adcdata4_4
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__18108\,
            I => buf_adcdata4_4
        );

    \I__1823\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__18092\,
            I => buf_data1_6
        );

    \I__1819\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__18080\,
            I => n4146
        );

    \I__1815\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__1813\ : Span4Mux_h
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__1812\ : Sp12to4
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__1811\ : Span12Mux_h
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__1810\ : Odrv12
    port map (
            O => \N__18062\,
            I => buf_data1_0
        );

    \I__1809\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__18056\,
            I => \N__18051\
        );

    \I__1807\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18048\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__18054\,
            I => \N__18045\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__18051\,
            I => \N__18042\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__18048\,
            I => \N__18039\
        );

    \I__1803\ : InMux
    port map (
            O => \N__18045\,
            I => \N__18036\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__18042\,
            I => cmd_rdadctmp_15_adj_1134
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__18039\,
            I => cmd_rdadctmp_15_adj_1134
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__18036\,
            I => cmd_rdadctmp_15_adj_1134
        );

    \I__1799\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18026\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18026\,
            I => \N__18023\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__1795\ : Sp12to4
    port map (
            O => \N__18017\,
            I => \N__18012\
        );

    \I__1794\ : InMux
    port map (
            O => \N__18016\,
            I => \N__18009\
        );

    \I__1793\ : InMux
    port map (
            O => \N__18015\,
            I => \N__18006\
        );

    \I__1792\ : Span12Mux_h
    port map (
            O => \N__18012\,
            I => \N__18003\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__18009\,
            I => \N__18000\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__18006\,
            I => buf_adcdata4_0
        );

    \I__1789\ : Odrv12
    port map (
            O => \N__18003\,
            I => buf_adcdata4_0
        );

    \I__1788\ : Odrv12
    port map (
            O => \N__18000\,
            I => buf_adcdata4_0
        );

    \I__1787\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__17987\,
            I => \N__17983\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__17986\,
            I => \N__17980\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__17983\,
            I => \N__17977\
        );

    \I__1782\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17973\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__17977\,
            I => \N__17970\
        );

    \I__1780\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17967\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__17973\,
            I => \N__17964\
        );

    \I__1778\ : Span12Mux_h
    port map (
            O => \N__17970\,
            I => \N__17961\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__17967\,
            I => buf_adcdata4_1
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__17964\,
            I => buf_adcdata4_1
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__17961\,
            I => buf_adcdata4_1
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__17954\,
            I => \N__17950\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__17953\,
            I => \N__17947\
        );

    \I__1772\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17939\
        );

    \I__1771\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17939\
        );

    \I__1770\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17939\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__17939\,
            I => cmd_rdadctmp_9_adj_1140
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__17936\,
            I => \N__17932\
        );

    \I__1767\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17924\
        );

    \I__1766\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17924\
        );

    \I__1765\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17924\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__17924\,
            I => cmd_rdadctmp_10_adj_1139
        );

    \I__1763\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17918\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__17918\,
            I => \N__17915\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__17915\,
            I => \N__17911\
        );

    \I__1760\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17907\
        );

    \I__1759\ : Sp12to4
    port map (
            O => \N__17911\,
            I => \N__17904\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__17910\,
            I => \N__17901\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__17907\,
            I => \N__17896\
        );

    \I__1756\ : Span12Mux_s11_h
    port map (
            O => \N__17904\,
            I => \N__17896\
        );

    \I__1755\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17893\
        );

    \I__1754\ : Span12Mux_h
    port map (
            O => \N__17896\,
            I => \N__17890\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__17893\,
            I => buf_adcdata4_2
        );

    \I__1752\ : Odrv12
    port map (
            O => \N__17890\,
            I => buf_adcdata4_2
        );

    \I__1751\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17881\
        );

    \I__1750\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17878\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__17881\,
            I => \N__17875\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__17878\,
            I => buf_adcdata2_4
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__17875\,
            I => buf_adcdata2_4
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__17870\,
            I => \N__17865\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__17869\,
            I => \N__17862\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__17868\,
            I => \N__17859\
        );

    \I__1743\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17856\
        );

    \I__1742\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17851\
        );

    \I__1741\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17851\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__17856\,
            I => cmd_rdadctmp_13_adj_1063
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__17851\,
            I => cmd_rdadctmp_13_adj_1063
        );

    \I__1738\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17839\
        );

    \I__1737\ : InMux
    port map (
            O => \N__17845\,
            I => \N__17839\
        );

    \I__1736\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17836\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__17839\,
            I => cmd_rdadctmp_14_adj_1062
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__17836\,
            I => cmd_rdadctmp_14_adj_1062
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__17831\,
            I => \N__17826\
        );

    \I__1732\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17823\
        );

    \I__1731\ : InMux
    port map (
            O => \N__17829\,
            I => \N__17818\
        );

    \I__1730\ : InMux
    port map (
            O => \N__17826\,
            I => \N__17818\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__17823\,
            I => cmd_rdadctmp_11_adj_1065
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__17818\,
            I => cmd_rdadctmp_11_adj_1065
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__17813\,
            I => \N__17809\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__17812\,
            I => \N__17805\
        );

    \I__1725\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17800\
        );

    \I__1724\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17800\
        );

    \I__1723\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17797\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__17800\,
            I => cmd_rdadctmp_12_adj_1064
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__17797\,
            I => cmd_rdadctmp_12_adj_1064
        );

    \I__1720\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__17789\,
            I => \N__17785\
        );

    \I__1718\ : InMux
    port map (
            O => \N__17788\,
            I => \N__17782\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__17785\,
            I => \N__17779\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__17782\,
            I => buf_adcdata1_5
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__17779\,
            I => buf_adcdata1_5
        );

    \I__1714\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__17771\,
            I => \N__17767\
        );

    \I__1712\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17764\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__17767\,
            I => \N__17761\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__17764\,
            I => buf_adcdata1_7
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__17761\,
            I => buf_adcdata1_7
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__1707\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17749\
        );

    \I__1706\ : InMux
    port map (
            O => \N__17752\,
            I => \N__17746\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17740\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__17746\,
            I => \N__17740\
        );

    \I__1703\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17737\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__17740\,
            I => \N__17734\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__17737\,
            I => buf_adcdata4_5
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__17734\,
            I => buf_adcdata4_5
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__17729\,
            I => \N__17724\
        );

    \I__1698\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17717\
        );

    \I__1697\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17717\
        );

    \I__1696\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17717\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__17717\,
            I => cmd_rdadctmp_13_adj_1136
        );

    \I__1694\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17711\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__17711\,
            I => \N__17706\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__17710\,
            I => \N__17703\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__17709\,
            I => \N__17700\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__17706\,
            I => \N__17697\
        );

    \I__1689\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17692\
        );

    \I__1688\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17692\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__17697\,
            I => cmd_rdadctmp_14_adj_1135
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__17692\,
            I => cmd_rdadctmp_14_adj_1135
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__1684\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__17681\,
            I => \N__17677\
        );

    \I__1682\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17674\
        );

    \I__1681\ : Span4Mux_h
    port map (
            O => \N__17677\,
            I => \N__17668\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__17674\,
            I => \N__17668\
        );

    \I__1679\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17665\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__17668\,
            I => \N__17662\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__17665\,
            I => buf_adcdata4_6
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__17662\,
            I => buf_adcdata4_6
        );

    \I__1675\ : InMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__17654\,
            I => \N__17650\
        );

    \I__1673\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17647\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__17650\,
            I => \N__17644\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__17647\,
            I => buf_adcdata2_5
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__17644\,
            I => buf_adcdata2_5
        );

    \I__1669\ : InMux
    port map (
            O => \N__17639\,
            I => \N__17635\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \N__17632\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__17635\,
            I => \N__17629\
        );

    \I__1666\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17626\
        );

    \I__1665\ : Span4Mux_h
    port map (
            O => \N__17629\,
            I => \N__17623\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__17626\,
            I => buf_adcdata2_6
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__17623\,
            I => buf_adcdata2_6
        );

    \I__1662\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17614\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__17617\,
            I => \N__17611\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__17614\,
            I => \N__17608\
        );

    \I__1659\ : InMux
    port map (
            O => \N__17611\,
            I => \N__17605\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__17608\,
            I => \N__17602\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__17605\,
            I => buf_adcdata2_7
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__17602\,
            I => buf_adcdata2_7
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__17597\,
            I => \N__17592\
        );

    \I__1654\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17585\
        );

    \I__1653\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17585\
        );

    \I__1652\ : InMux
    port map (
            O => \N__17592\,
            I => \N__17585\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__17585\,
            I => cmd_rdadctmp_15_adj_1061
        );

    \I__1650\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__17579\,
            I => \N__17576\
        );

    \I__1648\ : Span4Mux_v
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__1647\ : Span4Mux_v
    port map (
            O => \N__17573\,
            I => \N__17569\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__17572\,
            I => \N__17566\
        );

    \I__1645\ : Sp12to4
    port map (
            O => \N__17569\,
            I => \N__17563\
        );

    \I__1644\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17560\
        );

    \I__1643\ : Span12Mux_h
    port map (
            O => \N__17563\,
            I => \N__17557\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__17560\,
            I => buf_adcdata2_3
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__17557\,
            I => buf_adcdata2_3
        );

    \I__1640\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__17549\,
            I => n4301
        );

    \I__1638\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__17543\,
            I => \N__17540\
        );

    \I__1636\ : Sp12to4
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__1635\ : Span12Mux_v
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__1634\ : Span12Mux_h
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__1633\ : Odrv12
    port map (
            O => \N__17531\,
            I => buf_data2_0
        );

    \I__1632\ : InMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__17525\,
            I => \N__17522\
        );

    \I__1630\ : Span12Mux_h
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__17519\,
            I => buf_data2_1
        );

    \I__1628\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__1626\ : Span4Mux_v
    port map (
            O => \N__17510\,
            I => \N__17507\
        );

    \I__1625\ : Sp12to4
    port map (
            O => \N__17507\,
            I => \N__17504\
        );

    \I__1624\ : Span12Mux_h
    port map (
            O => \N__17504\,
            I => \N__17501\
        );

    \I__1623\ : Odrv12
    port map (
            O => \N__17501\,
            I => buf_data2_2
        );

    \I__1622\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17495\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__17495\,
            I => n4307
        );

    \I__1620\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17489\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__17489\,
            I => n4306
        );

    \I__1618\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17483\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__17483\,
            I => n4308
        );

    \I__1616\ : InMux
    port map (
            O => \N__17480\,
            I => \N__17477\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__17477\,
            I => buf_data2_6
        );

    \I__1614\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17469\
        );

    \I__1613\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17464\
        );

    \I__1612\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17464\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__17469\,
            I => buf_adcdata4_7
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__17464\,
            I => buf_adcdata4_7
        );

    \I__1609\ : InMux
    port map (
            O => \N__17459\,
            I => \N__17456\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__17456\,
            I => buf_data2_7
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__1606\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__17444\,
            I => buf_data2_4
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__17441\,
            I => \n4304_cascade_\
        );

    \I__1602\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17435\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__17435\,
            I => buf_data2_5
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__17432\,
            I => \n4303_cascade_\
        );

    \I__1599\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17426\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__17426\,
            I => n4302
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__17423\,
            I => \N__17419\
        );

    \I__1596\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17414\
        );

    \I__1595\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17414\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__17414\,
            I => cmd_rdadctmp_5_adj_1071
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__17411\,
            I => \N__17407\
        );

    \I__1592\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17402\
        );

    \I__1591\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17402\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__17402\,
            I => cmd_rdadctmp_3_adj_1073
        );

    \I__1589\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17393\
        );

    \I__1588\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17393\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__17393\,
            I => cmd_rdadctmp_4_adj_1072
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__17390\,
            I => \n14_adj_1035_cascade_\
        );

    \I__1585\ : IoInMux
    port map (
            O => \N__17387\,
            I => \N__17384\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__17384\,
            I => \N__17381\
        );

    \I__1583\ : IoSpan4Mux
    port map (
            O => \N__17381\,
            I => \N__17378\
        );

    \I__1582\ : Span4Mux_s2_h
    port map (
            O => \N__17378\,
            I => \N__17374\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \N__17371\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__17374\,
            I => \N__17368\
        );

    \I__1579\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__17368\,
            I => \M_CS2\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__17365\,
            I => \M_CS2\
        );

    \I__1576\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17356\
        );

    \I__1575\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__17356\,
            I => n15165
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__17353\,
            I => n15165
        );

    \I__1572\ : InMux
    port map (
            O => \N__17348\,
            I => \N__17345\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__17345\,
            I => \N__17342\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__17342\,
            I => \N__17339\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__17339\,
            I => \N__17336\
        );

    \I__1568\ : Span4Mux_h
    port map (
            O => \N__17336\,
            I => \N__17333\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__17333\,
            I => \M_MISO2\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__17330\,
            I => \n8302_cascade_\
        );

    \I__1565\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17323\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__17326\,
            I => \N__17320\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__17323\,
            I => \N__17317\
        );

    \I__1562\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__17317\,
            I => cmd_rdadctmp_2_adj_1074
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__17314\,
            I => cmd_rdadctmp_2_adj_1074
        );

    \I__1559\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17303\
        );

    \I__1558\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17303\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__17303\,
            I => cmd_rdadctmp_0_adj_1076
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__17300\,
            I => \N__17296\
        );

    \I__1555\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17291\
        );

    \I__1554\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17291\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__17291\,
            I => cmd_rdadctmp_1_adj_1075
        );

    \I__1552\ : InMux
    port map (
            O => \N__17288\,
            I => n14029
        );

    \I__1551\ : InMux
    port map (
            O => \N__17285\,
            I => n14030
        );

    \I__1550\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__17279\,
            I => \N__17272\
        );

    \I__1548\ : ClkMux
    port map (
            O => \N__17278\,
            I => \N__17261\
        );

    \I__1547\ : ClkMux
    port map (
            O => \N__17277\,
            I => \N__17261\
        );

    \I__1546\ : ClkMux
    port map (
            O => \N__17276\,
            I => \N__17261\
        );

    \I__1545\ : ClkMux
    port map (
            O => \N__17275\,
            I => \N__17261\
        );

    \I__1544\ : Glb2LocalMux
    port map (
            O => \N__17272\,
            I => \N__17261\
        );

    \I__1543\ : GlobalMux
    port map (
            O => \N__17261\,
            I => \clk_16MHz\
        );

    \I__1542\ : SRMux
    port map (
            O => \N__17258\,
            I => \N__17254\
        );

    \I__1541\ : SRMux
    port map (
            O => \N__17257\,
            I => \N__17251\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__17254\,
            I => \N__17247\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__17251\,
            I => \N__17244\
        );

    \I__1538\ : SRMux
    port map (
            O => \N__17250\,
            I => \N__17241\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__17247\,
            I => \N__17238\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__17244\,
            I => \N__17235\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__17241\,
            I => \N__17232\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__17238\,
            I => n10522
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__17235\,
            I => n10522
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__17232\,
            I => n10522
        );

    \I__1531\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__1529\ : Span4Mux_v
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__17216\,
            I => \N__17212\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__17215\,
            I => \N__17209\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__1525\ : InMux
    port map (
            O => \N__17209\,
            I => \N__17203\
        );

    \I__1524\ : Span12Mux_h
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__17203\,
            I => buf_adcdata2_0
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__17200\,
            I => buf_adcdata2_0
        );

    \I__1521\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17186\
        );

    \I__1520\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17186\
        );

    \I__1519\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17186\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__17186\,
            I => cmd_rdadctmp_8_adj_1068
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__1516\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17174\
        );

    \I__1515\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17174\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__17174\,
            I => cmd_rdadctmp_7_adj_1069
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__17171\,
            I => \N__17168\
        );

    \I__1512\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17161\
        );

    \I__1510\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17158\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__17161\,
            I => cmd_rdadctmp_6_adj_1070
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__17158\,
            I => cmd_rdadctmp_6_adj_1070
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__1506\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17146\
        );

    \I__1505\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17143\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__17146\,
            I => \N__17140\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__17143\,
            I => secclk_cnt_13
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__17140\,
            I => secclk_cnt_13
        );

    \I__1501\ : InMux
    port map (
            O => \N__17135\,
            I => n14021
        );

    \I__1500\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17128\
        );

    \I__1499\ : InMux
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__17128\,
            I => secclk_cnt_14
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__17125\,
            I => secclk_cnt_14
        );

    \I__1496\ : InMux
    port map (
            O => \N__17120\,
            I => n14022
        );

    \I__1495\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17113\
        );

    \I__1494\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17110\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__17113\,
            I => secclk_cnt_15
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__17110\,
            I => secclk_cnt_15
        );

    \I__1491\ : InMux
    port map (
            O => \N__17105\,
            I => n14023
        );

    \I__1490\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17098\
        );

    \I__1489\ : InMux
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__17098\,
            I => \N__17092\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__17095\,
            I => secclk_cnt_16
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__17092\,
            I => secclk_cnt_16
        );

    \I__1485\ : InMux
    port map (
            O => \N__17087\,
            I => \bfn_3_9_0_\
        );

    \I__1484\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17080\
        );

    \I__1483\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__17080\,
            I => secclk_cnt_17
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__17077\,
            I => secclk_cnt_17
        );

    \I__1480\ : InMux
    port map (
            O => \N__17072\,
            I => n14025
        );

    \I__1479\ : InMux
    port map (
            O => \N__17069\,
            I => \N__17065\
        );

    \I__1478\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17062\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__17065\,
            I => secclk_cnt_18
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__17062\,
            I => secclk_cnt_18
        );

    \I__1475\ : InMux
    port map (
            O => \N__17057\,
            I => n14026
        );

    \I__1474\ : InMux
    port map (
            O => \N__17054\,
            I => n14027
        );

    \I__1473\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17047\
        );

    \I__1472\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17044\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__17047\,
            I => secclk_cnt_20
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__17044\,
            I => secclk_cnt_20
        );

    \I__1469\ : InMux
    port map (
            O => \N__17039\,
            I => n14028
        );

    \I__1468\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__1467\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__17032\,
            I => secclk_cnt_4
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__17029\,
            I => secclk_cnt_4
        );

    \I__1464\ : InMux
    port map (
            O => \N__17024\,
            I => n14012
        );

    \I__1463\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17017\
        );

    \I__1462\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17014\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__17017\,
            I => secclk_cnt_5
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__17014\,
            I => secclk_cnt_5
        );

    \I__1459\ : InMux
    port map (
            O => \N__17009\,
            I => n14013
        );

    \I__1458\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17002\
        );

    \I__1457\ : InMux
    port map (
            O => \N__17005\,
            I => \N__16999\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__17002\,
            I => secclk_cnt_6
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__16999\,
            I => secclk_cnt_6
        );

    \I__1454\ : InMux
    port map (
            O => \N__16994\,
            I => n14014
        );

    \I__1453\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16987\
        );

    \I__1452\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16984\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__16987\,
            I => secclk_cnt_7
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__16984\,
            I => secclk_cnt_7
        );

    \I__1449\ : InMux
    port map (
            O => \N__16979\,
            I => n14015
        );

    \I__1448\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16972\
        );

    \I__1447\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16969\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__16972\,
            I => secclk_cnt_8
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__16969\,
            I => secclk_cnt_8
        );

    \I__1444\ : InMux
    port map (
            O => \N__16964\,
            I => \bfn_3_8_0_\
        );

    \I__1443\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16957\
        );

    \I__1442\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16954\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__16957\,
            I => secclk_cnt_9
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__16954\,
            I => secclk_cnt_9
        );

    \I__1439\ : InMux
    port map (
            O => \N__16949\,
            I => n14017
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__16946\,
            I => \N__16942\
        );

    \I__1437\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__1436\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__16939\,
            I => secclk_cnt_10
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__16936\,
            I => secclk_cnt_10
        );

    \I__1433\ : InMux
    port map (
            O => \N__16931\,
            I => n14018
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__16928\,
            I => \N__16924\
        );

    \I__1431\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16921\
        );

    \I__1430\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__16921\,
            I => secclk_cnt_11
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__16918\,
            I => secclk_cnt_11
        );

    \I__1427\ : InMux
    port map (
            O => \N__16913\,
            I => n14019
        );

    \I__1426\ : InMux
    port map (
            O => \N__16910\,
            I => n14020
        );

    \I__1425\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16904\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__16904\,
            I => n28
        );

    \I__1423\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16898\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__16898\,
            I => n26_adj_1180
        );

    \I__1421\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__16892\,
            I => n10
        );

    \I__1419\ : IoInMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__1417\ : Span4Mux_s2_v
    port map (
            O => \N__16883\,
            I => \N__16880\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__16880\,
            I => \N__16877\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__16877\,
            I => \DDS_MCLK1\
        );

    \I__1414\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16870\
        );

    \I__1413\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16867\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__16870\,
            I => secclk_cnt_0
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__16867\,
            I => secclk_cnt_0
        );

    \I__1410\ : InMux
    port map (
            O => \N__16862\,
            I => \bfn_3_7_0_\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__16859\,
            I => \N__16855\
        );

    \I__1408\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16852\
        );

    \I__1407\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__16852\,
            I => secclk_cnt_1
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__16849\,
            I => secclk_cnt_1
        );

    \I__1404\ : InMux
    port map (
            O => \N__16844\,
            I => n14009
        );

    \I__1403\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16837\
        );

    \I__1402\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16834\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__16837\,
            I => secclk_cnt_2
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__16834\,
            I => secclk_cnt_2
        );

    \I__1399\ : InMux
    port map (
            O => \N__16829\,
            I => n14010
        );

    \I__1398\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16822\
        );

    \I__1397\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16819\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__16822\,
            I => secclk_cnt_3
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__16819\,
            I => secclk_cnt_3
        );

    \I__1394\ : InMux
    port map (
            O => \N__16814\,
            I => n14011
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__16811\,
            I => \n25_cascade_\
        );

    \I__1392\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__16805\,
            I => n27_adj_1173
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__16802\,
            I => \n14114_cascade_\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__16799\,
            I => \n10522_cascade_\
        );

    \I__1388\ : IoInMux
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__16793\,
            I => \N__16790\
        );

    \I__1386\ : IoSpan4Mux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__1385\ : Span4Mux_s1_v
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__1384\ : Sp12to4
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__1383\ : Span12Mux_v
    port map (
            O => \N__16781\,
            I => \N__16777\
        );

    \I__1382\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16774\
        );

    \I__1381\ : Odrv12
    port map (
            O => \N__16777\,
            I => \TEST_LED\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__16774\,
            I => \TEST_LED\
        );

    \I__1379\ : IoInMux
    port map (
            O => \N__16769\,
            I => \N__16766\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__1377\ : IoSpan4Mux
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__1376\ : IoSpan4Mux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__16757\,
            I => \ICE_SYSCLK\
        );

    \I__1374\ : IoInMux
    port map (
            O => \N__16754\,
            I => \N__16750\
        );

    \I__1373\ : IoInMux
    port map (
            O => \N__16753\,
            I => \N__16746\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__16750\,
            I => \N__16742\
        );

    \I__1371\ : IoInMux
    port map (
            O => \N__16749\,
            I => \N__16739\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__16746\,
            I => \N__16736\
        );

    \I__1369\ : IoInMux
    port map (
            O => \N__16745\,
            I => \N__16733\
        );

    \I__1368\ : IoSpan4Mux
    port map (
            O => \N__16742\,
            I => \N__16730\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__16739\,
            I => \N__16727\
        );

    \I__1366\ : IoSpan4Mux
    port map (
            O => \N__16736\,
            I => \N__16722\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__16733\,
            I => \N__16722\
        );

    \I__1364\ : Span4Mux_s1_v
    port map (
            O => \N__16730\,
            I => \N__16719\
        );

    \I__1363\ : Span4Mux_s1_v
    port map (
            O => \N__16727\,
            I => \N__16716\
        );

    \I__1362\ : IoSpan4Mux
    port map (
            O => \N__16722\,
            I => \N__16713\
        );

    \I__1361\ : Sp12to4
    port map (
            O => \N__16719\,
            I => \N__16710\
        );

    \I__1360\ : Sp12to4
    port map (
            O => \N__16716\,
            I => \N__16707\
        );

    \I__1359\ : Span4Mux_s2_h
    port map (
            O => \N__16713\,
            I => \N__16704\
        );

    \I__1358\ : Span12Mux_s9_v
    port map (
            O => \N__16710\,
            I => \N__16701\
        );

    \I__1357\ : Span12Mux_h
    port map (
            O => \N__16707\,
            I => \N__16698\
        );

    \I__1356\ : Sp12to4
    port map (
            O => \N__16704\,
            I => \N__16695\
        );

    \I__1355\ : Span12Mux_v
    port map (
            O => \N__16701\,
            I => \N__16692\
        );

    \I__1354\ : Span12Mux_v
    port map (
            O => \N__16698\,
            I => \N__16689\
        );

    \I__1353\ : Span12Mux_v
    port map (
            O => \N__16695\,
            I => \N__16686\
        );

    \I__1352\ : Span12Mux_h
    port map (
            O => \N__16692\,
            I => \N__16683\
        );

    \I__1351\ : Span12Mux_v
    port map (
            O => \N__16689\,
            I => \N__16678\
        );

    \I__1350\ : Span12Mux_h
    port map (
            O => \N__16686\,
            I => \N__16678\
        );

    \I__1349\ : Odrv12
    port map (
            O => \N__16683\,
            I => \M_CLK4\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__16678\,
            I => \M_CLK4\
        );

    \I__1347\ : IoInMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__1345\ : IoSpan4Mux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__1344\ : Sp12to4
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__1343\ : Span12Mux_s3_v
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__1342\ : Span12Mux_h
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__16655\,
            I => \ICE_GPMO_2\
        );

    \INVcomm_spi.bit_cnt_1603__i3C\ : INV
    port map (
            O => \INVcomm_spi.bit_cnt_1603__i3C_net\,
            I => \N__42424\
        );

    \INVdata_count_i0_i8C\ : INV
    port map (
            O => \INVdata_count_i0_i8C_net\,
            I => \N__51309\
        );

    \INVdata_count_i0_i0C\ : INV
    port map (
            O => \INVdata_count_i0_i0C_net\,
            I => \N__51303\
        );

    \INVdata_cntvec_i0_i8C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i8C_net\,
            I => \N__51294\
        );

    \INVdata_cntvec_i0_i0C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i0C_net\,
            I => \N__51283\
        );

    \INVcomm_spi.MISO_48_7334_7335_setC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_7334_7335_setC_net\,
            I => \N__51131\
        );

    \INVcomm_spi.MISO_48_7334_7335_resetC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_7334_7335_resetC_net\,
            I => \N__51116\
        );

    \INVacadc_trig_329C\ : INV
    port map (
            O => \INVacadc_trig_329C_net\,
            I => \N__51281\
        );

    \INVcomm_spi.imiso_83_7340_7341_setC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_7340_7341_setC_net\,
            I => \N__42420\
        );

    \INVcomm_spi.data_valid_85C\ : INV
    port map (
            O => \INVcomm_spi.data_valid_85C_net\,
            I => \N__51123\
        );

    \INVacadc_skipcnt_i0_i9C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i9C_net\,
            I => \N__51268\
        );

    \INVacadc_skipcnt_i0_i1C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i1C_net\,
            I => \N__51252\
        );

    \INVacadc_skipcnt_i0_i0C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i0C_net\,
            I => \N__51236\
        );

    \INVeis_state_i0C\ : INV
    port map (
            O => \INVeis_state_i0C_net\,
            I => \N__51184\
        );

    \INVeis_end_328C\ : INV
    port map (
            O => \INVeis_end_328C_net\,
            I => \N__51166\
        );

    \INVcomm_spi.imiso_83_7340_7341_resetC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_7340_7341_resetC_net\,
            I => \N__42440\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged2WCLKN_net\,
            I => \N__51260\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged3WCLKN_net\,
            I => \N__51288\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged8WCLKN_net\,
            I => \N__51175\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged4WCLKN_net\,
            I => \N__51306\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged9WCLKN_net\,
            I => \N__51210\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged11WCLKN_net\,
            I => \N__51227\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged5WCLKN_net\,
            I => \N__51314\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged0WCLKN_net\,
            I => \N__51135\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged10WCLKN_net\,
            I => \N__51193\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged6WCLKN_net\,
            I => \N__51318\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged1WCLKN_net\,
            I => \N__51157\
        );

    \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN\ : INV
    port map (
            O => \INVraw_buf1_raw_buf4_merged_raw_buf3_merged_raw_buf2_merged7WCLKN_net\,
            I => \N__51320\
        );

    \IN_MUX_bfv_3_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_7_0_\
        );

    \IN_MUX_bfv_3_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n14016,
            carryinitout => \bfn_3_8_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n14024,
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \n13966_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13974,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13958,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n13949,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n14038,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n14047,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_6_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_16_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i11_4_lut_adj_191_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17005\,
            in1 => \N__17131\,
            in2 => \N__16946\,
            in3 => \N__16825\,
            lcout => n27_adj_1173,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17116\,
            in1 => \N__16975\,
            in2 => \N__16859\,
            in3 => \N__17020\,
            lcout => OPEN,
            ltout => \n25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_193_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16907\,
            in1 => \N__16901\,
            in2 => \N__16811\,
            in3 => \N__16808\,
            lcout => OPEN,
            ltout => \n14114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_194_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17050\,
            in1 => \N__16895\,
            in2 => \N__16802\,
            in3 => \N__18518\,
            lcout => n10522,
            ltout => \n10522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SecClk_321_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__16780\,
            in1 => \_gnd_net_\,
            in2 => \N__16799\,
            in3 => \_gnd_net_\,
            lcout => \TEST_LED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17277\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_189_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17068\,
            in1 => \N__16873\,
            in2 => \N__16928\,
            in3 => \N__17035\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_190_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17102\,
            in1 => \N__16990\,
            in2 => \N__17153\,
            in3 => \N__16840\,
            lcout => n26_adj_1180,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16960\,
            in2 => \_gnd_net_\,
            in3 => \N__17083\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_58_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36410\,
            in2 => \_gnd_net_\,
            in3 => \N__35617\,
            lcout => n15165,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_16MHz_I_0_1_lut_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DDS_MCLK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secclk_cnt_1601_1602__i1_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16874\,
            in2 => \_gnd_net_\,
            in3 => \N__16862\,
            lcout => secclk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_3_7_0_\,
            carryout => n14009,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i2_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16858\,
            in2 => \_gnd_net_\,
            in3 => \N__16844\,
            lcout => secclk_cnt_1,
            ltout => OPEN,
            carryin => n14009,
            carryout => n14010,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i3_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16841\,
            in2 => \_gnd_net_\,
            in3 => \N__16829\,
            lcout => secclk_cnt_2,
            ltout => OPEN,
            carryin => n14010,
            carryout => n14011,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i4_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16826\,
            in2 => \_gnd_net_\,
            in3 => \N__16814\,
            lcout => secclk_cnt_3,
            ltout => OPEN,
            carryin => n14011,
            carryout => n14012,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i5_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17036\,
            in2 => \_gnd_net_\,
            in3 => \N__17024\,
            lcout => secclk_cnt_4,
            ltout => OPEN,
            carryin => n14012,
            carryout => n14013,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i6_LC_3_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17021\,
            in2 => \_gnd_net_\,
            in3 => \N__17009\,
            lcout => secclk_cnt_5,
            ltout => OPEN,
            carryin => n14013,
            carryout => n14014,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i7_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17006\,
            in2 => \_gnd_net_\,
            in3 => \N__16994\,
            lcout => secclk_cnt_6,
            ltout => OPEN,
            carryin => n14014,
            carryout => n14015,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i8_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16991\,
            in2 => \_gnd_net_\,
            in3 => \N__16979\,
            lcout => secclk_cnt_7,
            ltout => OPEN,
            carryin => n14015,
            carryout => n14016,
            clk => \N__17275\,
            ce => 'H',
            sr => \N__17257\
        );

    \secclk_cnt_1601_1602__i9_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16976\,
            in2 => \_gnd_net_\,
            in3 => \N__16964\,
            lcout => secclk_cnt_8,
            ltout => OPEN,
            carryin => \bfn_3_8_0_\,
            carryout => n14017,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i10_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16961\,
            in2 => \_gnd_net_\,
            in3 => \N__16949\,
            lcout => secclk_cnt_9,
            ltout => OPEN,
            carryin => n14017,
            carryout => n14018,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i11_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16945\,
            in2 => \_gnd_net_\,
            in3 => \N__16931\,
            lcout => secclk_cnt_10,
            ltout => OPEN,
            carryin => n14018,
            carryout => n14019,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i12_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16927\,
            in2 => \_gnd_net_\,
            in3 => \N__16913\,
            lcout => secclk_cnt_11,
            ltout => OPEN,
            carryin => n14019,
            carryout => n14020,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i13_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18547\,
            in2 => \_gnd_net_\,
            in3 => \N__16910\,
            lcout => secclk_cnt_12,
            ltout => OPEN,
            carryin => n14020,
            carryout => n14021,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i14_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17149\,
            in2 => \_gnd_net_\,
            in3 => \N__17135\,
            lcout => secclk_cnt_13,
            ltout => OPEN,
            carryin => n14021,
            carryout => n14022,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i15_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17132\,
            in2 => \_gnd_net_\,
            in3 => \N__17120\,
            lcout => secclk_cnt_14,
            ltout => OPEN,
            carryin => n14022,
            carryout => n14023,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i16_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17117\,
            in2 => \_gnd_net_\,
            in3 => \N__17105\,
            lcout => secclk_cnt_15,
            ltout => OPEN,
            carryin => n14023,
            carryout => n14024,
            clk => \N__17276\,
            ce => 'H',
            sr => \N__17250\
        );

    \secclk_cnt_1601_1602__i17_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17101\,
            in2 => \_gnd_net_\,
            in3 => \N__17087\,
            lcout => secclk_cnt_16,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => n14025,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \secclk_cnt_1601_1602__i18_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17084\,
            in2 => \_gnd_net_\,
            in3 => \N__17072\,
            lcout => secclk_cnt_17,
            ltout => OPEN,
            carryin => n14025,
            carryout => n14026,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \secclk_cnt_1601_1602__i19_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17069\,
            in2 => \_gnd_net_\,
            in3 => \N__17057\,
            lcout => secclk_cnt_18,
            ltout => OPEN,
            carryin => n14026,
            carryout => n14027,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \secclk_cnt_1601_1602__i20_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18568\,
            in2 => \_gnd_net_\,
            in3 => \N__17054\,
            lcout => secclk_cnt_19,
            ltout => OPEN,
            carryin => n14027,
            carryout => n14028,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \secclk_cnt_1601_1602__i21_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17051\,
            in2 => \_gnd_net_\,
            in3 => \N__17039\,
            lcout => secclk_cnt_20,
            ltout => OPEN,
            carryin => n14028,
            carryout => n14029,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \secclk_cnt_1601_1602__i22_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18583\,
            in2 => \_gnd_net_\,
            in3 => \N__17288\,
            lcout => secclk_cnt_21,
            ltout => OPEN,
            carryin => n14029,
            carryout => n14030,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \secclk_cnt_1601_1602__i23_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18532\,
            in2 => \_gnd_net_\,
            in3 => \N__17285\,
            lcout => secclk_cnt_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__17278\,
            ce => 'H',
            sr => \N__17258\
        );

    \ADC_VAC2.ADC_DATA_i0_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53685\,
            in1 => \N__53436\,
            in2 => \N__17215\,
            in3 => \N__17195\,
            lcout => buf_adcdata2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i9_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46004\,
            in1 => \N__53437\,
            in2 => \N__42931\,
            in3 => \N__17194\,
            lcout => cmd_rdadctmp_9_adj_1067,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i8_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__46003\,
            in1 => \N__17193\,
            in2 => \N__17183\,
            in3 => \N__53438\,
            lcout => cmd_rdadctmp_8_adj_1068,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i7_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__53435\,
            in1 => \N__17179\,
            in2 => \N__17171\,
            in3 => \N__46002\,
            lcout => cmd_rdadctmp_7_adj_1069,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i10_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53434\,
            in1 => \N__42927\,
            in2 => \N__46696\,
            in3 => \N__46001\,
            lcout => cmd_rdadctmp_10_adj_1066,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51275\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_17_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36449\,
            in2 => \_gnd_net_\,
            in3 => \N__35616\,
            lcout => n15150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i6_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__53391\,
            in1 => \N__17164\,
            in2 => \N__46038\,
            in3 => \N__17422\,
            lcout => cmd_rdadctmp_6_adj_1070,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i3_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__17327\,
            in1 => \N__45993\,
            in2 => \N__17411\,
            in3 => \N__53392\,
            lcout => cmd_rdadctmp_3_adj_1073,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i5_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__17399\,
            in1 => \N__45997\,
            in2 => \N__17423\,
            in3 => \N__53393\,
            lcout => cmd_rdadctmp_5_adj_1071,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i4_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__53390\,
            in1 => \N__17410\,
            in2 => \N__46037\,
            in3 => \N__17398\,
            lcout => cmd_rdadctmp_4_adj_1072,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.adc_state_i2_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__36429\,
            in1 => \N__53335\,
            in2 => \_gnd_net_\,
            in3 => \N__35618\,
            lcout => \DTRIG_N_957_adj_1077\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51311\,
            ce => \N__35503\,
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_207_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__36428\,
            in1 => \N__53404\,
            in2 => \N__17377\,
            in3 => \N__35608\,
            lcout => OPEN,
            ltout => \n14_adj_1035_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.CS_37_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__53405\,
            in1 => \N__30185\,
            in2 => \N__17390\,
            in3 => \N__17360\,
            lcout => \M_CS2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i1_3_lut_adj_4_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__30186\,
            in1 => \N__17359\,
            in2 => \_gnd_net_\,
            in3 => \N__53403\,
            lcout => n8302,
            ltout => \n8302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i0_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__53406\,
            in1 => \N__17348\,
            in2 => \N__17330\,
            in3 => \N__17308\,
            lcout => cmd_rdadctmp_0_adj_1076,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i2_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__45949\,
            in1 => \N__17299\,
            in2 => \N__17326\,
            in3 => \N__53408\,
            lcout => cmd_rdadctmp_2_adj_1074,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i1_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53407\,
            in1 => \N__17309\,
            in2 => \N__17300\,
            in3 => \N__45948\,
            lcout => cmd_rdadctmp_1_adj_1075,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i7_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__27527\,
            in1 => \N__18059\,
            in2 => \N__25967\,
            in3 => \N__17473\,
            lcout => buf_adcdata4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1525_i7_4_lut_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__17480\,
            in1 => \N__48060\,
            in2 => \N__17687\,
            in3 => \N__47339\,
            lcout => n4302,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i3_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__20811\,
            in1 => \N__25962\,
            in2 => \N__18233\,
            in3 => \N__27528\,
            lcout => buf_adcdata4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1525_i8_4_lut_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__47338\,
            in1 => \N__17472\,
            in2 => \N__48085\,
            in3 => \N__17459\,
            lcout => n4301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1525_i5_4_lut_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__48072\,
            in1 => \N__18120\,
            in2 => \N__17453\,
            in3 => \N__47322\,
            lcout => OPEN,
            ltout => \n4304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i4_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39903\,
            in2 => \N__17441\,
            in3 => \N__50274\,
            lcout => comm_buf_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51176\,
            ce => \N__18325\,
            sr => \N__18298\
        );

    \mux_1525_i6_4_lut_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010000"
        )
    port map (
            in0 => \N__48073\,
            in1 => \N__17438\,
            in2 => \N__17756\,
            in3 => \N__47323\,
            lcout => OPEN,
            ltout => \n4303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i5_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39797\,
            in2 => \N__17432\,
            in3 => \N__50275\,
            lcout => comm_buf_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51176\,
            ce => \N__18325\,
            sr => \N__18298\
        );

    \comm_buf_5__i6_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40693\,
            in1 => \N__17429\,
            in2 => \_gnd_net_\,
            in3 => \N__50276\,
            lcout => comm_buf_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51176\,
            ce => \N__18325\,
            sr => \N__18298\
        );

    \comm_buf_5__i7_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39338\,
            in1 => \N__17552\,
            in2 => \_gnd_net_\,
            in3 => \N__50277\,
            lcout => comm_buf_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51176\,
            ce => \N__18325\,
            sr => \N__18298\
        );

    \comm_buf_2__i6_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40739\,
            in1 => \N__18089\,
            in2 => \_gnd_net_\,
            in3 => \N__50340\,
            lcout => comm_buf_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51194\,
            ce => \N__18377\,
            sr => \N__18613\
        );

    \comm_buf_2__i7_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18350\,
            in1 => \N__39397\,
            in2 => \_gnd_net_\,
            in3 => \N__50341\,
            lcout => comm_buf_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51194\,
            ce => \N__18377\,
            sr => \N__18613\
        );

    \mux_1525_i1_4_lut_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__17546\,
            in1 => \N__47230\,
            in2 => \N__48086\,
            in3 => \N__18016\,
            lcout => n4308,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1525_i2_4_lut_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__47231\,
            in1 => \N__48067\,
            in2 => \N__17986\,
            in3 => \N__17528\,
            lcout => n4307,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1525_i3_4_lut_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__17516\,
            in1 => \N__17914\,
            in2 => \N__47336\,
            in3 => \N__48068\,
            lcout => n4306,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i1_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44180\,
            in1 => \N__17498\,
            in2 => \_gnd_net_\,
            in3 => \N__50273\,
            lcout => comm_buf_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51211\,
            ce => \N__18329\,
            sr => \N__18299\
        );

    \comm_buf_5__i2_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50270\,
            in1 => \N__40124\,
            in2 => \_gnd_net_\,
            in3 => \N__17492\,
            lcout => comm_buf_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51211\,
            ce => \N__18329\,
            sr => \N__18299\
        );

    \comm_buf_5__i0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17486\,
            in1 => \N__50272\,
            in2 => \_gnd_net_\,
            in3 => \N__39215\,
            lcout => comm_buf_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51211\,
            ce => \N__18329\,
            sr => \N__18299\
        );

    \comm_buf_5__i3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50271\,
            in1 => \N__44921\,
            in2 => \_gnd_net_\,
            in3 => \N__20792\,
            lcout => comm_buf_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51211\,
            ce => \N__18329\,
            sr => \N__18299\
        );

    \ADC_VAC2.ADC_DATA_i5_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53702\,
            in1 => \N__17653\,
            in2 => \N__17870\,
            in3 => \N__53518\,
            lcout => buf_adcdata2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i6_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53515\,
            in1 => \N__53704\,
            in2 => \N__17638\,
            in3 => \N__17846\,
            lcout => buf_adcdata2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i7_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53703\,
            in1 => \N__53517\,
            in2 => \N__17617\,
            in3 => \N__17596\,
            lcout => buf_adcdata2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i15_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53516\,
            in1 => \N__17845\,
            in2 => \N__17597\,
            in3 => \N__46079\,
            lcout => cmd_rdadctmp_15_adj_1061,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i16_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46080\,
            in1 => \N__17595\,
            in2 => \N__20445\,
            in3 => \N__53519\,
            lcout => cmd_rdadctmp_16_adj_1060,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i3_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53695\,
            in1 => \N__53523\,
            in2 => \N__17572\,
            in3 => \N__17829\,
            lcout => buf_adcdata2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i11_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53520\,
            in1 => \N__46695\,
            in2 => \N__17831\,
            in3 => \N__46076\,
            lcout => cmd_rdadctmp_11_adj_1065,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i15_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__17714\,
            in1 => \N__27415\,
            in2 => \N__18054\,
            in3 => \N__26846\,
            lcout => cmd_rdadctmp_15_adj_1134,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i13_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53521\,
            in1 => \N__17808\,
            in2 => \N__17868\,
            in3 => \N__46077\,
            lcout => cmd_rdadctmp_13_adj_1063,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i4_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53696\,
            in1 => \N__17884\,
            in2 => \N__17813\,
            in3 => \N__53524\,
            lcout => buf_adcdata2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i14_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__53522\,
            in1 => \N__17844\,
            in2 => \N__17869\,
            in3 => \N__46078\,
            lcout => cmd_rdadctmp_14_adj_1062,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51244\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i12_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__17830\,
            in1 => \N__46058\,
            in2 => \N__17812\,
            in3 => \N__53356\,
            lcout => cmd_rdadctmp_12_adj_1064,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i5_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53049\,
            in1 => \N__17788\,
            in2 => \N__19595\,
            in3 => \N__52845\,
            lcout => buf_adcdata1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i7_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53051\,
            in1 => \N__17770\,
            in2 => \N__19793\,
            in3 => \N__52847\,
            lcout => buf_adcdata1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i5_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25940\,
            in1 => \N__17745\,
            in2 => \N__27515\,
            in3 => \N__17728\,
            lcout => buf_adcdata4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i13_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__27482\,
            in1 => \N__18151\,
            in2 => \N__17729\,
            in3 => \N__26839\,
            lcout => cmd_rdadctmp_13_adj_1136,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i14_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__26838\,
            in1 => \N__17727\,
            in2 => \N__17709\,
            in3 => \N__27485\,
            lcout => cmd_rdadctmp_14_adj_1135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i6_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25941\,
            in1 => \N__17673\,
            in2 => \N__17710\,
            in3 => \N__27484\,
            lcout => buf_adcdata4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i16_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__27483\,
            in1 => \N__18055\,
            in2 => \N__19441\,
            in3 => \N__26840\,
            lcout => cmd_rdadctmp_16_adj_1133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51276\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25937\,
            in1 => \N__18015\,
            in2 => \N__18275\,
            in3 => \N__27451\,
            lcout => buf_adcdata4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i1_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27447\,
            in1 => \N__25938\,
            in2 => \N__17954\,
            in3 => \N__17976\,
            lcout => buf_adcdata4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i9_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26843\,
            in1 => \N__17946\,
            in2 => \N__18274\,
            in3 => \N__27453\,
            lcout => cmd_rdadctmp_9_adj_1140,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i10_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__27449\,
            in1 => \N__17931\,
            in2 => \N__17953\,
            in3 => \N__26844\,
            lcout => cmd_rdadctmp_10_adj_1139,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i11_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26841\,
            in1 => \N__18219\,
            in2 => \N__17936\,
            in3 => \N__27452\,
            lcout => cmd_rdadctmp_11_adj_1138,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i2_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27448\,
            in1 => \N__25939\,
            in2 => \N__17910\,
            in3 => \N__17935\,
            lcout => buf_adcdata4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i5_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__26842\,
            in1 => \N__27450\,
            in2 => \N__18203\,
            in3 => \N__18253\,
            lcout => cmd_rdadctmp_5_adj_1144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i7_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__26834\,
            in1 => \N__18242\,
            in2 => \N__27514\,
            in3 => \N__18283\,
            lcout => cmd_rdadctmp_7_adj_1142,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i8_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__18267\,
            in1 => \N__27472\,
            in2 => \N__18287\,
            in3 => \N__26837\,
            lcout => cmd_rdadctmp_8_adj_1141,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i6_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26833\,
            in1 => \N__18241\,
            in2 => \N__27513\,
            in3 => \N__18254\,
            lcout => cmd_rdadctmp_6_adj_1143,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i12_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__18220\,
            in1 => \N__27470\,
            in2 => \N__18150\,
            in3 => \N__26835\,
            lcout => cmd_rdadctmp_12_adj_1137,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i4_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__26832\,
            in1 => \N__18187\,
            in2 => \N__27512\,
            in3 => \N__18202\,
            lcout => cmd_rdadctmp_4_adj_1145,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i3_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__18175\,
            in1 => \N__27471\,
            in2 => \N__18188\,
            in3 => \N__26836\,
            lcout => cmd_rdadctmp_3_adj_1146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19847\,
            in1 => \N__27459\,
            in2 => \N__18176\,
            in3 => \N__26845\,
            lcout => cmd_rdadctmp_2_adj_1147,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i4_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25966\,
            in1 => \N__18121\,
            in2 => \N__18161\,
            in3 => \N__27526\,
            lcout => buf_adcdata4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1481_i7_4_lut_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__47324\,
            in1 => \N__18101\,
            in2 => \N__19528\,
            in3 => \N__48087\,
            lcout => n4146,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1481_i1_4_lut_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__18077\,
            in1 => \N__47326\,
            in2 => \N__48092\,
            in3 => \N__43814\,
            lcout => n4152,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1481_i8_4_lut_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__18359\,
            in1 => \N__48091\,
            in2 => \N__18715\,
            in3 => \N__47325\,
            lcout => n4145,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50268\,
            in1 => \N__44155\,
            in2 => \_gnd_net_\,
            in3 => \N__27545\,
            lcout => comm_buf_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51148\,
            ce => \N__18375\,
            sr => \N__18614\
        );

    \comm_buf_2__i0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50269\,
            in1 => \N__18341\,
            in2 => \_gnd_net_\,
            in3 => \N__39214\,
            lcout => comm_buf_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51148\,
            ce => \N__18375\,
            sr => \N__18614\
        );

    \i1_2_lut_adj_270_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__49536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52310\,
            lcout => n15221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_3_lut_3_lut_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__52309\,
            in1 => \N__50267\,
            in2 => \_gnd_net_\,
            in3 => \N__49535\,
            lcout => n15131,
            ltout => \n15131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_195_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__25558\,
            in1 => \N__50604\,
            in2 => \N__18335\,
            in3 => \N__27809\,
            lcout => n8738,
            ltout => \n8738_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7484_2_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__52312\,
            in1 => \_gnd_net_\,
            in2 => \N__18332\,
            in3 => \_gnd_net_\,
            lcout => n10590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_233_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__42839\,
            in1 => \N__50605\,
            in2 => \N__25572\,
            in3 => \N__27734\,
            lcout => n8847,
            ltout => \n8847_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7505_2_lut_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__52313\,
            in1 => \_gnd_net_\,
            in2 => \N__18302\,
            in3 => \_gnd_net_\,
            lcout => n10611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_201_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__42838\,
            in1 => \N__50603\,
            in2 => \N__25571\,
            in3 => \N__27827\,
            lcout => n8787,
            ltout => \n8787_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7491_2_lut_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__52311\,
            in1 => \_gnd_net_\,
            in2 => \N__18428\,
            in3 => \_gnd_net_\,
            lcout => n10599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1481_i3_4_lut_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__18425\,
            in1 => \N__48069\,
            in2 => \N__18475\,
            in3 => \N__47319\,
            lcout => OPEN,
            ltout => \n4150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i2_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40122\,
            in1 => \_gnd_net_\,
            in2 => \N__18407\,
            in3 => \N__50088\,
            lcout => comm_buf_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51178\,
            ce => \N__18376\,
            sr => \N__18612\
        );

    \comm_buf_2__i3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44907\,
            in1 => \N__32582\,
            in2 => \_gnd_net_\,
            in3 => \N__50089\,
            lcout => comm_buf_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51178\,
            ce => \N__18376\,
            sr => \N__18612\
        );

    \mux_1481_i5_4_lut_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__18404\,
            in1 => \N__48070\,
            in2 => \N__18764\,
            in3 => \N__47320\,
            lcout => OPEN,
            ltout => \n4148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i4_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39947\,
            in1 => \_gnd_net_\,
            in2 => \N__18395\,
            in3 => \N__50090\,
            lcout => comm_buf_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51178\,
            ce => \N__18376\,
            sr => \N__18612\
        );

    \mux_1481_i6_4_lut_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__18392\,
            in1 => \N__48071\,
            in2 => \N__19565\,
            in3 => \N__47321\,
            lcout => OPEN,
            ltout => \n4147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i5_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39809\,
            in2 => \N__18380\,
            in3 => \N__50091\,
            lcout => comm_buf_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51178\,
            ce => \N__18376\,
            sr => \N__18612\
        );

    \i6_4_lut_adj_192_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18584\,
            in1 => \N__18569\,
            in2 => \N__18554\,
            in3 => \N__18533\,
            lcout => n14_adj_1163,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i0_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24305\,
            in1 => \N__50278\,
            in2 => \_gnd_net_\,
            in3 => \N__39213\,
            lcout => comm_buf_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51196\,
            ce => \N__25450\,
            sr => \N__20088\
        );

    \comm_buf_4__i1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44179\,
            in1 => \N__42632\,
            in2 => \_gnd_net_\,
            in3 => \N__50279\,
            lcout => comm_buf_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51196\,
            ce => \N__25450\,
            sr => \N__20088\
        );

    \mux_1457_i3_4_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__18506\,
            in1 => \N__48037\,
            in2 => \N__19709\,
            in3 => \N__47290\,
            lcout => OPEN,
            ltout => \n4062_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i2_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40123\,
            in2 => \N__18485\,
            in3 => \N__50280\,
            lcout => comm_buf_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51196\,
            ce => \N__25450\,
            sr => \N__20088\
        );

    \comm_buf_4__i3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44908\,
            in1 => \N__26516\,
            in2 => \_gnd_net_\,
            in3 => \N__50281\,
            lcout => comm_buf_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51213\,
            ce => \N__25457\,
            sr => \N__20102\
        );

    \ADC_VAC3.ADC_DATA_i2_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49190\,
            in1 => \N__44356\,
            in2 => \N__19472\,
            in3 => \N__18459\,
            lcout => buf_adcdata3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i11_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__49193\,
            in1 => \N__18438\,
            in2 => \N__19471\,
            in3 => \N__48840\,
            lcout => cmd_rdadctmp_11_adj_1101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i12_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__48839\,
            in1 => \N__18648\,
            in2 => \N__18443\,
            in3 => \N__49194\,
            lcout => cmd_rdadctmp_12_adj_1100,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i3_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__49191\,
            in1 => \N__44357\,
            in2 => \N__32619\,
            in3 => \N__18442\,
            lcout => buf_adcdata3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i3_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__52848\,
            in1 => \N__53015\,
            in2 => \N__20525\,
            in3 => \N__18778\,
            lcout => buf_adcdata1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i4_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49192\,
            in1 => \N__44358\,
            in2 => \N__18655\,
            in3 => \N__18753\,
            lcout => buf_adcdata3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51230\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i1_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52851\,
            in1 => \N__18665\,
            in2 => \N__18733\,
            in3 => \N__26115\,
            lcout => cmd_rdadctmp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i2_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52852\,
            in1 => \N__18856\,
            in2 => \N__18734\,
            in3 => \N__26116\,
            lcout => cmd_rdadctmp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i7_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__44355\,
            in1 => \N__18708\,
            in2 => \N__21680\,
            in3 => \N__49201\,
            lcout => buf_adcdata3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i0_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52849\,
            in1 => \N__18664\,
            in2 => \N__18686\,
            in3 => \N__26113\,
            lcout => cmd_rdadctmp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i13_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__18656\,
            in1 => \N__49200\,
            in2 => \N__20322\,
            in3 => \N__48814\,
            lcout => cmd_rdadctmp_13_adj_1099,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i13_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52850\,
            in1 => \N__19488\,
            in2 => \N__19590\,
            in3 => \N__26114\,
            lcout => cmd_rdadctmp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i4_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53050\,
            in1 => \N__18628\,
            in2 => \N__19493\,
            in3 => \N__52853\,
            lcout => buf_adcdata1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51246\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.CS_37_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__18929\,
            in1 => \N__18896\,
            in2 => \N__19648\,
            in3 => \N__52674\,
            lcout => \M_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i24_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52670\,
            in1 => \N__22715\,
            in2 => \N__48252\,
            in3 => \N__26069\,
            lcout => cmd_rdadctmp_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i8_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__26075\,
            in1 => \N__52677\,
            in2 => \N__22477\,
            in3 => \N__18845\,
            lcout => cmd_rdadctmp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52671\,
            in1 => \N__18857\,
            in2 => \N__18811\,
            in3 => \N__26070\,
            lcout => cmd_rdadctmp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i7_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26074\,
            in1 => \N__18844\,
            in2 => \N__18836\,
            in3 => \N__52676\,
            lcout => cmd_rdadctmp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i6_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52673\,
            in1 => \N__18832\,
            in2 => \N__18824\,
            in3 => \N__26073\,
            lcout => cmd_rdadctmp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i5_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26072\,
            in1 => \N__18820\,
            in2 => \N__18797\,
            in3 => \N__52675\,
            lcout => cmd_rdadctmp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i4_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52672\,
            in1 => \N__18793\,
            in2 => \N__18812\,
            in3 => \N__26071\,
            lcout => cmd_rdadctmp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.adc_state_i2_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__52605\,
            in1 => \N__20627\,
            in2 => \_gnd_net_\,
            in3 => \N__20569\,
            lcout => \DTRIG_N_957\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51277\,
            ce => \N__19604\,
            sr => \_gnd_net_\
        );

    \ADC_VAC1.adc_state_i1_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__20568\,
            in1 => \_gnd_net_\,
            in2 => \N__20643\,
            in3 => \N__52606\,
            lcout => adc_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51277\,
            ce => \N__19604\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_224_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20623\,
            in2 => \_gnd_net_\,
            in3 => \N__20566\,
            lcout => n15168,
            ltout => \n15168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i1_3_lut_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__19640\,
            in1 => \_gnd_net_\,
            in2 => \N__18923\,
            in3 => \N__52603\,
            lcout => n8272,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_222_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110010"
        )
    port map (
            in0 => \N__20567\,
            in1 => \N__18907\,
            in2 => \N__20642\,
            in3 => \N__52604\,
            lcout => n14_adj_1039,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_298_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20622\,
            in2 => \_gnd_net_\,
            in3 => \N__20565\,
            lcout => n15153,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.SCLK_35_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011100010"
        )
    port map (
            in0 => \N__20638\,
            in1 => \N__52678\,
            in2 => \N__18880\,
            in3 => \N__20576\,
            lcout => \M_SCLK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51290\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i1_4_lut_adj_6_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000010"
        )
    port map (
            in0 => \N__20574\,
            in1 => \N__52616\,
            in2 => \N__19647\,
            in3 => \N__20636\,
            lcout => \ADC_VAC1.n9312\,
            ltout => \ADC_VAC1.n9312_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i7561_2_lut_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__20637\,
            in1 => \_gnd_net_\,
            in2 => \N__18863\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC1.n10667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i12131_4_lut_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18976\,
            in1 => \N__18991\,
            in2 => \N__19025\,
            in3 => \N__19006\,
            lcout => OPEN,
            ltout => \ADC_VAC1.n15338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i12151_4_lut_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18943\,
            in1 => \N__19039\,
            in2 => \N__18860\,
            in3 => \N__19141\,
            lcout => OPEN,
            ltout => \ADC_VAC1.n15360_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i12914_4_lut_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20575\,
            in1 => \N__18962\,
            in2 => \N__19043\,
            in3 => \N__52617\,
            lcout => \ADC_VAC1.n15553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.bit_cnt_i0_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19040\,
            in2 => \_gnd_net_\,
            in3 => \N__19028\,
            lcout => \ADC_VAC1.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_6_16_0_\,
            carryout => \ADC_VAC1.n13981\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i1_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19024\,
            in2 => \_gnd_net_\,
            in3 => \N__19010\,
            lcout => \ADC_VAC1.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC1.n13981\,
            carryout => \ADC_VAC1.n13982\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i2_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19007\,
            in2 => \_gnd_net_\,
            in3 => \N__18995\,
            lcout => \ADC_VAC1.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC1.n13982\,
            carryout => \ADC_VAC1.n13983\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i3_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18992\,
            in2 => \_gnd_net_\,
            in3 => \N__18980\,
            lcout => \ADC_VAC1.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC1.n13983\,
            carryout => \ADC_VAC1.n13984\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i4_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18977\,
            in2 => \_gnd_net_\,
            in3 => \N__18965\,
            lcout => \ADC_VAC1.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC1.n13984\,
            carryout => \ADC_VAC1.n13985\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i5_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18961\,
            in2 => \_gnd_net_\,
            in3 => \N__18947\,
            lcout => \ADC_VAC1.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC1.n13985\,
            carryout => \ADC_VAC1.n13986\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i6_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18944\,
            in2 => \_gnd_net_\,
            in3 => \N__18932\,
            lcout => \ADC_VAC1.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC1.n13986\,
            carryout => \ADC_VAC1.n13987\,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \ADC_VAC1.bit_cnt_i7_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19142\,
            in2 => \_gnd_net_\,
            in3 => \N__19145\,
            lcout => \ADC_VAC1.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51300\,
            ce => \N__19130\,
            sr => \N__19121\
        );

    \comm_index_0__bdd_4_lut_13254_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__38848\,
            in1 => \N__23537\,
            in2 => \N__22205\,
            in3 => \N__33206\,
            lcout => OPEN,
            ltout => \n16470_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16470_bdd_4_lut_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33207\,
            in1 => \N__20147\,
            in2 => \N__19115\,
            in3 => \N__19112\,
            lcout => n16473,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13205_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__38849\,
            in1 => \N__19100\,
            in2 => \N__19052\,
            in3 => \N__33208\,
            lcout => OPEN,
            ltout => \n16416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16416_bdd_4_lut_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__37878\,
            in1 => \N__33205\,
            in2 => \N__19088\,
            in3 => \N__33785\,
            lcout => OPEN,
            ltout => \n16419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i981538_i1_3_lut_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19085\,
            in2 => \N__19079\,
            in3 => \N__33535\,
            lcout => OPEN,
            ltout => \n7_adj_1238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i5_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33536\,
            in1 => \N__20936\,
            in2 => \N__19076\,
            in3 => \N__33352\,
            lcout => comm_tx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51126\,
            ce => \N__43110\,
            sr => \N__22393\
        );

    \mux_1469_i6_4_lut_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__19073\,
            in1 => \N__48013\,
            in2 => \N__23177\,
            in3 => \N__47335\,
            lcout => OPEN,
            ltout => \n4103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i5_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39796\,
            in1 => \_gnd_net_\,
            in2 => \N__19055\,
            in3 => \N__50112\,
            lcout => comm_buf_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51138\,
            ce => \N__19202\,
            sr => \N__19178\
        );

    \comm_buf_3__i6_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40692\,
            in1 => \N__29045\,
            in2 => \_gnd_net_\,
            in3 => \N__50113\,
            lcout => comm_buf_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51138\,
            ce => \N__19202\,
            sr => \N__19178\
        );

    \comm_buf_3__i7_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39360\,
            in1 => \N__45836\,
            in2 => \_gnd_net_\,
            in3 => \N__50114\,
            lcout => comm_buf_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51138\,
            ce => \N__19202\,
            sr => \N__19178\
        );

    \comm_buf_3__i0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__46718\,
            in1 => \N__50337\,
            in2 => \_gnd_net_\,
            in3 => \N__39209\,
            lcout => comm_buf_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51149\,
            ce => \N__19201\,
            sr => \N__19174\
        );

    \mux_1469_i2_4_lut_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__19247\,
            in1 => \N__48006\,
            in2 => \N__25799\,
            in3 => \N__47088\,
            lcout => OPEN,
            ltout => \n4107_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i1_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__44171\,
            in1 => \_gnd_net_\,
            in2 => \N__19226\,
            in3 => \N__50338\,
            lcout => comm_buf_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51149\,
            ce => \N__19201\,
            sr => \N__19174\
        );

    \mux_1469_i3_4_lut_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__19223\,
            in1 => \N__48005\,
            in2 => \N__19285\,
            in3 => \N__47087\,
            lcout => \comm_buf_3_7_N_501_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39939\,
            in1 => \N__21554\,
            in2 => \_gnd_net_\,
            in3 => \N__50339\,
            lcout => comm_buf_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51149\,
            ce => \N__19201\,
            sr => \N__19174\
        );

    \i12238_3_lut_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22121\,
            in1 => \N__38840\,
            in2 => \_gnd_net_\,
            in3 => \N__23453\,
            lcout => n15448,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12178_3_lut_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__38842\,
            in1 => \_gnd_net_\,
            in2 => \N__19154\,
            in3 => \N__21125\,
            lcout => OPEN,
            ltout => \n15388_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16386_bdd_4_lut_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100110101000"
        )
    port map (
            in0 => \N__19301\,
            in1 => \N__33522\,
            in2 => \N__19331\,
            in3 => \N__29117\,
            lcout => OPEN,
            ltout => \n16389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i2_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33523\,
            in1 => \N__21029\,
            in2 => \N__19328\,
            in3 => \N__33347\,
            lcout => comm_tx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51161\,
            ce => \N__43127\,
            sr => \N__22348\
        );

    \i12237_3_lut_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19325\,
            in1 => \N__38841\,
            in2 => \_gnd_net_\,
            in3 => \N__19319\,
            lcout => OPEN,
            ltout => \n15447_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_13182_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__33521\,
            in1 => \N__19310\,
            in2 => \N__19304\,
            in3 => \N__33212\,
            lcout => n16386,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7554_3_lut_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__43078\,
            in1 => \N__52444\,
            in2 => \_gnd_net_\,
            in3 => \N__39263\,
            lcout => n10660,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i18_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25945\,
            in1 => \N__19278\,
            in2 => \N__25751\,
            in3 => \N__27511\,
            lcout => buf_adcdata4_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7498_2_lut_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52445\,
            in2 => \_gnd_net_\,
            in3 => \N__25448\,
            lcout => n10604,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9698_2_lut_3_lut_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__33971\,
            in1 => \N__50110\,
            in2 => \_gnd_net_\,
            in3 => \N__49537\,
            lcout => n14_adj_1169,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i1_3_lut_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33871\,
            in1 => \N__24512\,
            in2 => \_gnd_net_\,
            in3 => \N__48014\,
            lcout => n4209,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12187_3_lut_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21116\,
            in1 => \N__19259\,
            in2 => \_gnd_net_\,
            in3 => \N__38845\,
            lcout => n15397,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12213_3_lut_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__38843\,
            in1 => \N__19409\,
            in2 => \_gnd_net_\,
            in3 => \N__19403\,
            lcout => n15423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13230_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23672\,
            in1 => \N__33209\,
            in2 => \N__22025\,
            in3 => \N__38844\,
            lcout => OPEN,
            ltout => \n16440_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16440_bdd_4_lut_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33210\,
            in1 => \N__23288\,
            in2 => \N__19391\,
            in3 => \N__21092\,
            lcout => n16443,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_13225_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__33532\,
            in1 => \N__33211\,
            in2 => \N__19388\,
            in3 => \N__20981\,
            lcout => OPEN,
            ltout => \n16392_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16392_bdd_4_lut_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__31109\,
            in1 => \N__19379\,
            in2 => \N__19373\,
            in3 => \N__33533\,
            lcout => OPEN,
            ltout => \n16395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i3_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33534\,
            in1 => \N__19370\,
            in2 => \N__19364\,
            in3 => \N__33348\,
            lcout => comm_tx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51197\,
            ce => \N__43126\,
            sr => \N__22370\
        );

    \ADC_VAC2.cmd_rdadctmp_i31_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53354\,
            in1 => \N__48212\,
            in2 => \N__48139\,
            in3 => \N__46081\,
            lcout => cmd_rdadctmp_31_adj_1045,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.SCLK_35_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011100010"
        )
    port map (
            in0 => \N__36466\,
            in1 => \N__53355\,
            in2 => \N__19348\,
            in3 => \N__35609\,
            lcout => \M_SCLK2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i8_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__49195\,
            in1 => \N__43827\,
            in2 => \N__23999\,
            in3 => \N__48815\,
            lcout => cmd_rdadctmp_8_adj_1104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i1_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__44354\,
            in1 => \N__27571\,
            in2 => \N__20396\,
            in3 => \N__49196\,
            lcout => buf_adcdata3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51214\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i5_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__44352\,
            in1 => \N__19551\,
            in2 => \N__20326\,
            in3 => \N__49199\,
            lcout => buf_adcdata3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i6_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49197\,
            in1 => \N__44353\,
            in2 => \N__20297\,
            in3 => \N__19515\,
            lcout => buf_adcdata3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i12_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20514\,
            in1 => \N__52836\,
            in2 => \N__19492\,
            in3 => \N__26126\,
            lcout => cmd_rdadctmp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i10_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__49198\,
            in1 => \N__20392\,
            in2 => \N__19470\,
            in3 => \N__48763\,
            lcout => cmd_rdadctmp_10_adj_1102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i8_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27372\,
            in1 => \N__25926\,
            in2 => \N__24336\,
            in3 => \N__19448\,
            lcout => buf_adcdata4_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i9_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__25925\,
            in1 => \N__27376\,
            in2 => \N__42652\,
            in3 => \N__19423\,
            lcout => buf_adcdata4_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i17_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__27373\,
            in1 => \N__19447\,
            in2 => \N__19424\,
            in3 => \N__26855\,
            lcout => cmd_rdadctmp_17_adj_1132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i18_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__26854\,
            in1 => \N__19422\,
            in2 => \N__19726\,
            in3 => \N__27378\,
            lcout => cmd_rdadctmp_18_adj_1131,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i19_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__27374\,
            in1 => \N__19722\,
            in2 => \N__22500\,
            in3 => \N__26856\,
            lcout => cmd_rdadctmp_19_adj_1130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i10_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25924\,
            in1 => \N__19695\,
            in2 => \N__19727\,
            in3 => \N__27377\,
            lcout => buf_adcdata4_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i20_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__27375\,
            in1 => \N__22656\,
            in2 => \N__22501\,
            in3 => \N__26857\,
            lcout => cmd_rdadctmp_20_adj_1129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51247\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i1_4_lut_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__20632\,
            in1 => \N__52619\,
            in2 => \N__19658\,
            in3 => \N__30658\,
            lcout => OPEN,
            ltout => \ADC_VAC1.n15263_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i1_2_lut_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__20573\,
            in1 => \_gnd_net_\,
            in2 => \N__19673\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC1.n15264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.adc_state_i0_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__20580\,
            in1 => \N__52620\,
            in2 => \N__20644\,
            in3 => \N__19670\,
            lcout => adc_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51264\,
            ce => \N__19664\,
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i30_4_lut_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110000001"
        )
    port map (
            in0 => \N__30659\,
            in1 => \N__20631\,
            in2 => \N__20581\,
            in3 => \N__19657\,
            lcout => OPEN,
            ltout => \ADC_VAC1.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.i13056_2_lut_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19607\,
            in3 => \N__52618\,
            lcout => \ADC_VAC1.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i15_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26089\,
            in1 => \N__19782\,
            in2 => \N__52778\,
            in3 => \N__21723\,
            lcout => cmd_rdadctmp_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i14_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19591\,
            in1 => \N__52679\,
            in2 => \N__21727\,
            in3 => \N__26088\,
            lcout => cmd_rdadctmp_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i1_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19805\,
            in1 => \N__27460\,
            in2 => \N__19846\,
            in3 => \N__26858\,
            lcout => cmd_rdadctmp_1_adj_1148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i0_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19804\,
            in1 => \N__27468\,
            in2 => \N__19829\,
            in3 => \N__26797\,
            lcout => cmd_rdadctmp_0_adj_1149,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i16_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__19783\,
            in1 => \N__26127\,
            in2 => \N__32166\,
            in3 => \N__52774\,
            lcout => cmd_rdadctmp_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51291\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i17_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__20458\,
            in1 => \N__46062\,
            in2 => \N__46227\,
            in3 => \N__53402\,
            lcout => cmd_rdadctmp_17_adj_1059,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ICE_GPMO_0_I_0_1_lut_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32771\,
            lcout => \M_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_7348_7349_reset_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20924\,
            in1 => \N__20912\,
            in2 => \_gnd_net_\,
            in3 => \N__21617\,
            lcout => \comm_spi.n10460\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42466\,
            ce => 'H',
            sr => \N__20885\
        );

    \comm_tx_buf_i0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__20837\,
            in1 => \N__33520\,
            in2 => \N__20990\,
            in3 => \N__33353\,
            lcout => comm_tx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51119\,
            ce => \N__43134\,
            sr => \N__22394\
        );

    \i12201_3_lut_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25043\,
            in1 => \N__23615\,
            in2 => \_gnd_net_\,
            in3 => \N__38846\,
            lcout => n15411,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12181_3_lut_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19748\,
            in1 => \N__19739\,
            in2 => \_gnd_net_\,
            in3 => \N__38847\,
            lcout => n15391,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16410_bdd_4_lut_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__33106\,
            in1 => \N__33970\,
            in2 => \N__41897\,
            in3 => \N__19886\,
            lcout => OPEN,
            ltout => \n16413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10400_3_lut_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19880\,
            in2 => \N__19931\,
            in3 => \N__33349\,
            lcout => n13493,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__38810\,
            in1 => \N__22229\,
            in2 => \N__33168\,
            in3 => \N__23567\,
            lcout => OPEN,
            ltout => \n16518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16518_bdd_4_lut_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__19928\,
            in1 => \N__33110\,
            in2 => \N__19919\,
            in3 => \N__20135\,
            lcout => OPEN,
            ltout => \n16521_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i6_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__33350\,
            in1 => \N__19916\,
            in2 => \N__19910\,
            in3 => \N__33531\,
            lcout => comm_tx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51127\,
            ce => \N__43122\,
            sr => \N__22383\
        );

    \comm_index_0__bdd_4_lut_13200_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__19907\,
            in1 => \N__33104\,
            in2 => \N__19895\,
            in3 => \N__38809\,
            lcout => n16410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16488_bdd_4_lut_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__33105\,
            in1 => \N__23369\,
            in2 => \N__24794\,
            in3 => \N__25127\,
            lcout => n16491,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13195_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__19874\,
            in1 => \N__33182\,
            in2 => \N__19862\,
            in3 => \N__38839\,
            lcout => OPEN,
            ltout => \n16404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16404_bdd_4_lut_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33183\,
            in1 => \N__34560\,
            in2 => \N__19850\,
            in3 => \N__41105\,
            lcout => OPEN,
            ltout => \n16407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i979126_i1_3_lut_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19976\,
            in2 => \N__20006\,
            in3 => \N__33524\,
            lcout => n7_adj_1240,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16512_bdd_4_lut_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__33181\,
            in1 => \N__20003\,
            in2 => \N__19991\,
            in3 => \N__19970\,
            lcout => n16515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13284_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23774\,
            in1 => \N__33180\,
            in2 => \N__22091\,
            in3 => \N__38838\,
            lcout => n16512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16422_bdd_4_lut_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__33184\,
            in1 => \N__23645\,
            in2 => \N__24707\,
            in3 => \N__24980\,
            lcout => OPEN,
            ltout => \n16425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__33351\,
            in1 => \N__19964\,
            in2 => \N__19958\,
            in3 => \N__33525\,
            lcout => comm_tx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51139\,
            ce => \N__43138\,
            sr => \N__22392\
        );

    \comm_spi.data_tx_i7_7337_7338_set_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27668\,
            in1 => \N__27794\,
            in2 => \_gnd_net_\,
            in3 => \N__28994\,
            lcout => \comm_spi.n10448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42467\,
            ce => 'H',
            sr => \N__30779\
        );

    \i1_2_lut_adj_60_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36587\,
            in2 => \_gnd_net_\,
            in3 => \N__33566\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1457_i5_4_lut_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__19955\,
            in1 => \N__48035\,
            in2 => \N__20491\,
            in3 => \N__47291\,
            lcout => OPEN,
            ltout => \n4060_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i4_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39932\,
            in1 => \_gnd_net_\,
            in2 => \N__19934\,
            in3 => \N__50325\,
            lcout => comm_buf_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51162\,
            ce => \N__25449\,
            sr => \N__20095\
        );

    \comm_buf_4__i5_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39798\,
            in1 => \N__28595\,
            in2 => \_gnd_net_\,
            in3 => \N__50326\,
            lcout => comm_buf_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51162\,
            ce => \N__25449\,
            sr => \N__20095\
        );

    \comm_buf_4__i6_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40732\,
            in1 => \N__20258\,
            in2 => \_gnd_net_\,
            in3 => \N__50327\,
            lcout => comm_buf_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51162\,
            ce => \N__25449\,
            sr => \N__20095\
        );

    \mux_1457_i8_4_lut_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__20126\,
            in1 => \N__48036\,
            in2 => \N__26003\,
            in3 => \N__47292\,
            lcout => OPEN,
            ltout => \n4057_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i7_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39383\,
            in1 => \_gnd_net_\,
            in2 => \N__20105\,
            in3 => \N__50328\,
            lcout => comm_buf_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51162\,
            ce => \N__25449\,
            sr => \N__20095\
        );

    \ADC_VAC1.ADC_DATA_i17_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53075\,
            in1 => \N__20056\,
            in2 => \N__20207\,
            in3 => \N__52888\,
            lcout => buf_adcdata1_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i18_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52879\,
            in1 => \N__53076\,
            in2 => \N__20041\,
            in3 => \N__20020\,
            lcout => buf_adcdata1_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i26_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20202\,
            in1 => \N__52883\,
            in2 => \N__20021\,
            in3 => \N__26158\,
            lcout => cmd_rdadctmp_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i27_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26159\,
            in1 => \N__20247\,
            in2 => \N__52898\,
            in3 => \N__20019\,
            lcout => cmd_rdadctmp_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i28_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20248\,
            in1 => \N__52884\,
            in2 => \N__20374\,
            in3 => \N__26160\,
            lcout => cmd_rdadctmp_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i19_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52880\,
            in1 => \N__53077\,
            in2 => \N__20227\,
            in3 => \N__20249\,
            lcout => buf_adcdata1_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i25_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__48259\,
            in1 => \N__52882\,
            in2 => \N__20206\,
            in3 => \N__26157\,
            lcout => cmd_rdadctmp_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i20_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52881\,
            in1 => \N__53078\,
            in2 => \N__20182\,
            in3 => \N__20370\,
            lcout => buf_adcdata1_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_140_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100001"
        )
    port map (
            in0 => \N__45659\,
            in1 => \N__47077\,
            in2 => \N__39556\,
            in3 => \N__40884\,
            lcout => n84,
            ltout => \n84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12632_2_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20162\,
            in3 => \N__34550\,
            lcout => OPEN,
            ltout => \n15593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__44178\,
            in1 => \N__50345\,
            in2 => \N__20159\,
            in3 => \N__26012\,
            lcout => comm_buf_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51198\,
            ce => \N__25274\,
            sr => \N__24209\
        );

    \i1_4_lut_adj_150_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101000"
        )
    port map (
            in0 => \N__40252\,
            in1 => \N__23867\,
            in2 => \N__27617\,
            in3 => \N__45220\,
            lcout => OPEN,
            ltout => \n8045_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i7_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__50344\,
            in1 => \N__20153\,
            in2 => \N__20156\,
            in3 => \N__39396\,
            lcout => comm_buf_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51198\,
            ce => \N__25274\,
            sr => \N__24209\
        );

    \i12650_2_lut_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38904\,
            in2 => \_gnd_net_\,
            in3 => \N__32094\,
            lcout => n15573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i11_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__44464\,
            in1 => \N__52837\,
            in2 => \N__20518\,
            in3 => \N__26177\,
            lcout => cmd_rdadctmp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i12_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25920\,
            in1 => \N__20481\,
            in2 => \N__22666\,
            in3 => \N__27464\,
            lcout => buf_adcdata4_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i8_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53697\,
            in1 => \N__20410\,
            in2 => \N__20459\,
            in3 => \N__53294\,
            lcout => buf_adcdata2_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i9_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20391\,
            in1 => \N__49240\,
            in2 => \N__43840\,
            in3 => \N__48816\,
            lcout => cmd_rdadctmp_9_adj_1103,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i29_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__20375\,
            in1 => \N__21288\,
            in2 => \N__52889\,
            in3 => \N__26178\,
            lcout => cmd_rdadctmp_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51215\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i9_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24144\,
            in1 => \N__22476\,
            in2 => \N__52891\,
            in3 => \N__26161\,
            lcout => cmd_rdadctmp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i17_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53716\,
            in1 => \N__20344\,
            in2 => \N__43966\,
            in3 => \N__53276\,
            lcout => buf_adcdata2_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i15_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__48776\,
            in1 => \N__21663\,
            in2 => \N__49204\,
            in3 => \N__20292\,
            lcout => cmd_rdadctmp_15_adj_1097,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i14_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20330\,
            in1 => \N__49124\,
            in2 => \N__20296\,
            in3 => \N__48777\,
            lcout => cmd_rdadctmp_14_adj_1098,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51232\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1457_i7_4_lut_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__20276\,
            in1 => \N__48074\,
            in2 => \N__24103\,
            in3 => \N__47311\,
            lcout => n4058,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_200_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001110"
        )
    port map (
            in0 => \N__23062\,
            in1 => \N__49107\,
            in2 => \N__20695\,
            in3 => \N__22978\,
            lcout => OPEN,
            ltout => \n14_adj_1031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.CS_37_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__49108\,
            in1 => \N__23123\,
            in2 => \N__20711\,
            in3 => \N__20723\,
            lcout => \M_CS3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i25_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__21327\,
            in1 => \N__46063\,
            in2 => \N__43962\,
            in3 => \N__53277\,
            lcout => cmd_rdadctmp_25_adj_1051,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i24_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__34475\,
            in1 => \N__46039\,
            in2 => \N__21331\,
            in3 => \N__53278\,
            lcout => cmd_rdadctmp_24_adj_1052,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.SCLK_35_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__49225\,
            in1 => \N__22979\,
            in2 => \N__20674\,
            in3 => \N__23058\,
            lcout => \M_SCLK3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i2_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20749\,
            in1 => \N__49226\,
            in2 => \N__21538\,
            in3 => \N__48734\,
            lcout => cmd_rdadctmp_2_adj_1110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i4_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__48733\,
            in1 => \N__21521\,
            in2 => \N__49256\,
            in3 => \N__20656\,
            lcout => cmd_rdadctmp_4_adj_1108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i5_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20657\,
            in1 => \N__49227\,
            in2 => \N__24286\,
            in3 => \N__48735\,
            lcout => cmd_rdadctmp_5_adj_1107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.DTRIG_39_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__20648\,
            in1 => \N__20585\,
            in2 => \N__52890\,
            in3 => \N__21482\,
            lcout => acadc_dtrig1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20758\,
            in1 => \N__49129\,
            in2 => \N__20780\,
            in3 => \N__48678\,
            lcout => cmd_rdadctmp_0_adj_1112,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i1_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20759\,
            in1 => \N__49130\,
            in2 => \N__20750\,
            in3 => \N__48679\,
            lcout => cmd_rdadctmp_1_adj_1111,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51279\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i13060_2_lut_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49128\,
            in2 => \_gnd_net_\,
            in3 => \N__22553\,
            lcout => \ADC_VAC3.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_32_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22956\,
            in2 => \_gnd_net_\,
            in3 => \N__23042\,
            lcout => n15147,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.adc_state_i2_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__49122\,
            in1 => \N__22955\,
            in2 => \_gnd_net_\,
            in3 => \N__23040\,
            lcout => \DTRIG_N_957_adj_1114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51292\,
            ce => \N__20735\,
            sr => \_gnd_net_\
        );

    \ADC_VAC3.adc_state_i1_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__49121\,
            in1 => \N__22954\,
            in2 => \_gnd_net_\,
            in3 => \N__23041\,
            lcout => adc_state_1_adj_1079,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51292\,
            ce => \N__20735\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_50_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22953\,
            in2 => \_gnd_net_\,
            in3 => \N__23039\,
            lcout => n15162,
            ltout => \n15162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i1_3_lut_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23111\,
            in2 => \N__20714\,
            in3 => \N__49120\,
            lcout => n8332,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_7322_7323_set_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28752\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n10433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42464\,
            ce => 'H',
            sr => \N__20876\
        );

    \comm_spi.RESET_I_0_98_2_lut_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46607\,
            lcout => \comm_spi.data_tx_7__N_811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13117_4_lut_3_lut_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46610\,
            in1 => \N__20923\,
            in2 => \_gnd_net_\,
            in3 => \N__21598\,
            lcout => \comm_spi.n16911\,
            ltout => \comm_spi.n16911_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_7348_7349_set_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20911\,
            in1 => \_gnd_net_\,
            in2 => \N__20900\,
            in3 => \N__21610\,
            lcout => \comm_spi.n10459\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42465\,
            ce => 'H',
            sr => \N__20897\
        );

    \comm_spi.RESET_I_0_106_2_lut_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20868\,
            lcout => \comm_spi.data_tx_7__N_831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_99_2_lut_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21597\,
            lcout => \comm_spi.data_tx_7__N_812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13082_4_lut_3_lut_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20870\,
            in1 => \N__23235\,
            in2 => \_gnd_net_\,
            in3 => \N__46609\,
            lcout => \comm_spi.n16908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_13249_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__20852\,
            in1 => \N__33330\,
            in2 => \N__20969\,
            in3 => \N__33176\,
            lcout => OPEN,
            ltout => \n16446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16446_bdd_4_lut_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33331\,
            in1 => \N__29102\,
            in2 => \N__20846\,
            in3 => \N__20843\,
            lcout => n16449,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1525_i4_4_lut_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__20831\,
            in1 => \N__48012\,
            in2 => \N__20818\,
            in3 => \N__47337\,
            lcout => n4305,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16428_bdd_4_lut_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__33175\,
            in1 => \N__24737\,
            in2 => \N__23261\,
            in3 => \N__21572\,
            lcout => n16431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13279_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__38825\,
            in1 => \N__23801\,
            in2 => \N__21860\,
            in3 => \N__33173\,
            lcout => OPEN,
            ltout => \n16506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16506_bdd_4_lut_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33174\,
            in1 => \N__21017\,
            in2 => \N__21005\,
            in3 => \N__21002\,
            lcout => n16509,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12214_3_lut_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38823\,
            in1 => \N__22151\,
            in2 => \_gnd_net_\,
            in3 => \N__23486\,
            lcout => n15424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12202_3_lut_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21914\,
            in1 => \N__23894\,
            in2 => \_gnd_net_\,
            in3 => \N__38821\,
            lcout => n15412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12240_3_lut_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38822\,
            in1 => \N__20960\,
            in2 => \_gnd_net_\,
            in3 => \N__20951\,
            lcout => n15450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13259_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__38824\,
            in1 => \N__25370\,
            in2 => \N__21983\,
            in3 => \N__33171\,
            lcout => OPEN,
            ltout => \n16482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16482_bdd_4_lut_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__33172\,
            in1 => \N__23342\,
            in2 => \N__20939\,
            in3 => \N__24824\,
            lcout => n16485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imiso_83_7340_7341_reset_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29128\,
            in1 => \N__29156\,
            in2 => \_gnd_net_\,
            in3 => \N__30845\,
            lcout => \comm_spi.n10452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_7340_7341_resetC_net\,
            ce => 'H',
            sr => \N__31007\
        );

    \comm_buf_3__i2_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40121\,
            in1 => \N__21137\,
            in2 => \_gnd_net_\,
            in3 => \N__49896\,
            lcout => comm_buf_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51140\,
            ce => \N__25175\,
            sr => \N__30736\
        );

    \comm_buf_3__i3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49895\,
            in1 => \N__44909\,
            in2 => \_gnd_net_\,
            in3 => \N__43001\,
            lcout => comm_buf_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51140\,
            ce => \N__25175\,
            sr => \N__30736\
        );

    \comm_buf_9__i3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44910\,
            in1 => \N__21104\,
            in2 => \_gnd_net_\,
            in3 => \N__50330\,
            lcout => comm_buf_9_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51150\,
            ce => \N__27707\,
            sr => \N__30743\
        );

    \comm_buf_9__i4_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50329\,
            in1 => \N__39940\,
            in2 => \_gnd_net_\,
            in3 => \N__21077\,
            lcout => comm_buf_9_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51150\,
            ce => \N__27707\,
            sr => \N__30743\
        );

    \i132_4_lut_adj_100_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100000001000"
        )
    port map (
            in0 => \N__48041\,
            in1 => \N__41258\,
            in2 => \N__45317\,
            in3 => \N__29581\,
            lcout => OPEN,
            ltout => \n66_adj_1153_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i123_3_lut_adj_105_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29300\,
            in2 => \N__21062\,
            in3 => \N__47268\,
            lcout => n96_adj_1159,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12672_2_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33752\,
            lcout => n15578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i20_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44351\,
            in1 => \N__49123\,
            in2 => \N__24251\,
            in3 => \N__24060\,
            lcout => buf_adcdata3_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.SCLK_27_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010011010001"
        )
    port map (
            in0 => \N__35765\,
            in1 => \N__48363\,
            in2 => \N__21046\,
            in3 => \N__48544\,
            lcout => \DDS_SCK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.MOSI_31_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31046\,
            in1 => \N__21214\,
            in2 => \_gnd_net_\,
            in3 => \N__48543\,
            lcout => \DDS_MOSI1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.bit_cnt_i0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__48545\,
            in1 => \N__25495\,
            in2 => \_gnd_net_\,
            in3 => \N__31189\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12726_2_lut_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48040\,
            in2 => \_gnd_net_\,
            in3 => \N__32216\,
            lcout => n15522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12666_2_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__31430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48042\,
            lcout => n15523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_13215_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__45219\,
            in1 => \N__21203\,
            in2 => \N__21197\,
            in3 => \N__47260\,
            lcout => OPEN,
            ltout => \n16398_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16398_bdd_4_lut_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47261\,
            in1 => \N__34046\,
            in2 => \N__21188\,
            in3 => \N__27749\,
            lcout => OPEN,
            ltout => \n16401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i108_4_lut_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__45660\,
            in1 => \N__34253\,
            in2 => \N__21185\,
            in3 => \N__47262\,
            lcout => OPEN,
            ltout => \n109_adj_1155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_123_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__31292\,
            in1 => \N__39543\,
            in2 => \N__21182\,
            in3 => \N__40251\,
            lcout => OPEN,
            ltout => \n8048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i5_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__39808\,
            in1 => \N__50323\,
            in2 => \N__21179\,
            in3 => \N__21176\,
            lcout => comm_buf_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51181\,
            ce => \N__25269\,
            sr => \N__24205\
        );

    \ADC_VAC1.ADC_DATA_i21_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52831\,
            in1 => \N__53127\,
            in2 => \N__21157\,
            in3 => \N__21290\,
            lcout => buf_adcdata1_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i22_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53126\,
            in1 => \N__52834\,
            in2 => \N__21355\,
            in3 => \N__21274\,
            lcout => buf_adcdata1_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i16_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53698\,
            in1 => \N__21304\,
            in2 => \N__21335\,
            in3 => \N__53293\,
            lcout => buf_adcdata2_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i31_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__26180\,
            in1 => \N__21273\,
            in2 => \N__22753\,
            in3 => \N__52835\,
            lcout => cmd_rdadctmp_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i30_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52832\,
            in1 => \N__21289\,
            in2 => \N__21275\,
            in3 => \N__26179\,
            lcout => cmd_rdadctmp_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53125\,
            in1 => \N__21250\,
            in2 => \N__24154\,
            in3 => \N__52833\,
            lcout => buf_adcdata1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.bit_cnt_i0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21383\,
            in2 => \_gnd_net_\,
            in3 => \N__21236\,
            lcout => \ADC_VAC2.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \ADC_VAC2.n13988\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21439\,
            in2 => \_gnd_net_\,
            in3 => \N__21233\,
            lcout => \ADC_VAC2.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC2.n13988\,
            carryout => \ADC_VAC2.n13989\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22601\,
            in2 => \_gnd_net_\,
            in3 => \N__21230\,
            lcout => \ADC_VAC2.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC2.n13989\,
            carryout => \ADC_VAC2.n13990\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22628\,
            in2 => \_gnd_net_\,
            in3 => \N__21227\,
            lcout => \ADC_VAC2.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC2.n13990\,
            carryout => \ADC_VAC2.n13991\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22640\,
            in2 => \_gnd_net_\,
            in3 => \N__21452\,
            lcout => \ADC_VAC2.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC2.n13991\,
            carryout => \ADC_VAC2.n13992\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22615\,
            in2 => \_gnd_net_\,
            in3 => \N__21449\,
            lcout => \ADC_VAC2.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC2.n13992\,
            carryout => \ADC_VAC2.n13993\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i6_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21397\,
            in2 => \_gnd_net_\,
            in3 => \N__21446\,
            lcout => \ADC_VAC2.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC2.n13993\,
            carryout => \ADC_VAC2.n13994\,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.bit_cnt_i7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21427\,
            in2 => \_gnd_net_\,
            in3 => \N__21443\,
            lcout => \ADC_VAC2.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51216\,
            ce => \N__36505\,
            sr => \N__36377\
        );

    \ADC_VAC2.i12780_4_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21440\,
            in1 => \N__21371\,
            in2 => \N__21428\,
            in3 => \N__22589\,
            lcout => \ADC_VAC2.n15595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i1_4_lut_adj_5_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__36456\,
            in1 => \N__53222\,
            in2 => \N__30214\,
            in3 => \N__30656\,
            lcout => OPEN,
            ltout => \ADC_VAC2.n15261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i1_2_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21413\,
            in3 => \N__35598\,
            lcout => \ADC_VAC2.n15262\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.adc_state_i0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__35599\,
            in1 => \N__53223\,
            in2 => \N__36470\,
            in3 => \N__21410\,
            lcout => adc_state_0_adj_1044,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51233\,
            ce => \N__21404\,
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i6_4_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__53221\,
            in1 => \N__35595\,
            in2 => \N__21398\,
            in3 => \N__21382\,
            lcout => \ADC_VAC2.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i30_4_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000110001"
        )
    port map (
            in0 => \N__35597\,
            in1 => \N__36434\,
            in2 => \N__30215\,
            in3 => \N__30657\,
            lcout => OPEN,
            ltout => \ADC_VAC2.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i13058_2_lut_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__53220\,
            in1 => \_gnd_net_\,
            in2 => \N__21542\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC2.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i1_4_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000110"
        )
    port map (
            in0 => \N__35596\,
            in1 => \N__36433\,
            in2 => \N__30213\,
            in3 => \N__53219\,
            lcout => \ADC_VAC2.n9413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i1_2_lut_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23057\,
            in2 => \_gnd_net_\,
            in3 => \N__22559\,
            lcout => \ADC_VAC3.n15260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.DTRIG_39_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011100000"
        )
    port map (
            in0 => \N__53275\,
            in1 => \N__35568\,
            in2 => \N__21502\,
            in3 => \N__36474\,
            lcout => acadc_dtrig2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i3_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21539\,
            in1 => \N__49012\,
            in2 => \N__21520\,
            in3 => \N__48757\,
            lcout => cmd_rdadctmp_3_adj_1109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_127_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21460\,
            in1 => \N__21469\,
            in2 => \N__21503\,
            in3 => \N__21481\,
            lcout => n14087,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.DTRIG_39_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101000"
        )
    port map (
            in0 => \N__21470\,
            in1 => \N__27115\,
            in2 => \N__27467\,
            in3 => \N__27034\,
            lcout => acadc_dtrig4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.DTRIG_39_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010101000"
        )
    port map (
            in0 => \N__21461\,
            in1 => \N__49231\,
            in2 => \N__22980\,
            in3 => \N__23049\,
            lcout => acadc_dtrig3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i6_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53063\,
            in1 => \N__21694\,
            in2 => \N__21734\,
            in3 => \N__52846\,
            lcout => buf_adcdata1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i18_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__46228\,
            in1 => \N__46072\,
            in2 => \N__38283\,
            in3 => \N__53325\,
            lcout => cmd_rdadctmp_18_adj_1058,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i16_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21676\,
            in1 => \N__49029\,
            in2 => \N__38193\,
            in3 => \N__48680\,
            lcout => cmd_rdadctmp_16_adj_1096,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.SCLK_35_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__27336\,
            in1 => \N__27116\,
            in2 => \N__21634\,
            in3 => \N__27035\,
            lcout => \M_SCLK4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51280\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_7322_7323_reset_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28751\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n10434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42463\,
            ce => 'H',
            sr => \N__21581\
        );

    \comm_spi.data_tx_i2_7352_7353_set_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23236\,
            in1 => \N__23215\,
            in2 => \_gnd_net_\,
            in3 => \N__23200\,
            lcout => \comm_spi.n10463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42448\,
            ce => 'H',
            sr => \N__24905\
        );

    \comm_spi.RESET_I_0_2_lut_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21599\,
            in2 => \_gnd_net_\,
            in3 => \N__46605\,
            lcout => \comm_spi.data_tx_7__N_834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13220_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23705\,
            in1 => \N__33170\,
            in2 => \N__21746\,
            in3 => \N__38837\,
            lcout => n16428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1469_i5_4_lut_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__21566\,
            in1 => \N__48083\,
            in2 => \N__24652\,
            in3 => \N__47293\,
            lcout => n4104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12172_3_lut_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21827\,
            in1 => \N__21818\,
            in2 => \_gnd_net_\,
            in3 => \N__38828\,
            lcout => OPEN,
            ltout => \n15382_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16380_bdd_4_lut_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__38582\,
            in1 => \N__21782\,
            in2 => \N__21806\,
            in3 => \N__33490\,
            lcout => OPEN,
            ltout => \n16383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i7_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33491\,
            in1 => \N__21797\,
            in2 => \N__21803\,
            in3 => \N__33346\,
            lcout => comm_tx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51114\,
            ce => \N__43139\,
            sr => \N__22384\
        );

    \comm_index_0__bdd_4_lut_13274_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33130\,
            in1 => \N__23930\,
            in2 => \N__21944\,
            in3 => \N__38827\,
            lcout => OPEN,
            ltout => \n16494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16494_bdd_4_lut_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__24764\,
            in1 => \N__33132\,
            in2 => \N__21800\,
            in3 => \N__23390\,
            lcout => n16497,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12241_3_lut_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21887\,
            in1 => \N__23588\,
            in2 => \_gnd_net_\,
            in3 => \N__38826\,
            lcout => OPEN,
            ltout => \n15451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_13177_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__21791\,
            in1 => \N__33131\,
            in2 => \N__21785\,
            in3 => \N__33489\,
            lcout => n16380,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_11__i1_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__50258\,
            in1 => \N__21776\,
            in2 => \_gnd_net_\,
            in3 => \N__44159\,
            lcout => comm_buf_11_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i2_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40118\,
            in1 => \N__21764\,
            in2 => \_gnd_net_\,
            in3 => \N__50264\,
            lcout => comm_buf_11_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i3_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50259\,
            in1 => \N__44887\,
            in2 => \_gnd_net_\,
            in3 => \N__22043\,
            lcout => comm_buf_11_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i4_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39928\,
            in1 => \N__22010\,
            in2 => \_gnd_net_\,
            in3 => \N__50265\,
            lcout => comm_buf_11_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i5_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50260\,
            in1 => \N__39804\,
            in2 => \_gnd_net_\,
            in3 => \N__21995\,
            lcout => comm_buf_11_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i6_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21974\,
            in1 => \N__50263\,
            in2 => \_gnd_net_\,
            in3 => \N__40706\,
            lcout => comm_buf_11_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i7_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50261\,
            in1 => \N__39394\,
            in2 => \_gnd_net_\,
            in3 => \N__21959\,
            lcout => comm_buf_11_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_11__i0_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21932\,
            in1 => \N__50262\,
            in2 => \_gnd_net_\,
            in3 => \N__39188\,
            lcout => comm_buf_11_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51120\,
            ce => \N__23837\,
            sr => \N__23822\
        );

    \comm_buf_7__i7_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49892\,
            in1 => \N__39395\,
            in2 => \_gnd_net_\,
            in3 => \N__21908\,
            lcout => comm_buf_7_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i0_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21878\,
            in1 => \N__49893\,
            in2 => \_gnd_net_\,
            in3 => \N__39205\,
            lcout => comm_buf_7_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i6_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49891\,
            in1 => \N__40730\,
            in2 => \_gnd_net_\,
            in3 => \N__21848\,
            lcout => comm_buf_7_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i5_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49898\,
            in1 => \N__22217\,
            in2 => \_gnd_net_\,
            in3 => \N__39803\,
            lcout => comm_buf_7_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i4_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49890\,
            in1 => \N__39915\,
            in2 => \_gnd_net_\,
            in3 => \N__22190\,
            lcout => comm_buf_7_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i3_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__49897\,
            in1 => \N__22169\,
            in2 => \_gnd_net_\,
            in3 => \N__44886\,
            lcout => comm_buf_7_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i2_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__49889\,
            in1 => \N__40120\,
            in2 => \_gnd_net_\,
            in3 => \N__22142\,
            lcout => comm_buf_7_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \comm_buf_7__i1_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44157\,
            in1 => \N__22112\,
            in2 => \_gnd_net_\,
            in3 => \N__49894\,
            lcout => comm_buf_7_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51128\,
            ce => \N__23855\,
            sr => \N__23846\
        );

    \i12193_3_lut_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38836\,
            in1 => \N__22076\,
            in2 => \_gnd_net_\,
            in3 => \N__22061\,
            lcout => OPEN,
            ltout => \n15403_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16476_bdd_4_lut_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__29339\,
            in1 => \N__22244\,
            in2 => \N__22049\,
            in3 => \N__33484\,
            lcout => OPEN,
            ltout => \n16479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i4_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__33485\,
            in1 => \N__22283\,
            in2 => \N__22046\,
            in3 => \N__33321\,
            lcout => comm_tx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51141\,
            ce => \N__43109\,
            sr => \N__22385\
        );

    \i12190_3_lut_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22307\,
            in1 => \N__23510\,
            in2 => \_gnd_net_\,
            in3 => \N__38833\,
            lcout => n15400,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13244_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__38835\,
            in1 => \N__22301\,
            in2 => \N__23960\,
            in3 => \N__33177\,
            lcout => OPEN,
            ltout => \n16452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16452_bdd_4_lut_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__23318\,
            in1 => \N__22292\,
            in2 => \N__22286\,
            in3 => \N__33179\,
            lcout => n16455,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12189_3_lut_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38834\,
            in1 => \N__22277\,
            in2 => \_gnd_net_\,
            in3 => \N__22262\,
            lcout => OPEN,
            ltout => \n15399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__22253\,
            in1 => \N__33483\,
            in2 => \N__22247\,
            in3 => \N__33178\,
            lcout => n16476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12674_2_lut_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48039\,
            in2 => \_gnd_net_\,
            in3 => \N__34037\,
            lcout => OPEN,
            ltout => \n15633_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_13269_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__22424\,
            in1 => \N__45309\,
            in2 => \N__22238\,
            in3 => \N__47272\,
            lcout => OPEN,
            ltout => \n16458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16458_bdd_4_lut_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47273\,
            in1 => \N__29198\,
            in2 => \N__22235\,
            in3 => \N__28013\,
            lcout => OPEN,
            ltout => \n16461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_117_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110100"
        )
    port map (
            in0 => \N__39568\,
            in1 => \N__24038\,
            in2 => \N__22232\,
            in3 => \N__45654\,
            lcout => OPEN,
            ltout => \n76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_118_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__36960\,
            in1 => \N__22541\,
            in2 => \N__22430\,
            in3 => \N__40253\,
            lcout => OPEN,
            ltout => \n4_adj_1195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i4_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__36887\,
            in1 => \N__39922\,
            in2 => \N__22427\,
            in3 => \N__50291\,
            lcout => comm_buf_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51151\,
            ce => \N__25266\,
            sr => \N__24192\
        );

    \i12816_2_lut_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48038\,
            in2 => \_gnd_net_\,
            in3 => \N__30062\,
            lcout => n15632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i2_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__22418\,
            in1 => \N__40053\,
            in2 => \N__50324\,
            in3 => \N__22400\,
            lcout => comm_buf_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51164\,
            ce => \N__25268\,
            sr => \N__24186\
        );

    \i127_4_lut_adj_96_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__47254\,
            in1 => \N__27887\,
            in2 => \N__36734\,
            in3 => \N__45647\,
            lcout => n130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12699_2_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34373\,
            in2 => \_gnd_net_\,
            in3 => \N__32108\,
            lcout => n15589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i131_3_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26458\,
            in1 => \N__34819\,
            in2 => \_gnd_net_\,
            in3 => \N__47255\,
            lcout => OPEN,
            ltout => \n87_adj_1165_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i124_4_lut_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__47256\,
            in1 => \N__26257\,
            in2 => \N__22412\,
            in3 => \N__45648\,
            lcout => OPEN,
            ltout => \n69_adj_1161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_97_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__39542\,
            in1 => \N__40241\,
            in2 => \N__22409\,
            in3 => \N__22406\,
            lcout => n8050,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_116_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__45661\,
            in1 => \N__39569\,
            in2 => \N__47315\,
            in3 => \N__40886\,
            lcout => n8089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12691_2_lut_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43532\,
            in2 => \_gnd_net_\,
            in3 => \N__32118\,
            lcout => n15587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i127_4_lut_adj_107_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__45662\,
            in1 => \N__40565\,
            in2 => \N__22532\,
            in3 => \N__47274\,
            lcout => OPEN,
            ltout => \n130_adj_1156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_110_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__39570\,
            in1 => \N__40211\,
            in2 => \N__22520\,
            in3 => \N__24113\,
            lcout => OPEN,
            ltout => \n8051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i3_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__44917\,
            in1 => \N__22517\,
            in2 => \N__22511\,
            in3 => \N__50343\,
            lcout => comm_buf_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51182\,
            ce => \N__25270\,
            sr => \N__24193\
        );

    \ADC_VAC4.ADC_DATA_i11_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25897\,
            in1 => \N__26541\,
            in2 => \N__22508\,
            in3 => \N__27380\,
            lcout => buf_adcdata4_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i22_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__37461\,
            in1 => \N__52875\,
            in2 => \N__44602\,
            in3 => \N__26162\,
            lcout => cmd_rdadctmp_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i23_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__26163\,
            in1 => \N__37462\,
            in2 => \N__22710\,
            in3 => \N__52877\,
            lcout => cmd_rdadctmp_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53123\,
            in1 => \N__22444\,
            in2 => \N__22478\,
            in3 => \N__52876\,
            lcout => buf_adcdata1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i15_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__52874\,
            in1 => \N__53124\,
            in2 => \N__22711\,
            in3 => \N__22684\,
            lcout => buf_adcdata1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i21_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__26404\,
            in1 => \N__27379\,
            in2 => \N__22670\,
            in3 => \N__26850\,
            lcout => cmd_rdadctmp_21_adj_1128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i12926_4_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__22639\,
            in1 => \N__22627\,
            in2 => \N__22616\,
            in3 => \N__22600\,
            lcout => \ADC_VAC2.n15596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i12127_4_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22819\,
            in1 => \N__22834\,
            in2 => \N__22868\,
            in3 => \N__22849\,
            lcout => OPEN,
            ltout => \ADC_VAC3.n15334_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i12149_4_lut_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22789\,
            in1 => \N__22882\,
            in2 => \N__22583\,
            in3 => \N__22771\,
            lcout => OPEN,
            ltout => \ADC_VAC3.n15358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i12787_4_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23066\,
            in1 => \N__22804\,
            in2 => \N__22580\,
            in3 => \N__49007\,
            lcout => OPEN,
            ltout => \ADC_VAC3.n15602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.adc_state_i0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__22983\,
            in1 => \N__23067\,
            in2 => \N__22577\,
            in3 => \N__48943\,
            lcout => adc_state_0_adj_1080,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51217\,
            ce => \N__22574\,
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i1_4_lut_adj_7_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__22982\,
            in1 => \N__48942\,
            in2 => \N__23129\,
            in3 => \N__30654\,
            lcout => \ADC_VAC3.n15259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i30_4_lut_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110000001"
        )
    port map (
            in0 => \N__30655\,
            in1 => \N__22981\,
            in2 => \N__23069\,
            in3 => \N__23128\,
            lcout => \ADC_VAC3.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.bit_cnt_i0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22883\,
            in2 => \_gnd_net_\,
            in3 => \N__22871\,
            lcout => \ADC_VAC3.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \ADC_VAC3.n13995\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22867\,
            in2 => \_gnd_net_\,
            in3 => \N__22853\,
            lcout => \ADC_VAC3.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC3.n13995\,
            carryout => \ADC_VAC3.n13996\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22850\,
            in2 => \_gnd_net_\,
            in3 => \N__22838\,
            lcout => \ADC_VAC3.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC3.n13996\,
            carryout => \ADC_VAC3.n13997\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i3_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22835\,
            in2 => \_gnd_net_\,
            in3 => \N__22823\,
            lcout => \ADC_VAC3.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC3.n13997\,
            carryout => \ADC_VAC3.n13998\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i4_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22820\,
            in2 => \_gnd_net_\,
            in3 => \N__22808\,
            lcout => \ADC_VAC3.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC3.n13998\,
            carryout => \ADC_VAC3.n13999\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i5_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22805\,
            in2 => \_gnd_net_\,
            in3 => \N__22793\,
            lcout => \ADC_VAC3.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC3.n13999\,
            carryout => \ADC_VAC3.n14000\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i6_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22790\,
            in2 => \_gnd_net_\,
            in3 => \N__22778\,
            lcout => \ADC_VAC3.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC3.n14000\,
            carryout => \ADC_VAC3.n14001\,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC3.bit_cnt_i7_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22772\,
            in2 => \_gnd_net_\,
            in3 => \N__22775\,
            lcout => \ADC_VAC3.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51234\,
            ce => \N__22991\,
            sr => \N__22913\
        );

    \ADC_VAC1.ADC_DATA_i23_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53064\,
            in1 => \N__22729\,
            in2 => \N__22760\,
            in3 => \N__52844\,
            lcout => buf_adcdata1_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51250\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i1_4_lut_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000100"
        )
    port map (
            in0 => \N__49020\,
            in1 => \N__22984\,
            in2 => \N__23124\,
            in3 => \N__23068\,
            lcout => \ADC_VAC3.n9514\,
            ltout => \ADC_VAC3.n9514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.i7638_2_lut_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__22985\,
            in1 => \_gnd_net_\,
            in2 => \N__22916\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC3.n10744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_67_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27105\,
            in2 => \_gnd_net_\,
            in3 => \N__27033\,
            lcout => n15144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.bit_cnt_i0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24413\,
            in2 => \_gnd_net_\,
            in3 => \N__22901\,
            lcout => \ADC_VAC4.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \ADC_VAC4.n14002\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i1_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24454\,
            in2 => \_gnd_net_\,
            in3 => \N__22898\,
            lcout => \ADC_VAC4.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC4.n14002\,
            carryout => \ADC_VAC4.n14003\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i2_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24440\,
            in2 => \_gnd_net_\,
            in3 => \N__22895\,
            lcout => \ADC_VAC4.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC4.n14003\,
            carryout => \ADC_VAC4.n14004\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i3_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24467\,
            in2 => \_gnd_net_\,
            in3 => \N__22892\,
            lcout => \ADC_VAC4.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC4.n14004\,
            carryout => \ADC_VAC4.n14005\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i4_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24479\,
            in2 => \_gnd_net_\,
            in3 => \N__22889\,
            lcout => \ADC_VAC4.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC4.n14005\,
            carryout => \ADC_VAC4.n14006\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i5_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24691\,
            in2 => \_gnd_net_\,
            in3 => \N__22886\,
            lcout => \ADC_VAC4.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC4.n14006\,
            carryout => \ADC_VAC4.n14007\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i6_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24427\,
            in2 => \_gnd_net_\,
            in3 => \N__23246\,
            lcout => \ADC_VAC4.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC4.n14007\,
            carryout => \ADC_VAC4.n14008\,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.bit_cnt_i7_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24398\,
            in2 => \_gnd_net_\,
            in3 => \N__23243\,
            lcout => \ADC_VAC4.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51267\,
            ce => \N__24668\,
            sr => \N__24659\
        );

    \ADC_VAC4.ADC_DATA_i22_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25961\,
            in1 => \N__29061\,
            in2 => \N__23438\,
            in3 => \N__27352\,
            lcout => buf_adcdata4_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i2_7352_7353_reset_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23240\,
            in1 => \N__23219\,
            in2 => \_gnd_net_\,
            in3 => \N__23204\,
            lcout => \comm_spi.n10464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42455\,
            ce => 'H',
            sr => \N__23186\
        );

    \ADC_VAC4.ADC_DATA_i19_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25942\,
            in1 => \N__43017\,
            in2 => \N__25655\,
            in3 => \N__27524\,
            lcout => buf_adcdata4_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_105_2_lut_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46604\,
            in2 => \_gnd_net_\,
            in3 => \N__24928\,
            lcout => \comm_spi.data_tx_7__N_828\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i21_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25943\,
            in1 => \N__23166\,
            in2 => \N__23144\,
            in3 => \N__27525\,
            lcout => buf_adcdata4_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i29_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26851\,
            in1 => \N__23139\,
            in2 => \N__27529\,
            in3 => \N__25624\,
            lcout => cmd_rdadctmp_29_adj_1120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i30_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__23140\,
            in1 => \N__27517\,
            in2 => \N__23434\,
            in3 => \N__26853\,
            lcout => cmd_rdadctmp_30_adj_1119,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i31_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26852\,
            in1 => \N__23413\,
            in2 => \N__27530\,
            in3 => \N__23430\,
            lcout => cmd_rdadctmp_31_adj_1118,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i23_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27516\,
            in1 => \N__25944\,
            in2 => \N__45867\,
            in3 => \N__23414\,
            lcout => buf_adcdata4_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51109\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_8__i7_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50316\,
            in1 => \N__39334\,
            in2 => \_gnd_net_\,
            in3 => \N__23405\,
            lcout => comm_buf_8_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i6_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23381\,
            in1 => \N__40691\,
            in2 => \_gnd_net_\,
            in3 => \N__50320\,
            lcout => comm_buf_8_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i5_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50315\,
            in1 => \_gnd_net_\,
            in2 => \N__39795\,
            in3 => \N__23357\,
            lcout => comm_buf_8_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i4_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39859\,
            in1 => \N__23333\,
            in2 => \_gnd_net_\,
            in3 => \N__50319\,
            lcout => comm_buf_8_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50314\,
            in1 => \N__44856\,
            in2 => \_gnd_net_\,
            in3 => \N__23306\,
            lcout => comm_buf_8_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i2_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23273\,
            in1 => \N__40076\,
            in2 => \_gnd_net_\,
            in3 => \N__50318\,
            lcout => comm_buf_8_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50313\,
            in1 => \N__44099\,
            in2 => \_gnd_net_\,
            in3 => \N__23660\,
            lcout => comm_buf_8_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_8__i0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23633\,
            in1 => \N__50317\,
            in2 => \_gnd_net_\,
            in3 => \N__39177\,
            lcout => comm_buf_8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51112\,
            ce => \N__25082\,
            sr => \N__25067\
        );

    \comm_buf_6__i7_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39390\,
            in1 => \N__23603\,
            in2 => \_gnd_net_\,
            in3 => \N__50257\,
            lcout => comm_buf_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51115\,
            ce => \N__23762\,
            sr => \N__23743\
        );

    \comm_buf_6__i6_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50254\,
            in1 => \_gnd_net_\,
            in2 => \N__40722\,
            in3 => \N__23582\,
            lcout => comm_buf_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51115\,
            ce => \N__23762\,
            sr => \N__23743\
        );

    \comm_buf_6__i5_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39785\,
            in1 => \N__23552\,
            in2 => \_gnd_net_\,
            in3 => \N__50256\,
            lcout => comm_buf_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51115\,
            ce => \N__23762\,
            sr => \N__23743\
        );

    \comm_buf_6__i4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50253\,
            in1 => \N__39887\,
            in2 => \_gnd_net_\,
            in3 => \N__23525\,
            lcout => comm_buf_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51115\,
            ce => \N__23762\,
            sr => \N__23743\
        );

    \comm_buf_6__i3_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__44885\,
            in2 => \_gnd_net_\,
            in3 => \N__50255\,
            lcout => comm_buf_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51115\,
            ce => \N__23762\,
            sr => \N__23743\
        );

    \comm_buf_6__i2_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50252\,
            in1 => \N__40117\,
            in2 => \_gnd_net_\,
            in3 => \N__23474\,
            lcout => comm_buf_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51115\,
            ce => \N__23762\,
            sr => \N__23743\
        );

    \i1_4_lut_adj_237_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__38787\,
            in1 => \N__42798\,
            in2 => \N__38559\,
            in3 => \N__25399\,
            lcout => n8907,
            ltout => \n8907_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7512_2_lut_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23858\,
            in3 => \N__52450\,
            lcout => n10618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_247_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__38788\,
            in1 => \N__42799\,
            in2 => \N__38560\,
            in3 => \N__25400\,
            lcout => n8943,
            ltout => \n8943_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7519_2_lut_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23849\,
            in3 => \N__52451\,
            lcout => n10625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_275_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__38789\,
            in1 => \N__42800\,
            in2 => \N__38561\,
            in3 => \N__25154\,
            lcout => n9123,
            ltout => \n9123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7547_2_lut_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23825\,
            in3 => \N__52452\,
            lcout => n10653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39179\,
            in1 => \N__23816\,
            in2 => \_gnd_net_\,
            in3 => \N__50312\,
            lcout => comm_buf_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51121\,
            ce => \N__23761\,
            sr => \N__23744\
        );

    \comm_buf_6__i1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50311\,
            in1 => \N__44156\,
            in2 => \_gnd_net_\,
            in3 => \N__23789\,
            lcout => comm_buf_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51121\,
            ce => \N__23761\,
            sr => \N__23744\
        );

    \comm_buf_10__i2_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40119\,
            in1 => \N__23723\,
            in2 => \_gnd_net_\,
            in3 => \N__50303\,
            lcout => comm_buf_10_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51129\,
            ce => \N__25356\,
            sr => \N__25319\
        );

    \comm_buf_10__i3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50300\,
            in1 => \N__44888\,
            in2 => \_gnd_net_\,
            in3 => \N__23693\,
            lcout => comm_buf_10_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51129\,
            ce => \N__25356\,
            sr => \N__25319\
        );

    \comm_buf_10__i4_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39914\,
            in1 => \N__23978\,
            in2 => \_gnd_net_\,
            in3 => \N__50304\,
            lcout => comm_buf_10_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51129\,
            ce => \N__25356\,
            sr => \N__25319\
        );

    \comm_buf_10__i7_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50301\,
            in1 => \_gnd_net_\,
            in2 => \N__39401\,
            in3 => \N__23951\,
            lcout => comm_buf_10_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51129\,
            ce => \N__25356\,
            sr => \N__25319\
        );

    \comm_buf_10__i0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39180\,
            in1 => \N__23915\,
            in2 => \_gnd_net_\,
            in3 => \N__50302\,
            lcout => comm_buf_10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51129\,
            ce => \N__25356\,
            sr => \N__25319\
        );

    \comm_cmd_1__bdd_4_lut_13235_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__28052\,
            in1 => \N__45289\,
            in2 => \N__31307\,
            in3 => \N__47251\,
            lcout => OPEN,
            ltout => \n16434_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16434_bdd_4_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47252\,
            in1 => \N__27980\,
            in2 => \N__23882\,
            in3 => \N__29168\,
            lcout => OPEN,
            ltout => \n16437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i108_4_lut_adj_132_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__30902\,
            in1 => \N__45538\,
            in2 => \N__23879\,
            in3 => \N__47253\,
            lcout => n109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_136_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__23876\,
            in1 => \N__42968\,
            in2 => \N__39581\,
            in3 => \N__40240\,
            lcout => OPEN,
            ltout => \n8054_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__40731\,
            in1 => \N__27758\,
            in2 => \N__23870\,
            in3 => \N__50305\,
            lcout => comm_buf_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51142\,
            ce => \N__25265\,
            sr => \N__24187\
        );

    \i106_4_lut_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__47921\,
            in1 => \N__25757\,
            in2 => \N__41633\,
            in3 => \N__45646\,
            lcout => n59,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i16_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44359\,
            in1 => \N__49110\,
            in2 => \N__28493\,
            in3 => \N__26355\,
            lcout => buf_adcdata3_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51152\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i17_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49109\,
            in1 => \N__44360\,
            in2 => \N__24014\,
            in3 => \N__27954\,
            lcout => buf_adcdata3_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51152\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i25_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__28489\,
            in1 => \N__24009\,
            in2 => \N__48831\,
            in3 => \N__49111\,
            lcout => cmd_rdadctmp_25_adj_1087,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51152\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i26_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__24010\,
            in1 => \N__48805\,
            in2 => \N__49202\,
            in3 => \N__26481\,
            lcout => cmd_rdadctmp_26_adj_1086,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51152\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7470_2_lut_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52453\,
            in2 => \_gnd_net_\,
            in3 => \N__25224\,
            lcout => n10576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i7_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__48824\,
            in1 => \N__24269\,
            in2 => \N__49203\,
            in3 => \N__23992\,
            lcout => cmd_rdadctmp_7_adj_1105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51152\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i27_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__26847\,
            in1 => \N__25741\,
            in2 => \N__25651\,
            in3 => \N__27466\,
            lcout => cmd_rdadctmp_27_adj_1122,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51152\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_13289_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__26432\,
            in1 => \N__45308\,
            in2 => \N__31394\,
            in3 => \N__47247\,
            lcout => OPEN,
            ltout => \n16500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16500_bdd_4_lut_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47248\,
            in1 => \N__27995\,
            in2 => \N__23981\,
            in3 => \N__27971\,
            lcout => OPEN,
            ltout => \n16503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_293_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__31349\,
            in1 => \N__45657\,
            in2 => \N__24221\,
            in3 => \N__47249\,
            lcout => n4_adj_1280,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_295_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__40210\,
            in1 => \N__24218\,
            in2 => \N__39580\,
            in3 => \N__24386\,
            lcout => OPEN,
            ltout => \n8047_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__39201\,
            in1 => \N__32069\,
            in2 => \N__24212\,
            in3 => \N__50342\,
            lcout => comm_buf_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51165\,
            ce => \N__25267\,
            sr => \N__24188\
        );

    \ADC_VAC1.cmd_rdadctmp_i10_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24155\,
            in1 => \N__52813\,
            in2 => \N__44451\,
            in3 => \N__26182\,
            lcout => cmd_rdadctmp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_3__358_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__39650\,
            in1 => \N__43533\,
            in2 => \N__24128\,
            in3 => \N__41169\,
            lcout => buf_control_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i124_4_lut_adj_108_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__26192\,
            in1 => \N__45658\,
            in2 => \N__24127\,
            in3 => \N__47250\,
            lcout => n69_adj_1029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i14_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25882\,
            in1 => \N__24096\,
            in2 => \N__27353\,
            in3 => \N__26392\,
            lcout => buf_adcdata4_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i112_4_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__24074\,
            in1 => \N__45655\,
            in2 => \N__24026\,
            in3 => \N__47243\,
            lcout => n61,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_4__357_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__41171\,
            in1 => \N__39655\,
            in2 => \N__36989\,
            in3 => \N__24025\,
            lcout => buf_control_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i127_4_lut_adj_294_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__26333\,
            in1 => \N__45656\,
            in2 => \N__24376\,
            in3 => \N__47244\,
            lcout => n69,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_0__361_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__39654\,
            in1 => \N__34118\,
            in2 => \N__24377\,
            in3 => \N__41170\,
            lcout => buf_control_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i28_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__48978\,
            in1 => \N__24237\,
            in2 => \N__25708\,
            in3 => \N__48785\,
            lcout => cmd_rdadctmp_28_adj_1084,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i9_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__34590\,
            in1 => \N__29227\,
            in2 => \N__41527\,
            in3 => \N__41380\,
            lcout => buf_dds_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i27_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__48977\,
            in1 => \N__26488\,
            in2 => \N__25707\,
            in3 => \N__48784\,
            lcout => cmd_rdadctmp_27_adj_1085,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1457_i1_4_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__24362\,
            in1 => \N__48004\,
            in2 => \N__24346\,
            in3 => \N__47246\,
            lcout => n4064,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i6_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__48755\,
            in1 => \N__24262\,
            in2 => \N__24290\,
            in3 => \N__49011\,
            lcout => cmd_rdadctmp_6_adj_1106,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i29_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__24244\,
            in1 => \N__36861\,
            in2 => \N__49119\,
            in3 => \N__48756\,
            lcout => cmd_rdadctmp_29_adj_1083,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i13_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27288\,
            in1 => \N__25883\,
            in2 => \N__26420\,
            in3 => \N__28616\,
            lcout => buf_adcdata4_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i17_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__32173\,
            in1 => \N__52809\,
            in2 => \N__24575\,
            in3 => \N__26183\,
            lcout => cmd_rdadctmp_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i19_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__26184\,
            in1 => \N__24552\,
            in2 => \N__52878\,
            in3 => \N__52917\,
            lcout => cmd_rdadctmp_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51218\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i9_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52795\,
            in1 => \N__53085\,
            in2 => \N__24595\,
            in3 => \N__24574\,
            lcout => buf_adcdata1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i18_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__52796\,
            in1 => \N__24573\,
            in2 => \N__52921\,
            in3 => \N__26185\,
            lcout => cmd_rdadctmp_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i20_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__52797\,
            in1 => \N__46272\,
            in2 => \N__24557\,
            in3 => \N__26186\,
            lcout => cmd_rdadctmp_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i11_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53084\,
            in1 => \N__52798\,
            in2 => \N__24532\,
            in3 => \N__24556\,
            lcout => buf_adcdata1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i8_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44302\,
            in1 => \N__49118\,
            in2 => \N__38207\,
            in3 => \N__24501\,
            lcout => buf_adcdata3_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51235\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i12123_4_lut_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24478\,
            in1 => \N__24466\,
            in2 => \N__24455\,
            in3 => \N__24439\,
            lcout => OPEN,
            ltout => \ADC_VAC4.n15330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i12146_4_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24428\,
            in1 => \N__24412\,
            in2 => \N__24401\,
            in3 => \N__24397\,
            lcout => \ADC_VAC4.n15354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i12804_4_lut_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27250\,
            in1 => \N__27009\,
            in2 => \N__24692\,
            in3 => \N__24677\,
            lcout => OPEN,
            ltout => \ADC_VAC4.n15619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.adc_state_i0_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__27010\,
            in1 => \N__27251\,
            in2 => \N__24671\,
            in3 => \N__27110\,
            lcout => adc_state_0_adj_1117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51251\,
            ce => \N__26681\,
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i30_4_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001010001"
        )
    port map (
            in0 => \N__27109\,
            in1 => \N__27008\,
            in2 => \N__26669\,
            in3 => \N__30647\,
            lcout => \ADC_VAC4.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i1_4_lut_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000100"
        )
    port map (
            in0 => \N__27238\,
            in1 => \N__27111\,
            in2 => \N__26665\,
            in3 => \N__27007\,
            lcout => \ADC_VAC4.n9631\,
            ltout => \ADC_VAC4.n9631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i7677_2_lut_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__27112\,
            in1 => \_gnd_net_\,
            in2 => \N__24662\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC4.n10783\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i20_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25960\,
            in1 => \N__24639\,
            in2 => \N__25625\,
            in3 => \N__27489\,
            lcout => buf_adcdata4_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_96_2_lut_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30954\,
            lcout => \comm_spi.data_tx_7__N_809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13092_4_lut_3_lut_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24935\,
            in1 => \N__24889\,
            in2 => \_gnd_net_\,
            in3 => \N__46603\,
            lcout => \comm_spi.n16905\,
            ltout => \comm_spi.n16905_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_7356_7357_set_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24871\,
            in2 => \N__24617\,
            in3 => \N__24853\,
            lcout => \comm_spi.n10467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42447\,
            ce => 'H',
            sr => \N__24614\
        );

    \comm_spi.RESET_I_0_97_2_lut_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24934\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46602\,
            lcout => \comm_spi.data_tx_7__N_810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_103_2_lut_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46640\,
            in2 => \_gnd_net_\,
            in3 => \N__46600\,
            lcout => \comm_spi.data_tx_7__N_822\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_7356_7357_reset_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24890\,
            in1 => \N__24878\,
            in2 => \_gnd_net_\,
            in3 => \N__24854\,
            lcout => \comm_spi.n10468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42459\,
            ce => 'H',
            sr => \N__30932\
        );

    \comm_buf_9__i5_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39766\,
            in1 => \N__24842\,
            in2 => \_gnd_net_\,
            in3 => \N__50309\,
            lcout => comm_buf_9_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51108\,
            ce => \N__25031\,
            sr => \N__25012\
        );

    \comm_buf_9__i6_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50307\,
            in1 => \N__40690\,
            in2 => \_gnd_net_\,
            in3 => \N__24812\,
            lcout => comm_buf_9_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51108\,
            ce => \N__25031\,
            sr => \N__25012\
        );

    \comm_buf_9__i7_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39333\,
            in1 => \N__24782\,
            in2 => \_gnd_net_\,
            in3 => \N__50310\,
            lcout => comm_buf_9_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51108\,
            ce => \N__25031\,
            sr => \N__25012\
        );

    \comm_buf_9__i2_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50306\,
            in1 => \N__40075\,
            in2 => \_gnd_net_\,
            in3 => \N__24755\,
            lcout => comm_buf_9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51108\,
            ce => \N__25031\,
            sr => \N__25012\
        );

    \comm_buf_9__i1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44098\,
            in1 => \N__24725\,
            in2 => \_gnd_net_\,
            in3 => \N__50308\,
            lcout => comm_buf_9_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51108\,
            ce => \N__25031\,
            sr => \N__25012\
        );

    \i7533_2_lut_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52385\,
            in2 => \_gnd_net_\,
            in3 => \N__25029\,
            lcout => n10639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_231_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__50601\,
            in1 => \N__33294\,
            in2 => \N__33488\,
            in3 => \N__27861\,
            lcout => n13470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_234_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__27862\,
            in1 => \N__25192\,
            in2 => \N__33328\,
            in3 => \N__33460\,
            lcout => OPEN,
            ltout => \n15161_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_268_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__50602\,
            in1 => \N__38534\,
            in2 => \N__25085\,
            in3 => \N__42795\,
            lcout => n9027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_255_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__42796\,
            in1 => \N__25421\,
            in2 => \N__38548\,
            in3 => \N__25166\,
            lcout => n8997,
            ltout => \n8997_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7526_2_lut_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__52386\,
            in1 => \_gnd_net_\,
            in2 => \N__25070\,
            in3 => \_gnd_net_\,
            lcout => n10632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_429_i6_2_lut_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__33295\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33459\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_9__i0_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25061\,
            in1 => \N__50266\,
            in2 => \_gnd_net_\,
            in3 => \N__39178\,
            lcout => comm_buf_9_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51111\,
            ce => \N__25030\,
            sr => \N__25013\
        );

    \comm_index_0__bdd_4_lut_13210_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__33102\,
            in1 => \N__24941\,
            in2 => \N__24995\,
            in3 => \N__38785\,
            lcout => n16422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_10__i1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50215\,
            in1 => \N__44151\,
            in2 => \_gnd_net_\,
            in3 => \N__24965\,
            lcout => comm_buf_10_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51113\,
            ce => \N__25357\,
            sr => \N__25317\
        );

    \i12638_2_lut_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33100\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38784\,
            lcout => n15670,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_243_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__52449\,
            in1 => \N__31055\,
            in2 => \N__51928\,
            in3 => \N__31124\,
            lcout => n8763,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_273_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33101\,
            in2 => \_gnd_net_\,
            in3 => \N__25165\,
            lcout => n13497,
            ltout => \n13497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_269_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__38558\,
            in1 => \N__38786\,
            in2 => \N__25148\,
            in3 => \N__42797\,
            lcout => n9045,
            ltout => \n9045_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7540_2_lut_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25145\,
            in3 => \N__52448\,
            lcout => n10646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_13264_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__25094\,
            in1 => \N__33097\,
            in2 => \N__25142\,
            in3 => \N__38781\,
            lcout => n16488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_10__i6_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50201\,
            in1 => \_gnd_net_\,
            in2 => \N__25115\,
            in3 => \N__40723\,
            lcout => comm_buf_10_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51118\,
            ce => \N__25355\,
            sr => \N__25313\
        );

    \i1_3_lut_4_lut_adj_260_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__50597\,
            in1 => \N__33249\,
            in2 => \N__33449\,
            in3 => \N__27856\,
            lcout => n13457,
            ltout => \n13457_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12761_2_lut_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25088\,
            in3 => \N__25417\,
            lcout => OPEN,
            ltout => \n15565_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i20_4_lut_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__50598\,
            in1 => \N__50200\,
            in2 => \N__25463\,
            in3 => \N__33626\,
            lcout => OPEN,
            ltout => \n13_adj_1257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_219_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25581\,
            in2 => \N__25460\,
            in3 => \N__42856\,
            lcout => n8823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i61_2_lut_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33096\,
            in2 => \_gnd_net_\,
            in3 => \N__38780\,
            lcout => n41,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_245_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25406\,
            lcout => n13458,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_10__i5_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50211\,
            in1 => \_gnd_net_\,
            in2 => \N__39802\,
            in3 => \N__25391\,
            lcout => comm_buf_10_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51125\,
            ce => \N__25358\,
            sr => \N__25318\
        );

    \equal_436_i5_2_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33099\,
            in2 => \_gnd_net_\,
            in3 => \N__38782\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_256_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__38783\,
            in1 => \N__33103\,
            in2 => \N__50322\,
            in3 => \N__31074\,
            lcout => OPEN,
            ltout => \n11_adj_1279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_142_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__42862\,
            in1 => \N__25582\,
            in2 => \N__25277\,
            in3 => \N__50599\,
            lcout => n8654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i36_4_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__50210\,
            in1 => \N__37079\,
            in2 => \N__25196\,
            in3 => \N__31075\,
            lcout => OPEN,
            ltout => \n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_179_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__42863\,
            in1 => \N__25583\,
            in2 => \N__25532\,
            in3 => \N__50600\,
            lcout => n8702,
            ltout => \n8702_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7477_2_lut_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25529\,
            in3 => \N__52376\,
            lcout => n10583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.i4_4_lut_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25525\,
            in1 => \N__25515\,
            in2 => \N__25504\,
            in3 => \N__48381\,
            lcout => n10_adj_1172,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.bit_cnt_i3_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__25517\,
            in1 => \N__25526\,
            in2 => \N__25505\,
            in3 => \N__31144\,
            lcout => bit_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51136\,
            ce => \N__48548\,
            sr => \N__31193\
        );

    \CLOCK_DDS.bit_cnt_i2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__31142\,
            in1 => \N__25500\,
            in2 => \_gnd_net_\,
            in3 => \N__25516\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51136\,
            ce => \N__48548\,
            sr => \N__31193\
        );

    \CLOCK_DDS.bit_cnt_i1_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25499\,
            in2 => \_gnd_net_\,
            in3 => \N__31143\,
            lcout => bit_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51136\,
            ce => \N__48548\,
            sr => \N__31193\
        );

    \comm_cmd_1__bdd_4_lut_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__31772\,
            in1 => \N__45218\,
            in2 => \N__28004\,
            in3 => \N__47140\,
            lcout => OPEN,
            ltout => \n16524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16524_bdd_4_lut_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47141\,
            in1 => \N__29183\,
            in2 => \N__25469\,
            in3 => \N__29405\,
            lcout => OPEN,
            ltout => \n16527_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_78_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__33989\,
            in1 => \N__45645\,
            in2 => \N__25466\,
            in3 => \N__47142\,
            lcout => OPEN,
            ltout => \n4_adj_1264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_82_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__39541\,
            in1 => \N__40239\,
            in2 => \N__26015\,
            in3 => \N__27893\,
            lcout => n8055,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i15_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__25921\,
            in1 => \N__26326\,
            in2 => \N__25995\,
            in3 => \N__27398\,
            lcout => buf_adcdata4_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i16_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__27393\,
            in1 => \N__26309\,
            in2 => \N__47359\,
            in3 => \N__25923\,
            lcout => buf_adcdata4_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.ADC_DATA_i17_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25922\,
            in1 => \N__25779\,
            in2 => \N__26294\,
            in3 => \N__27399\,
            lcout => buf_adcdata4_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i109_3_lut_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25668\,
            in1 => \N__28027\,
            in2 => \_gnd_net_\,
            in3 => \N__47238\,
            lcout => n71,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i26_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__26289\,
            in1 => \N__27394\,
            in2 => \N__25740\,
            in3 => \N__26849\,
            lcout => cmd_rdadctmp_26_adj_1123,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i19_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44367\,
            in1 => \N__49233\,
            in2 => \N__25715\,
            in3 => \N__26212\,
            lcout => buf_adcdata3_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i23_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49232\,
            in1 => \N__44368\,
            in2 => \N__29396\,
            in3 => \N__25669\,
            lcout => buf_adcdata3_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i28_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__25647\,
            in1 => \N__25605\,
            in2 => \N__27465\,
            in3 => \N__26848\,
            lcout => cmd_rdadctmp_28_adj_1121,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i24_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__26810\,
            in1 => \N__26325\,
            in2 => \N__27469\,
            in3 => \N__26307\,
            lcout => cmd_rdadctmp_24_adj_1125,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51160\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i23_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__26393\,
            in1 => \N__27410\,
            in2 => \N__26327\,
            in3 => \N__26811\,
            lcout => cmd_rdadctmp_23_adj_1126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51160\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3181_3_lut_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31617\,
            in1 => \N__29904\,
            in2 => \_gnd_net_\,
            in3 => \N__40528\,
            lcout => n8_adj_1227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_279_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__32812\,
            in1 => \N__28226\,
            in2 => \N__32912\,
            in3 => \N__28523\,
            lcout => n8_adj_1212,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i25_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__26308\,
            in1 => \N__27411\,
            in2 => \N__26293\,
            in3 => \N__26812\,
            lcout => cmd_rdadctmp_25_adj_1124,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51160\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_2__359_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__39640\,
            in1 => \N__34408\,
            in2 => \N__26253\,
            in3 => \N__41167\,
            lcout => \M_POW\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51160\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i131_3_lut_adj_102_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26211\,
            in1 => \N__34787\,
            in2 => \_gnd_net_\,
            in3 => \N__47245\,
            lcout => n87,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.cmd_rdadctmp_i21_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__44583\,
            in1 => \N__52793\,
            in2 => \N__46285\,
            in3 => \N__26181\,
            lcout => cmd_rdadctmp_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i6_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__33962\,
            in1 => \N__34617\,
            in2 => \N__41526\,
            in3 => \N__41373\,
            lcout => buf_dds_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_1__360_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__27915\,
            in1 => \N__34591\,
            in2 => \N__39663\,
            in3 => \N__41168\,
            lcout => \M_DCSEL\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i18_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44369\,
            in1 => \N__49189\,
            in2 => \N__26492\,
            in3 => \N__26451\,
            lcout => buf_adcdata3_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12630_2_lut_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47917\,
            lcout => n15811,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i23_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__49237\,
            in1 => \N__41585\,
            in2 => \N__36793\,
            in3 => \N__48804\,
            lcout => cmd_rdadctmp_23_adj_1089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__34407\,
            in1 => \N__31869\,
            in2 => \N__51897\,
            in3 => \N__28554\,
            lcout => \M_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i9_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44331\,
            in1 => \N__49238\,
            in2 => \N__44549\,
            in3 => \N__42087\,
            lcout => buf_adcdata3_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.cmd_rdadctmp_i22_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__26416\,
            in1 => \N__27403\,
            in2 => \N__26388\,
            in3 => \N__26753\,
            lcout => cmd_rdadctmp_22_adj_1127,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i130_3_lut_adj_291_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26362\,
            in1 => \N__34888\,
            in2 => \_gnd_net_\,
            in3 => \N__47239\,
            lcout => n90,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.adc_state_i2_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000100010"
        )
    port map (
            in0 => \N__27023\,
            in1 => \N__27097\,
            in2 => \_gnd_net_\,
            in3 => \N__27230\,
            lcout => \DTRIG_N_957_adj_1150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51212\,
            ce => \N__26962\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_218_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__27096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27022\,
            lcout => n15156,
            ltout => \n15156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i1_3_lut_adj_9_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__26657\,
            in1 => \_gnd_net_\,
            in2 => \N__26861\,
            in3 => \N__27229\,
            lcout => n9694,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i18_3_lut_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27095\,
            in2 => \N__26664\,
            in3 => \N__30636\,
            lcout => \ADC_VAC4.n15278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i1_4_lut_adj_8_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__27235\,
            in1 => \N__26637\,
            in2 => \N__27114\,
            in3 => \N__30648\,
            lcout => OPEN,
            ltout => \ADC_VAC4.n15257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i1_2_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26684\,
            in3 => \N__27018\,
            lcout => \ADC_VAC4.n15258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i1_3_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101010"
        )
    port map (
            in0 => \N__27017\,
            in1 => \_gnd_net_\,
            in2 => \N__27322\,
            in3 => \N__26675\,
            lcout => \ADC_VAC4.n14930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_198_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__27104\,
            in1 => \N__27236\,
            in2 => \N__26581\,
            in3 => \N__27016\,
            lcout => OPEN,
            ltout => \n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.CS_37_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__27237\,
            in1 => \N__26636\,
            in2 => \N__26606\,
            in3 => \N__26603\,
            lcout => \M_CS4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1457_i4_4_lut_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__26564\,
            in1 => \N__47944\,
            in2 => \N__26548\,
            in3 => \N__47310\,
            lcout => n4061,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.i13062_2_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__27234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26498\,
            lcout => \ADC_VAC4.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC4.adc_state_i1_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27252\,
            in2 => \_gnd_net_\,
            in3 => \N__27113\,
            lcout => adc_state_1_adj_1116,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51245\,
            ce => \N__26963\,
            sr => \N__26948\
        );

    \CONSTANT_ONE_LUT4_LC_13_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i4_7360_7361_set_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29029\,
            in1 => \N__26939\,
            in2 => \_gnd_net_\,
            in3 => \N__26927\,
            lcout => \comm_spi.n10471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42460\,
            ce => 'H',
            sr => \N__46655\
        );

    \comm_spi.data_tx_i4_7360_7361_reset_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29030\,
            in1 => \N__26938\,
            in2 => \_gnd_net_\,
            in3 => \N__26923\,
            lcout => \comm_spi.n10472\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42462\,
            ce => 'H',
            sr => \N__26912\
        );

    \comm_spi.i13077_4_lut_3_lut_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26877\,
            in1 => \N__30835\,
            in2 => \_gnd_net_\,
            in3 => \N__46575\,
            lcout => \comm_spi.n10444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.CS_28_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__35746\,
            in1 => \N__48388\,
            in2 => \_gnd_net_\,
            in3 => \N__48537\,
            lcout => \DDS_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51110\,
            ce => \N__31166\,
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_100_2_lut_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26878\,
            lcout => \comm_spi.data_tx_7__N_813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_92_2_lut_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46574\,
            lcout => \comm_spi.data_tx_7__N_805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_101_2_lut_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__46577\,
            in1 => \N__27687\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_93_2_lut_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27688\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46578\,
            lcout => \comm_spi.data_tx_7__N_806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13112_4_lut_3_lut_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46579\,
            in1 => \N__27689\,
            in2 => \_gnd_net_\,
            in3 => \N__27657\,
            lcout => \comm_spi.n16884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i7_7337_7338_reset_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__27658\,
            in1 => \N__27787\,
            in2 => \_gnd_net_\,
            in3 => \N__28984\,
            lcout => \comm_spi.n10449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42461\,
            ce => 'H',
            sr => \N__30996\
        );

    \i1_2_lut_adj_289_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47989\,
            in2 => \_gnd_net_\,
            in3 => \N__45298\,
            lcout => OPEN,
            ltout => \n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12648_4_lut_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__27641\,
            in1 => \N__45650\,
            in2 => \N__27623\,
            in3 => \N__29513\,
            lcout => OPEN,
            ltout => \n15466_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i103_4_lut_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__45651\,
            in1 => \N__27599\,
            in2 => \N__27620\,
            in3 => \N__47085\,
            lcout => n104,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i110_4_lut_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100000001000"
        )
    port map (
            in0 => \N__45297\,
            in1 => \N__29360\,
            in2 => \N__48046\,
            in3 => \N__31460\,
            lcout => n56,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1481_i2_4_lut_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__47086\,
            in1 => \N__27586\,
            in2 => \N__48047\,
            in3 => \N__27557\,
            lcout => n4151,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12765_2_lut_3_lut_4_lut_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33116\,
            in1 => \N__38832\,
            in2 => \N__33329\,
            in3 => \N__27860\,
            lcout => OPEN,
            ltout => \n15567_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i22_4_lut_adj_232_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50321\,
            in1 => \N__33487\,
            in2 => \N__27737\,
            in3 => \N__33632\,
            lcout => n7_adj_1255,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_196_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__43450\,
            in1 => \N__39256\,
            in2 => \_gnd_net_\,
            in3 => \N__43238\,
            lcout => n5_adj_1235,
            ltout => \n5_adj_1235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12752_4_lut_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__27722\,
            in1 => \N__33117\,
            in2 => \N__27716\,
            in3 => \N__38763\,
            lcout => OPEN,
            ltout => \n15535_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i30_4_lut_adj_265_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__49880\,
            in1 => \N__43643\,
            in2 => \N__27713\,
            in3 => \N__41936\,
            lcout => OPEN,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_178_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__52380\,
            in1 => \N__31123\,
            in2 => \N__27710\,
            in3 => \N__51898\,
            lcout => n9021,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i6_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__52384\,
            in1 => \N__51899\,
            in2 => \N__30410\,
            in3 => \N__30431\,
            lcout => data_index_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_3_lut_4_lut_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011000010"
        )
    port map (
            in0 => \N__50582\,
            in1 => \N__49479\,
            in2 => \N__52454\,
            in3 => \N__49881\,
            lcout => n8561,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i2_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27695\,
            lcout => comm_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51130\,
            ce => \N__32518\,
            sr => \N__33704\
        );

    \i1704_2_lut_3_lut_4_lut_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__38831\,
            in1 => \N__43454\,
            in2 => \N__33169\,
            in3 => \N__43281\,
            lcout => n4814,
            ltout => \n4814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i3_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__33251\,
            in1 => \_gnd_net_\,
            in2 => \N__27866\,
            in3 => \N__33448\,
            lcout => comm_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51130\,
            ce => \N__32518\,
            sr => \N__33704\
        );

    \i1_2_lut_3_lut_adj_261_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33414\,
            in2 => \N__27863\,
            in3 => \N__33250\,
            lcout => n13475,
            ltout => \n13475_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12972_2_lut_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27833\,
            in3 => \N__33111\,
            lcout => OPEN,
            ltout => \n15802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i30_4_lut_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__38830\,
            in1 => \N__50202\,
            in2 => \N__27830\,
            in3 => \N__33627\,
            lcout => n10_adj_1249,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12743_2_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38829\,
            in2 => \_gnd_net_\,
            in3 => \N__31073\,
            lcout => OPEN,
            ltout => \n15657_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i33_4_lut_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__33112\,
            in1 => \N__50203\,
            in2 => \N__27812\,
            in3 => \N__33628\,
            lcout => n13_adj_1042,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_7368_7369_set_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28907\,
            in1 => \N__28934\,
            in2 => \_gnd_net_\,
            in3 => \N__29012\,
            lcout => \comm_spi.n10479\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42438\,
            ce => 'H',
            sr => \N__27770\
        );

    \i12661_2_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41863\,
            in2 => \_gnd_net_\,
            in3 => \N__32126\,
            lcout => n15576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12670_2_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47914\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31805\,
            lcout => n15691,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12678_2_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27877\,
            in2 => \_gnd_net_\,
            in3 => \N__47915\,
            lcout => n15475,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12701_2_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__47912\,
            in1 => \N__29489\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n15835,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12746_2_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33851\,
            in2 => \_gnd_net_\,
            in3 => \N__47911\,
            lcout => n15542,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12851_2_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47913\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29545\,
            lcout => n15679,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12713_2_lut_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28065\,
            in2 => \_gnd_net_\,
            in3 => \N__47916\,
            lcout => n15543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i130_3_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27955\,
            in1 => \N__34856\,
            in2 => \_gnd_net_\,
            in3 => \N__47138\,
            lcout => OPEN,
            ltout => \n90_adj_1023_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i127_4_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__47139\,
            in1 => \N__27925\,
            in2 => \N__27896\,
            in3 => \N__45639\,
            lcout => n69_adj_1113,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i123_3_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28535\,
            in1 => \N__34154\,
            in2 => \_gnd_net_\,
            in3 => \N__47137\,
            lcout => n96,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i5_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__31846\,
            in1 => \N__36994\,
            in2 => \N__51770\,
            in3 => \N__27878\,
            lcout => buf_device_acadc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i1_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28066\,
            in1 => \N__37272\,
            in2 => \_gnd_net_\,
            in3 => \N__31847\,
            lcout => \M_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i15_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37583\,
            in1 => \N__40457\,
            in2 => \_gnd_net_\,
            in3 => \N__29511\,
            lcout => req_data_cnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__52345\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50596\,
            lcout => n8062,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12984_2_lut_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47909\,
            in2 => \_gnd_net_\,
            in3 => \N__41708\,
            lcout => n15555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_49_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32877\,
            in2 => \_gnd_net_\,
            in3 => \N__38090\,
            lcout => n3,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_280_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__32809\,
            in1 => \N__32736\,
            in2 => \N__28040\,
            in3 => \N__28028\,
            lcout => OPEN,
            ltout => \n10_adj_1242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_328_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__32735\,
            in1 => \N__38092\,
            in2 => \N__28037\,
            in3 => \N__28034\,
            lcout => eis_end,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_end_328C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i3_3_lut_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31946\,
            in1 => \N__40325\,
            in2 => \_gnd_net_\,
            in3 => \N__47910\,
            lcout => n4219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_149_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32808\,
            in2 => \_gnd_net_\,
            in3 => \N__38091\,
            lcout => n15171,
            ltout => \n15171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_3_lut_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__32878\,
            in1 => \_gnd_net_\,
            in2 => \N__28016\,
            in3 => \N__32737\,
            lcout => \raw_buf1_N_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__32813\,
            in1 => \N__28508\,
            in2 => \N__32916\,
            in3 => \N__29699\,
            lcout => eis_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__28187\,
            sr => \N__32753\
        );

    \i17_4_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__41037\,
            in1 => \N__34508\,
            in2 => \N__32923\,
            in3 => \N__28225\,
            lcout => OPEN,
            ltout => \n15356_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13047_3_lut_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32810\,
            in2 => \N__28208\,
            in3 => \N__38095\,
            lcout => n8459,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12862_2_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32911\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28522\,
            lcout => OPEN,
            ltout => \n15695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i2_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__32814\,
            in1 => \N__38096\,
            in2 => \N__28205\,
            in3 => \N__28202\,
            lcout => \eis_end_N_770\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__28187\,
            sr => \N__32753\
        );

    \i12861_3_lut_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__41038\,
            in1 => \_gnd_net_\,
            in2 => \N__32924\,
            in3 => \N__29710\,
            lcout => n15696,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12776_2_lut_3_lut_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__29711\,
            in1 => \N__38094\,
            in2 => \_gnd_net_\,
            in3 => \N__41039\,
            lcout => OPEN,
            ltout => \n15700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i1_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010011111110"
        )
    port map (
            in0 => \N__32811\,
            in1 => \N__32899\,
            in2 => \N__28196\,
            in3 => \N__28193\,
            lcout => eis_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__28187\,
            sr => \N__32753\
        );

    \comm_state_3__I_0_394_Mux_4_i15_4_lut_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52430\,
            in1 => \N__28501\,
            in2 => \N__51766\,
            in3 => \N__29887\,
            lcout => \data_index_9_N_258_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_I_3_3_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__34502\,
            in1 => \N__29459\,
            in2 => \_gnd_net_\,
            in3 => \N__31742\,
            lcout => \eis_end_N_773\,
            ltout => \eis_end_N_773_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12717_3_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__38097\,
            in1 => \_gnd_net_\,
            in2 => \N__28511\,
            in3 => \N__32889\,
            lcout => n15510,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i4_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__41826\,
            in1 => \N__51668\,
            in2 => \N__31625\,
            in3 => \N__31885\,
            lcout => \acadc_skipCount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i2_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__34593\,
            in1 => \N__31862\,
            in2 => \N__51767\,
            in3 => \N__29424\,
            lcout => \M_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i1_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__41825\,
            in1 => \N__41101\,
            in2 => \N__42187\,
            in3 => \N__51675\,
            lcout => \acadc_skipCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i4_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52431\,
            in1 => \N__28502\,
            in2 => \N__51768\,
            in3 => \N__29888\,
            lcout => data_index_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51202\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_69_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__28679\,
            in1 => \N__31884\,
            in2 => \N__28655\,
            in3 => \N__42177\,
            lcout => n18_adj_1276,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i24_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__36789\,
            in1 => \N__49239\,
            in2 => \N__28483\,
            in3 => \N__48803\,
            lcout => cmd_rdadctmp_24_adj_1088,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_1_i15_4_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52434\,
            in1 => \N__28577\,
            in2 => \N__51829\,
            in3 => \N__29959\,
            lcout => \data_index_9_N_258_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1457_i6_4_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__47860\,
            in1 => \N__28628\,
            in2 => \N__47307\,
            in3 => \N__28614\,
            lcout => n4059,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3209_3_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41092\,
            in1 => \N__29978\,
            in2 => \_gnd_net_\,
            in3 => \N__40544\,
            lcout => n8_adj_1233,
            ltout => \n8_adj_1233_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i1_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__29960\,
            in1 => \N__52435\,
            in2 => \N__28571\,
            in3 => \N__51725\,
            lcout => data_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i132_4_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__34348\,
            in1 => \N__47859\,
            in2 => \N__28558\,
            in3 => \N__45294\,
            lcout => n66_adj_1166,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i0_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29755\,
            in2 => \_gnd_net_\,
            in3 => \N__28526\,
            lcout => acadc_skipcnt_0,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => n13966,
            clk => \INVacadc_skipcnt_i0_i0C_net\,
            ce => \N__32367\,
            sr => \N__30686\
        );

    \add_58_2_THRU_CRY_0_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28767\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => n13966,
            carryout => \n13966_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_58_2_THRU_CRY_1_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28771\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n13966_THRU_CRY_0_THRU_CO\,
            carryout => \n13966_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_58_2_THRU_CRY_2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28768\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n13966_THRU_CRY_1_THRU_CO\,
            carryout => \n13966_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_58_2_THRU_CRY_3_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28772\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n13966_THRU_CRY_2_THRU_CO\,
            carryout => \n13966_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_58_2_THRU_CRY_4_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28769\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n13966_THRU_CRY_3_THRU_CO\,
            carryout => \n13966_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_58_2_THRU_CRY_5_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28773\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n13966_THRU_CRY_4_THRU_CO\,
            carryout => \n13966_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_58_2_THRU_CRY_6_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28770\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n13966_THRU_CRY_5_THRU_CO\,
            carryout => \n13966_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i1_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28678\,
            in2 => \_gnd_net_\,
            in3 => \N__28664\,
            lcout => acadc_skipcnt_1,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => n13967,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32005\,
            in2 => \_gnd_net_\,
            in3 => \N__28661\,
            lcout => acadc_skipcnt_2,
            ltout => OPEN,
            carryin => n13967,
            carryout => n13968,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i3_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32324\,
            in2 => \_gnd_net_\,
            in3 => \N__28658\,
            lcout => acadc_skipcnt_3,
            ltout => OPEN,
            carryin => n13968,
            carryout => n13969,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i4_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28651\,
            in2 => \_gnd_net_\,
            in3 => \N__28637\,
            lcout => acadc_skipcnt_4,
            ltout => OPEN,
            carryin => n13969,
            carryout => n13970,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i5_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32305\,
            in2 => \_gnd_net_\,
            in3 => \N__28634\,
            lcout => acadc_skipcnt_5,
            ltout => OPEN,
            carryin => n13970,
            carryout => n13971,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29737\,
            in2 => \_gnd_net_\,
            in3 => \N__28631\,
            lcout => acadc_skipcnt_6,
            ltout => OPEN,
            carryin => n13971,
            carryout => n13972,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i7_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31960\,
            in2 => \_gnd_net_\,
            in3 => \N__28880\,
            lcout => acadc_skipcnt_7,
            ltout => OPEN,
            carryin => n13972,
            carryout => n13973,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i8_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32290\,
            in2 => \_gnd_net_\,
            in3 => \N__28877\,
            lcout => acadc_skipcnt_8,
            ltout => OPEN,
            carryin => n13973,
            carryout => n13974,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__32371\,
            sr => \N__30707\
        );

    \acadc_skipcnt_i0_i9_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31507\,
            in2 => \_gnd_net_\,
            in3 => \N__28874\,
            lcout => acadc_skipcnt_9,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => n13975,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \acadc_skipcnt_i0_i10_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30076\,
            in2 => \_gnd_net_\,
            in3 => \N__28871\,
            lcout => acadc_skipcnt_10,
            ltout => OPEN,
            carryin => n13975,
            carryout => n13976,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \acadc_skipcnt_i0_i11_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30121\,
            in2 => \_gnd_net_\,
            in3 => \N__28868\,
            lcout => acadc_skipcnt_11,
            ltout => OPEN,
            carryin => n13976,
            carryout => n13977,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \acadc_skipcnt_i0_i12_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30028\,
            in2 => \_gnd_net_\,
            in3 => \N__28865\,
            lcout => acadc_skipcnt_12,
            ltout => OPEN,
            carryin => n13977,
            carryout => n13978,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \acadc_skipcnt_i0_i13_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32230\,
            in2 => \_gnd_net_\,
            in3 => \N__28862\,
            lcout => acadc_skipcnt_13,
            ltout => OPEN,
            carryin => n13978,
            carryout => n13979,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \acadc_skipcnt_i0_i14_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30139\,
            in2 => \_gnd_net_\,
            in3 => \N__28859\,
            lcout => acadc_skipcnt_14,
            ltout => OPEN,
            carryin => n13979,
            carryout => n13980,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \acadc_skipcnt_i0_i15_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31486\,
            in2 => \_gnd_net_\,
            in3 => \N__28856\,
            lcout => acadc_skipcnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__32375\,
            sr => \N__30703\
        );

    \mux_1469_i7_4_lut_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__29087\,
            in1 => \N__48084\,
            in2 => \N__29074\,
            in3 => \N__47084\,
            lcout => n4102,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13097_4_lut_3_lut_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29028\,
            in1 => \N__30971\,
            in2 => \_gnd_net_\,
            in3 => \N__46599\,
            lcout => \comm_spi.n16902\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i5_7364_7365_reset_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46397\,
            in1 => \N__28945\,
            in2 => \_gnd_net_\,
            in3 => \N__28963\,
            lcout => \comm_spi.n10476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42404\,
            ce => 'H',
            sr => \N__32537\
        );

    \comm_spi.data_tx_i6_7368_7369_reset_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28927\,
            in1 => \N__28897\,
            in2 => \_gnd_net_\,
            in3 => \N__29005\,
            lcout => \comm_spi.n10480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42439\,
            ce => 'H',
            sr => \N__28973\
        );

    \comm_spi.data_tx_i5_7364_7365_set_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28967\,
            in1 => \N__46396\,
            in2 => \_gnd_net_\,
            in3 => \N__28949\,
            lcout => \comm_spi.n10475\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42431\,
            ce => 'H',
            sr => \N__28916\
        );

    \comm_spi.RESET_I_0_94_2_lut_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__32562\,
            in1 => \N__46582\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13107_4_lut_3_lut_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46583\,
            in1 => \N__32563\,
            in2 => \_gnd_net_\,
            in3 => \N__28896\,
            lcout => \comm_spi.n16896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_91_2_lut_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__51404\,
            in1 => \N__46581\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.iclk_N_802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12653_2_lut_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32038\,
            lcout => n15474,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12656_2_lut_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47983\,
            in2 => \_gnd_net_\,
            in3 => \N__29239\,
            lcout => n15478,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12659_2_lut_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__47984\,
            in1 => \N__31382\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n15680,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_valid_85_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__38384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38423\,
            lcout => comm_data_vld,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.data_valid_85C_net\,
            ce => 'H',
            sr => \N__46580\
        );

    \comm_spi.imiso_83_7340_7341_set_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30843\,
            in1 => \N__29152\,
            in2 => \_gnd_net_\,
            in3 => \N__29135\,
            lcout => \comm_spi.n10451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_7340_7341_setC_net\,
            ce => 'H',
            sr => \N__30768\
        );

    \i12177_3_lut_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38765\,
            in1 => \N__39995\,
            in2 => \_gnd_net_\,
            in3 => \N__34396\,
            lcout => n15387,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12180_3_lut_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36712\,
            in1 => \N__34119\,
            in2 => \_gnd_net_\,
            in3 => \N__38764\,
            lcout => n15390,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9624_2_lut_3_lut_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__34120\,
            in1 => \N__49875\,
            in2 => \_gnd_net_\,
            in3 => \N__49543\,
            lcout => n14_adj_1211,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9632_2_lut_3_lut_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__38924\,
            in1 => \N__49879\,
            in2 => \_gnd_net_\,
            in3 => \N__49545\,
            lcout => n14_adj_1205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9637_2_lut_3_lut_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__49544\,
            in1 => \_gnd_net_\,
            in2 => \N__50111\,
            in3 => \N__41096\,
            lcout => n14_adj_1198,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i10_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__35747\,
            in1 => \N__48525\,
            in2 => \N__29213\,
            in3 => \N__34352\,
            lcout => \CLOCK_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i11_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48526\,
            in1 => \N__35748\,
            in2 => \N__29285\,
            in3 => \N__41257\,
            lcout => \CLOCK_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i12_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__32039\,
            in1 => \N__29276\,
            in2 => \N__35763\,
            in3 => \N__48527\,
            lcout => \CLOCK_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i13_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48528\,
            in1 => \N__35752\,
            in2 => \N__29270\,
            in3 => \N__34067\,
            lcout => \CLOCK_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i14_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__35753\,
            in1 => \N__48529\,
            in2 => \N__29258\,
            in3 => \N__29546\,
            lcout => \CLOCK_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i15_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__31456\,
            in1 => \N__29249\,
            in2 => \N__48546\,
            in3 => \N__35754\,
            lcout => tmp_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i9_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__29243\,
            in1 => \N__29204\,
            in2 => \N__35764\,
            in3 => \N__48536\,
            lcout => \CLOCK_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i8_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__33849\,
            in1 => \N__31217\,
            in2 => \N__48547\,
            in3 => \N__35755\,
            lcout => \CLOCK_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51143\,
            ce => \N__31210\,
            sr => \_gnd_net_\
        );

    \mux_1513_i5_4_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__45293\,
            in1 => \N__47308\,
            in2 => \N__29372\,
            in3 => \N__41600\,
            lcout => OPEN,
            ltout => \n4260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i4_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39904\,
            in1 => \_gnd_net_\,
            in2 => \N__29342\,
            in3 => \N__50131\,
            lcout => comm_buf_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51154\,
            ce => \N__44698\,
            sr => \N__44645\
        );

    \i9633_2_lut_3_lut_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__49542\,
            in1 => \N__31598\,
            in2 => \N__50290\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_1196,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9630_2_lut_3_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36967\,
            in1 => \N__50127\,
            in2 => \_gnd_net_\,
            in3 => \N__49541\,
            lcout => n14_adj_1207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12192_3_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38779\,
            in1 => \N__31597\,
            in2 => \_gnd_net_\,
            in3 => \N__36968\,
            lcout => n15402,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i11_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__30106\,
            in1 => \N__51679\,
            in2 => \N__43561\,
            in3 => \N__41827\,
            lcout => \acadc_skipCount_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_28_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__34010\,
            in1 => \N__52349\,
            in2 => \N__51769\,
            in3 => \N__50609\,
            lcout => n9224,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i8_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40464\,
            in1 => \N__37273\,
            in2 => \_gnd_net_\,
            in3 => \N__31409\,
            lcout => req_data_cnt_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i130_3_lut_adj_98_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29327\,
            in1 => \N__45216\,
            in2 => \_gnd_net_\,
            in3 => \N__30105\,
            lcout => OPEN,
            ltout => \n90_adj_1154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i125_4_lut_adj_99_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__45217\,
            in1 => \N__47864\,
            in2 => \N__29303\,
            in3 => \N__37427\,
            lcout => n72,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12629_2_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__47865\,
            in1 => \N__29428\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n15479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i30_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__36878\,
            in1 => \N__49205\,
            in2 => \N__43738\,
            in3 => \N__48818\,
            lcout => cmd_rdadctmp_30_adj_1082,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i31_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__48817\,
            in1 => \N__29386\,
            in2 => \N__49241\,
            in3 => \N__43734\,
            lcout => cmd_rdadctmp_31_adj_1081,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51167\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3157_3_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__38977\,
            in1 => \N__30258\,
            in2 => \_gnd_net_\,
            in3 => \N__40505\,
            lcout => n8_adj_1221,
            ltout => \n8_adj_1221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i7_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51636\,
            in1 => \N__52350\,
            in2 => \N__29375\,
            in3 => \N__30542\,
            lcout => data_index_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_90_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__34925\,
            in1 => \N__40324\,
            in2 => \N__31337\,
            in3 => \N__34688\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i5_3_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31576\,
            in1 => \N__40784\,
            in2 => \_gnd_net_\,
            in3 => \N__47822\,
            lcout => n4205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i9_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37238\,
            in1 => \N__40455\,
            in2 => \_gnd_net_\,
            in3 => \N__29488\,
            lcout => req_data_cnt_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i8_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__38925\,
            in1 => \N__29356\,
            in2 => \N__51738\,
            in3 => \N__31849\,
            lcout => buf_device_acadc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9631_2_lut_3_lut_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49540\,
            in1 => \N__41886\,
            in2 => \_gnd_net_\,
            in3 => \N__50288\,
            lcout => n14_adj_1206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i14_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__41887\,
            in1 => \N__29544\,
            in2 => \N__41518\,
            in3 => \N__41369\,
            lcout => buf_dds_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i3_3_lut_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29522\,
            in1 => \N__45652\,
            in2 => \_gnd_net_\,
            in3 => \N__31517\,
            lcout => n4252,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_75_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__29512\,
            in2 => \N__35402\,
            in3 => \N__29484\,
            lcout => OPEN,
            ltout => \n24_adj_1216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_113_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29468\,
            in1 => \N__31895\,
            in2 => \N__29462\,
            in3 => \N__31631\,
            lcout => n30_adj_1278,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3754_2_lut_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__49539\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50287\,
            lcout => n6791,
            ltout => \n6791_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i0_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__36715\,
            in1 => \N__41785\,
            in2 => \N__29453\,
            in3 => \N__34318\,
            lcout => \acadc_skipCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2358_3_lut_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30004\,
            in1 => \N__36714\,
            in2 => \_gnd_net_\,
            in3 => \N__40532\,
            lcout => n8_adj_1178,
            ltout => \n8_adj_1178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i0_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51664\,
            in1 => \N__52426\,
            in2 => \N__29450\,
            in3 => \N__29447\,
            lcout => data_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2356_3_lut_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30003\,
            in1 => \N__31673\,
            in2 => \_gnd_net_\,
            in3 => \N__29987\,
            lcout => n7_adj_1177,
            ltout => \n7_adj_1177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_0_i15_4_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51663\,
            in1 => \N__52425\,
            in2 => \N__29873\,
            in3 => \N__29870\,
            lcout => \data_index_9_N_258_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3201_3_lut_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__39997\,
            in1 => \N__29946\,
            in2 => \_gnd_net_\,
            in3 => \N__40533\,
            lcout => n8_adj_1231,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_70_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__29759\,
            in1 => \N__34760\,
            in2 => \N__29741\,
            in3 => \N__34314\,
            lcout => OPEN,
            ltout => \n17_adj_1277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29723\,
            in1 => \N__32246\,
            in2 => \N__29714\,
            in3 => \N__30086\,
            lcout => n31,
            ltout => \n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_304_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__38093\,
            in1 => \_gnd_net_\,
            in2 => \N__29702\,
            in3 => \N__41045\,
            lcout => n15187,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i2_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52433\,
            in1 => \N__29693\,
            in2 => \N__51844\,
            in3 => \N__29927\,
            lcout => data_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_2_i15_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52432\,
            in1 => \N__29692\,
            in2 => \N__51842\,
            in3 => \N__29926\,
            lcout => \data_index_9_N_258_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i12_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__36990\,
            in1 => \N__41824\,
            in2 => \N__30058\,
            in3 => \N__51749\,
            lcout => \acadc_skipCount_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i4_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__29565\,
            in1 => \N__43558\,
            in2 => \N__51843\,
            in3 => \N__31871\,
            lcout => \M_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__41704\,
            in1 => \N__30143\,
            in2 => \N__30125\,
            in3 => \N__30107\,
            lcout => OPEN,
            ltout => \n23_adj_1199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31472\,
            in1 => \N__31919\,
            in2 => \N__30089\,
            in3 => \N__30014\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__30080\,
            in1 => \N__30048\,
            in2 => \N__30032\,
            in3 => \N__34206\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_2_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43616\,
            in2 => \N__30008\,
            in3 => \_gnd_net_\,
            lcout => \data_index_9_N_647_0\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => n14031,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_3_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__29977\,
            in1 => \N__29976\,
            in2 => \N__31699\,
            in3 => \N__29951\,
            lcout => n7_adj_1232,
            ltout => OPEN,
            carryin => n14031,
            carryout => n14032,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_4_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__29947\,
            in2 => \N__31703\,
            in3 => \N__29918\,
            lcout => n7_adj_1230,
            ltout => OPEN,
            carryin => n14032,
            carryout => n14033,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_5_lut_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__30232\,
            in1 => \N__30231\,
            in2 => \N__31700\,
            in3 => \N__29915\,
            lcout => n7_adj_1228,
            ltout => OPEN,
            carryin => n14033,
            carryout => n14034,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_6_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__29912\,
            in1 => \N__29911\,
            in2 => \N__31704\,
            in3 => \N__29876\,
            lcout => n7_adj_1226,
            ltout => OPEN,
            carryin => n14034,
            carryout => n14035,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_7_lut_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32056\,
            in1 => \N__32055\,
            in2 => \N__31701\,
            in3 => \N__30266\,
            lcout => n7_adj_1224,
            ltout => OPEN,
            carryin => n14035,
            carryout => n14036,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_8_lut_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__30577\,
            in1 => \N__30576\,
            in2 => \N__31705\,
            in3 => \N__30263\,
            lcout => n7_adj_1222,
            ltout => OPEN,
            carryin => n14036,
            carryout => n14037,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_9_lut_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__30260\,
            in1 => \N__30259\,
            in2 => \N__31702\,
            in3 => \N__30239\,
            lcout => n7_adj_1220,
            ltout => OPEN,
            carryin => n14037,
            carryout => n14038,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1443_10_lut_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32657\,
            in1 => \N__32656\,
            in2 => \N__31712\,
            in3 => \N__30236\,
            lcout => n7_adj_1218,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i19_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__38284\,
            in1 => \N__46089\,
            in2 => \N__46164\,
            in3 => \N__53474\,
            lcout => cmd_rdadctmp_19_adj_1057,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3145_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32655\,
            in1 => \N__34124\,
            in2 => \_gnd_net_\,
            in3 => \N__40545\,
            lcout => n8_adj_1219,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3193_3_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40546\,
            in1 => \N__44776\,
            in2 => \_gnd_net_\,
            in3 => \N__30233\,
            lcout => n8_adj_1229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i3_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52442\,
            in1 => \N__32501\,
            in2 => \N__51918\,
            in3 => \N__32489\,
            lcout => data_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51269\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.i18_3_lut_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30212\,
            in1 => \N__36475\,
            in2 => \_gnd_net_\,
            in3 => \N__30604\,
            lcout => \ADC_VAC2.n15280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13029_2_lut_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32345\,
            lcout => n10532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13050_2_lut_3_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32729\,
            in1 => \N__32836\,
            in2 => \_gnd_net_\,
            in3 => \N__38122\,
            lcout => n15344,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17_3_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__38123\,
            in1 => \N__32925\,
            in2 => \N__32840\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n15328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_trig_329_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__32728\,
            in1 => \N__30674\,
            in2 => \N__30662\,
            in3 => \N__30618\,
            lcout => acadc_trig,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_329C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3165_3_lut_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33969\,
            in1 => \N__30578\,
            in2 => \_gnd_net_\,
            in3 => \N__40547\,
            lcout => n8_adj_1223,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_7_i15_4_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52467\,
            in1 => \N__30551\,
            in2 => \N__51909\,
            in3 => \N__30541\,
            lcout => \data_index_9_N_258_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_6_i15_4_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__52468\,
            in1 => \N__30424\,
            in2 => \N__30397\,
            in3 => \N__51851\,
            lcout => \data_index_9_N_258_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i7336_3_lut_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30788\,
            in1 => \N__30272\,
            in2 => \_gnd_net_\,
            in3 => \N__30844\,
            lcout => \ICE_SPI_MISO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.MISO_48_7334_7335_reset_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30890\,
            in1 => \N__30863\,
            in2 => \_gnd_net_\,
            in3 => \N__30834\,
            lcout => \comm_spi.n10446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_7334_7335_resetC_net\,
            ce => 'H',
            sr => \N__31000\
        );

    \comm_spi.RESET_I_0_104_2_lut_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30967\,
            lcout => \comm_spi.data_tx_7__N_825\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i105_4_lut_adj_131_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010001000"
        )
    port map (
            in0 => \N__45285\,
            in1 => \N__30917\,
            in2 => \N__37610\,
            in3 => \N__47855\,
            lcout => n66,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.MISO_48_7334_7335_set_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30886\,
            in1 => \N__30856\,
            in2 => \_gnd_net_\,
            in3 => \N__30842\,
            lcout => \comm_spi.n10445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_7334_7335_setC_net\,
            ce => 'H',
            sr => \N__30778\
        );

    \i1_2_lut_3_lut_adj_176_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__52238\,
            in1 => \N__49996\,
            in2 => \_gnd_net_\,
            in3 => \N__49504\,
            lcout => n15204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_181_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__49505\,
            in1 => \_gnd_net_\,
            in2 => \N__50219\,
            in3 => \N__52239\,
            lcout => n10640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_216_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__52240\,
            in1 => \N__50000\,
            in2 => \_gnd_net_\,
            in3 => \N__49507\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9642_2_lut_3_lut_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__37883\,
            in1 => \N__50004\,
            in2 => \_gnd_net_\,
            in3 => \N__49508\,
            lcout => n14_adj_1213,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9697_2_lut_3_lut_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__49506\,
            in1 => \_gnd_net_\,
            in2 => \N__50220\,
            in3 => \N__38976\,
            lcout => n14_adj_1168,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_262_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49471\,
            in2 => \_gnd_net_\,
            in3 => \N__50580\,
            lcout => n15176,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12186_3_lut_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__38766\,
            in1 => \N__44774\,
            in2 => \_gnd_net_\,
            in3 => \N__43560\,
            lcout => n15396,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12817_4_lut_4_lut_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000010000"
        )
    port map (
            in0 => \N__49868\,
            in1 => \N__49470\,
            in2 => \N__43439\,
            in3 => \N__43255\,
            lcout => n15527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__49473\,
            in1 => \N__52360\,
            in2 => \_gnd_net_\,
            in3 => \N__49870\,
            lcout => n8133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i34_4_lut_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__49874\,
            in1 => \N__33625\,
            in2 => \N__31094\,
            in3 => \N__31082\,
            lcout => n15_adj_1203,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_3_lut_4_lut_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000111100000"
        )
    port map (
            in0 => \N__49869\,
            in1 => \N__49472\,
            in2 => \N__52446\,
            in3 => \N__50581\,
            lcout => n10566,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i0_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__48518\,
            in1 => \N__35734\,
            in2 => \N__33875\,
            in3 => \N__31036\,
            lcout => \CLOCK_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i1_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__35735\,
            in1 => \N__48519\,
            in2 => \N__31025\,
            in3 => \N__42125\,
            lcout => \CLOCK_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i2_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48520\,
            in1 => \N__35736\,
            in2 => \N__31016\,
            in3 => \N__43685\,
            lcout => \CLOCK_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.i1_4_lut_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100110"
        )
    port map (
            in0 => \N__35733\,
            in1 => \N__48387\,
            in2 => \N__33908\,
            in3 => \N__48517\,
            lcout => \CLOCK_DDS.n9759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i3_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48521\,
            in1 => \N__35737\,
            in2 => \N__31262\,
            in3 => \N__40969\,
            lcout => \CLOCK_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i4_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__31577\,
            in1 => \N__31253\,
            in2 => \N__35759\,
            in3 => \N__48522\,
            lcout => \CLOCK_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i5_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48523\,
            in1 => \N__35741\,
            in2 => \N__31244\,
            in3 => \N__34233\,
            lcout => \CLOCK_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i6_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__35742\,
            in1 => \N__48524\,
            in2 => \N__31235\,
            in3 => \N__34628\,
            lcout => \CLOCK_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51155\,
            ce => \N__31209\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.tmp_buf_i7_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__48506\,
            in1 => \N__35732\,
            in2 => \N__31226\,
            in3 => \N__31730\,
            lcout => \CLOCK_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51168\,
            ce => \N__31211\,
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.i7713_3_lut_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__35728\,
            in1 => \N__48383\,
            in2 => \_gnd_net_\,
            in3 => \N__48503\,
            lcout => n10823,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.i23_4_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000010101"
        )
    port map (
            in0 => \N__48505\,
            in1 => \N__33896\,
            in2 => \N__48389\,
            in3 => \N__35731\,
            lcout => \CLOCK_DDS.n9_adj_1021\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.i13064_4_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__35730\,
            in1 => \N__48382\,
            in2 => \N__33903\,
            in3 => \N__48504\,
            lcout => \CLOCK_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12766_2_lut_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31151\,
            in2 => \_gnd_net_\,
            in3 => \N__35729\,
            lcout => n15640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i8_3_lut_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31729\,
            in1 => \N__36763\,
            in2 => \_gnd_net_\,
            in3 => \N__47702\,
            lcout => n4202,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i8_3_lut_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31316\,
            in1 => \_gnd_net_\,
            in2 => \N__45653\,
            in3 => \N__33806\,
            lcout => n4247,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i7_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37318\,
            in1 => \N__40434\,
            in2 => \_gnd_net_\,
            in3 => \N__31336\,
            lcout => req_data_cnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i7_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__41818\,
            in1 => \N__51915\,
            in2 => \N__38971\,
            in3 => \N__31986\,
            lcout => \acadc_skipCount_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12655_2_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47810\,
            in2 => \_gnd_net_\,
            in3 => \N__31911\,
            lcout => n15556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i14_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31912\,
            in1 => \_gnd_net_\,
            in2 => \N__40460\,
            in3 => \N__37630\,
            lcout => req_data_cnt_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51186\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i111_4_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__36843\,
            in1 => \N__45598\,
            in2 => \N__31553\,
            in3 => \N__47150\,
            lcout => n60_adj_1157,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i3_4_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__47151\,
            in1 => \N__45306\,
            in2 => \N__43661\,
            in3 => \N__31280\,
            lcout => n4262,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_299_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101111"
        )
    port map (
            in0 => \N__50561\,
            in1 => \_gnd_net_\,
            in2 => \N__49538\,
            in3 => \N__49966\,
            lcout => n7567,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i8_4_lut_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000010000"
        )
    port map (
            in0 => \N__47152\,
            in1 => \N__45307\,
            in2 => \N__31271\,
            in3 => \N__31466\,
            lcout => n4257,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__34889\,
            in1 => \N__31422\,
            in2 => \N__35453\,
            in3 => \N__31407\,
            lcout => n19_adj_1234,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i15_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__31452\,
            in1 => \N__38926\,
            in2 => \N__41511\,
            in3 => \N__41356\,
            lcout => buf_dds_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i13_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37663\,
            in1 => \N__40454\,
            in2 => \_gnd_net_\,
            in3 => \N__31423\,
            lcout => req_data_cnt_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12710_2_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__31408\,
            in1 => \_gnd_net_\,
            in2 => \N__47918\,
            in3 => \_gnd_net_\,
            lcout => n15812,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i7_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__41896\,
            in1 => \N__31848\,
            in2 => \N__51739\,
            in3 => \N__31378\,
            lcout => buf_device_acadc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_292_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010001000"
        )
    port map (
            in0 => \N__47816\,
            in1 => \N__40982\,
            in2 => \N__31364\,
            in3 => \N__41935\,
            lcout => n99,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i8_3_lut_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47815\,
            in1 => \N__31335\,
            in2 => \_gnd_net_\,
            in3 => \N__31991\,
            lcout => n4214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i4_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40471\,
            in1 => \N__37400\,
            in2 => \_gnd_net_\,
            in3 => \N__34658\,
            lcout => req_data_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i10_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37190\,
            in1 => \N__40472\,
            in2 => \_gnd_net_\,
            in3 => \N__34177\,
            lcout => req_data_cnt_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i7_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38972\,
            in1 => \N__31728\,
            in2 => \N__41506\,
            in3 => \N__41361\,
            lcout => buf_dds_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_288_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110111011"
        )
    port map (
            in0 => \N__52443\,
            in1 => \N__31674\,
            in2 => \N__51737\,
            in3 => \N__40543\,
            lcout => n9187,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_94_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__34030\,
            in1 => \N__34820\,
            in2 => \N__35477\,
            in3 => \N__34176\,
            lcout => n21_adj_1204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i4_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__31624\,
            in1 => \N__31575\,
            in2 => \N__41505\,
            in3 => \N__41360\,
            lcout => buf_dds_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_5__356_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__39662\,
            in1 => \N__31549\,
            in2 => \N__33794\,
            in3 => \N__41151\,
            lcout => buf_control_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51221\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1494_i3_3_lut_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47805\,
            in1 => \N__37039\,
            in2 => \_gnd_net_\,
            in3 => \N__34684\,
            lcout => OPEN,
            ltout => \n4195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i3_4_lut_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__31535\,
            in1 => \N__47806\,
            in2 => \N__31520\,
            in3 => \N__45239\,
            lcout => n4232,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__31511\,
            in1 => \N__41656\,
            in2 => \N__31493\,
            in3 => \N__31782\,
            lcout => n24_adj_1174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i9_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__31784\,
            in1 => \N__34594\,
            in2 => \N__41828\,
            in3 => \N__51853\,
            lcout => \acadc_skipCount_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51238\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_92_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__34786\,
            in1 => \N__31913\,
            in2 => \N__35429\,
            in3 => \N__37423\,
            lcout => n23_adj_1194,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i5_3_lut_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47811\,
            in1 => \N__34653\,
            in2 => \_gnd_net_\,
            in3 => \N__31889\,
            lcout => n4217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__51852\,
            in1 => \N__33789\,
            in2 => \N__31870\,
            in3 => \N__31798\,
            lcout => buf_device_acadc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51238\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13004_2_lut_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47804\,
            lcout => n15834,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i8_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__41789\,
            in1 => \N__51880\,
            in2 => \N__34141\,
            in3 => \N__32271\,
            lcout => \acadc_skipCount_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i2_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51879\,
            in1 => \N__41790\,
            in2 => \N__31945\,
            in3 => \N__39996\,
            lcout => \acadc_skipCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3173_3_lut_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32057\,
            in1 => \N__37870\,
            in2 => \_gnd_net_\,
            in3 => \N__40534\,
            lcout => n8_adj_1225,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_103_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38166\,
            in1 => \N__38332\,
            in2 => \N__37771\,
            in3 => \N__42015\,
            lcout => OPEN,
            ltout => \n20_adj_1253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34634\,
            in1 => \N__31760\,
            in2 => \N__31745\,
            in3 => \N__34298\,
            lcout => n29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12715_2_lut_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34134\,
            in2 => \_gnd_net_\,
            in3 => \N__32125\,
            lcout => n15546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i23_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__53605\,
            in1 => \N__46082\,
            in2 => \N__34470\,
            in3 => \N__53481\,
            lcout => cmd_rdadctmp_23_adj_1053,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i5_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__51508\,
            in1 => \N__51869\,
            in2 => \N__52489\,
            in3 => \N__52184\,
            lcout => data_index_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i6_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41820\,
            in1 => \N__33961\,
            in2 => \N__51917\,
            in3 => \N__34759\,
            lcout => \acadc_skipCount_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i12_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__36995\,
            in1 => \N__41510\,
            in2 => \N__32031\,
            in3 => \N__41374\,
            lcout => buf_dds_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32009\,
            in1 => \N__31987\,
            in2 => \N__31967\,
            in3 => \N__31935\,
            lcout => n22_adj_1170,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i3_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51867\,
            in1 => \N__40470\,
            in2 => \N__44775\,
            in3 => \N__38170\,
            lcout => req_data_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i10_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41819\,
            in1 => \N__34424\,
            in2 => \N__51916\,
            in3 => \N__34210\,
            lcout => \acadc_skipCount_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i13_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51866\,
            in1 => \N__41821\,
            in2 => \N__32215\,
            in3 => \N__33793\,
            lcout => \acadc_skipCount_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51270\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_3_i15_4_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52466\,
            in1 => \N__32500\,
            in2 => \N__51913\,
            in3 => \N__32488\,
            lcout => \data_index_9_N_258_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13054_3_lut_4_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__32833\,
            in1 => \N__32926\,
            in2 => \N__32767\,
            in3 => \N__38127\,
            lcout => n8456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i3_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51868\,
            in1 => \N__41822\,
            in2 => \N__44777\,
            in3 => \N__38146\,
            lcout => \acadc_skipCount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i5_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__37741\,
            in1 => \N__37882\,
            in2 => \N__51914\,
            in3 => \N__41823\,
            lcout => \acadc_skipCount_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51282\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__32323\,
            in1 => \N__37740\,
            in2 => \N__32309\,
            in3 => \N__38145\,
            lcout => OPEN,
            ltout => \n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__32291\,
            in1 => \N__32272\,
            in2 => \N__32249\,
            in3 => \N__32189\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_46_i14_2_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32234\,
            in2 => \_gnd_net_\,
            in3 => \N__32205\,
            lcout => n14_adj_1160,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i8_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53101\,
            in1 => \N__32140\,
            in2 => \N__32183\,
            in3 => \N__52897\,
            lcout => buf_adcdata1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__32930\,
            in1 => \N__32834\,
            in2 => \N__32763\,
            in3 => \N__38132\,
            lcout => n9790,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i8_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__52469\,
            in1 => \N__42580\,
            in2 => \N__51931\,
            in3 => \N__42601\,
            lcout => data_index_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.dds_state_i2_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35669\,
            in2 => \_gnd_net_\,
            in3 => \N__48420\,
            lcout => dds_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1481_i4_4_lut_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__48048\,
            in2 => \N__47309\,
            in3 => \N__32623\,
            lcout => n4149,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_102_2_lut_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32564\,
            in2 => \_gnd_net_\,
            in3 => \N__46561\,
            lcout => \comm_spi.data_tx_7__N_819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i1_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100100000"
        )
    port map (
            in0 => \N__43298\,
            in1 => \N__43441\,
            in2 => \N__38693\,
            in3 => \N__33020\,
            lcout => comm_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51132\,
            ce => \N__32522\,
            sr => \N__33693\
        );

    \comm_index_i0_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__43440\,
            in1 => \N__38642\,
            in2 => \_gnd_net_\,
            in3 => \N__43297\,
            lcout => comm_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51132\,
            ce => \N__32522\,
            sr => \N__33693\
        );

    \i12636_3_lut_4_lut_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__40237\,
            in1 => \N__45302\,
            in2 => \N__33559\,
            in3 => \N__47236\,
            lcout => n15463,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12637_3_lut_4_lut_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__47237\,
            in1 => \N__33371\,
            in2 => \N__45313\,
            in3 => \N__40238\,
            lcout => OPEN,
            ltout => \n15460_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i39_4_lut_adj_64_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__33649\,
            in1 => \N__33372\,
            in2 => \N__33596\,
            in3 => \N__45604\,
            lcout => OPEN,
            ltout => \n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i3_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__33373\,
            in1 => \N__47852\,
            in2 => \N__33593\,
            in3 => \N__36586\,
            lcout => comm_length_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51144\,
            ce => \N__50660\,
            sr => \N__33700\
        );

    \i39_4_lut_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__33555\,
            in1 => \N__33590\,
            in2 => \N__33650\,
            in3 => \N__45603\,
            lcout => OPEN,
            ltout => \n19_adj_1151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i2_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111111011"
        )
    port map (
            in0 => \N__33584\,
            in1 => \N__38996\,
            in2 => \N__33569\,
            in3 => \N__47853\,
            lcout => comm_length_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51144\,
            ce => \N__50660\,
            sr => \N__33700\
        );

    \i2_4_lut_adj_281_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__33551\,
            in1 => \N__33486\,
            in2 => \N__33374\,
            in3 => \N__33320\,
            lcout => OPEN,
            ltout => \n6_adj_1281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_283_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111110"
        )
    port map (
            in0 => \N__33715\,
            in1 => \N__32948\,
            in2 => \N__33215\,
            in3 => \N__38630\,
            lcout => n7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_200_i2_2_lut_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32938\,
            in2 => \_gnd_net_\,
            in3 => \N__33085\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_55_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__32939\,
            in1 => \N__40910\,
            in2 => \N__39475\,
            in3 => \N__41221\,
            lcout => OPEN,
            ltout => \n15119_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i1_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__36605\,
            in1 => \N__40925\,
            in2 => \N__32942\,
            in3 => \N__33728\,
            lcout => comm_length_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51156\,
            ce => \N__50656\,
            sr => \N__33692\
        );

    \i1_2_lut_3_lut_4_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101010"
        )
    port map (
            in0 => \N__40880\,
            in1 => \N__44969\,
            in2 => \N__47232\,
            in3 => \N__43198\,
            lcout => n5_adj_1282,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_209_i13_2_lut_3_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__43197\,
            in1 => \N__47095\,
            in2 => \_gnd_net_\,
            in3 => \N__40879\,
            lcout => n13,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_54_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33731\,
            in3 => \N__38995\,
            lcout => n6_adj_1273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i0_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110111111111"
        )
    port map (
            in0 => \N__33722\,
            in1 => \N__33716\,
            in2 => \N__39476\,
            in3 => \N__41166\,
            lcout => comm_length_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51156\,
            ce => \N__50656\,
            sr => \N__33692\
        );

    \i1_4_lut_adj_209_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010000"
        )
    port map (
            in0 => \N__50536\,
            in1 => \N__33656\,
            in2 => \N__52447\,
            in3 => \N__51841\,
            lcout => n8253,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9554_2_lut_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__47047\,
            in1 => \N__45229\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n12649,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_250_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__52217\,
            in1 => \N__49531\,
            in2 => \N__42755\,
            in3 => \N__36595\,
            lcout => n8525,
            ltout => \n8525_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i5_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__37369\,
            in1 => \N__34234\,
            in2 => \N__33635\,
            in3 => \N__52218\,
            lcout => buf_dds_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_230_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__40212\,
            in1 => \N__39590\,
            in2 => \N__36566\,
            in3 => \N__47046\,
            lcout => n4075,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds_333_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__36596\,
            in1 => \N__33914\,
            in2 => \N__33907\,
            in3 => \N__41498\,
            lcout => trig_dds,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i0_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__36716\,
            in1 => \N__33870\,
            in2 => \N__41520\,
            in3 => \N__41313\,
            lcout => buf_dds_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i8_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__41312\,
            in1 => \N__34133\,
            in2 => \N__33850\,
            in3 => \N__41497\,
            lcout => buf_dds_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1494_i8_3_lut_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37298\,
            in1 => \N__47700\,
            in2 => \_gnd_net_\,
            in3 => \N__34921\,
            lcout => OPEN,
            ltout => \n4190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i8_4_lut_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__47701\,
            in1 => \N__33821\,
            in2 => \N__33809\,
            in3 => \N__45240\,
            lcout => n4227,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i2_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40116\,
            in1 => \N__50123\,
            in2 => \_gnd_net_\,
            in3 => \N__33800\,
            lcout => comm_buf_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51187\,
            ce => \N__44711\,
            sr => \N__44653\
        );

    \i9634_2_lut_3_lut_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49546\,
            in1 => \N__39970\,
            in2 => \_gnd_net_\,
            in3 => \N__50120\,
            lcout => n14_adj_1197,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9627_2_lut_3_lut_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__50121\,
            in1 => \N__34592\,
            in2 => \_gnd_net_\,
            in3 => \N__49547\,
            lcout => n14_adj_1210,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9628_2_lut_3_lut_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49548\,
            in1 => \N__34409\,
            in2 => \_gnd_net_\,
            in3 => \N__50122\,
            lcout => n14_adj_1209,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9638_2_lut_3_lut_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__49819\,
            in1 => \N__33775\,
            in2 => \_gnd_net_\,
            in3 => \N__49549\,
            lcout => n14_adj_1202,
            ltout => \n14_adj_1202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i13_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__52300\,
            in1 => \N__34060\,
            in2 => \N__34070\,
            in3 => \N__41346\,
            lcout => buf_dds_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12856_2_lut_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47824\,
            lcout => n15690,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i12_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40433\,
            in1 => \N__37718\,
            in2 => \_gnd_net_\,
            in3 => \N__34029\,
            lcout => req_data_cnt_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_206_i13_2_lut_3_lut_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__43199\,
            in1 => \N__47027\,
            in2 => \_gnd_net_\,
            in3 => \N__40875\,
            lcout => n13_adj_1026,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_71_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__34507\,
            in1 => \N__45597\,
            in2 => \N__37214\,
            in3 => \N__45264\,
            lcout => OPEN,
            ltout => \n78_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_77_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011000000"
        )
    port map (
            in0 => \N__34001\,
            in1 => \N__47823\,
            in2 => \N__33992\,
            in3 => \N__41931\,
            lcout => n99_adj_1024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i7_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39361\,
            in1 => \N__50152\,
            in2 => \_gnd_net_\,
            in3 => \N__33977\,
            lcout => comm_buf_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51222\,
            ce => \N__44712\,
            sr => \N__44641\
        );

    \comm_buf_1__i0_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50149\,
            in1 => \N__39187\,
            in2 => \_gnd_net_\,
            in3 => \N__37088\,
            lcout => comm_buf_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51222\,
            ce => \N__44712\,
            sr => \N__44641\
        );

    \comm_buf_1__i6_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40715\,
            in1 => \N__50151\,
            in2 => \_gnd_net_\,
            in3 => \N__34703\,
            lcout => comm_buf_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51222\,
            ce => \N__44712\,
            sr => \N__44641\
        );

    \comm_buf_1__i1_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50150\,
            in1 => \N__44158\,
            in2 => \_gnd_net_\,
            in3 => \N__42137\,
            lcout => comm_buf_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51222\,
            ce => \N__44712\,
            sr => \N__44641\
        );

    \i105_4_lut_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__45233\,
            in1 => \N__37649\,
            in2 => \N__34268\,
            in3 => \N__47744\,
            lcout => n66_adj_1158,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i6_3_lut_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47745\,
            in1 => \_gnd_net_\,
            in2 => \N__34238\,
            in3 => \N__37512\,
            lcout => n4204,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_228_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__45231\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47742\,
            lcout => n93,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i130_3_lut_adj_85_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34186\,
            in1 => \N__45230\,
            in2 => \_gnd_net_\,
            in3 => \N__34214\,
            lcout => n90_adj_1167,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_adj_215_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__44963\,
            in1 => \N__47174\,
            in2 => \N__39664\,
            in3 => \N__40885\,
            lcout => n7485,
            ltout => \n7485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tacadc_rst_364_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34187\,
            in1 => \_gnd_net_\,
            in2 => \N__34190\,
            in3 => \N__34419\,
            lcout => tacadc_rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i125_4_lut_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__45232\,
            in1 => \N__34178\,
            in2 => \N__34163\,
            in3 => \N__47743\,
            lcout => n72_adj_1162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_start_366_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34142\,
            in1 => \N__34519\,
            in2 => \_gnd_net_\,
            in3 => \N__41044\,
            lcout => eis_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51239\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_109_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__42159\,
            in1 => \N__37811\,
            in2 => \N__34657\,
            in3 => \N__38228\,
            lcout => n18_adj_1217,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i7_3_lut_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47920\,
            in1 => \_gnd_net_\,
            in2 => \N__34624\,
            in3 => \N__41557\,
            lcout => n4203,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_stop_365_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34595\,
            in1 => \N__34523\,
            in2 => \_gnd_net_\,
            in3 => \N__34506\,
            lcout => eis_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i15_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53809\,
            in1 => \N__34441\,
            in2 => \N__34474\,
            in3 => \N__53433\,
            lcout => buf_adcdata2_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i10_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__34423\,
            in1 => \N__41525\,
            in2 => \N__41381\,
            in3 => \N__34341\,
            lcout => buf_dds_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i1_3_lut_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47919\,
            in1 => \N__34322\,
            in2 => \_gnd_net_\,
            in3 => \N__34285\,
            lcout => n4221,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_112_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__34945\,
            in1 => \N__36648\,
            in2 => \N__37922\,
            in3 => \N__34284\,
            lcout => n17_adj_1214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i5_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__40458\,
            in1 => \N__37874\,
            in2 => \N__37772\,
            in3 => \N__51895\,
            lcout => req_data_cnt_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i0_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51894\,
            in1 => \N__40459\,
            in2 => \N__34292\,
            in3 => \N__36713\,
            lcout => req_data_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51271\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i7_3_lut_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47922\,
            in1 => \N__34758\,
            in2 => \_gnd_net_\,
            in3 => \N__37921\,
            lcout => n4215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1494_i7_3_lut_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37346\,
            in1 => \N__47923\,
            in2 => \_gnd_net_\,
            in3 => \N__34944\,
            lcout => OPEN,
            ltout => \n4191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i7_4_lut_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__47924\,
            in1 => \N__34739\,
            in2 => \N__34724\,
            in3 => \N__45295\,
            lcout => OPEN,
            ltout => \n4228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i7_3_lut_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34721\,
            in2 => \N__34715\,
            in3 => \N__45649\,
            lcout => OPEN,
            ltout => \n4248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i7_4_lut_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__34712\,
            in1 => \N__47173\,
            in2 => \N__34706\,
            in3 => \N__45296\,
            lcout => n4258,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_cntvec_i0_i0_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36649\,
            in2 => \_gnd_net_\,
            in3 => \N__34694\,
            lcout => data_cntvec_0,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => n13951,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i1_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38227\,
            in2 => \_gnd_net_\,
            in3 => \N__34691\,
            lcout => data_cntvec_1,
            ltout => OPEN,
            carryin => n13951,
            carryout => n13952,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i2_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34683\,
            in2 => \_gnd_net_\,
            in3 => \N__34661\,
            lcout => data_cntvec_2,
            ltout => OPEN,
            carryin => n13952,
            carryout => n13953,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i3_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42016\,
            in2 => \_gnd_net_\,
            in3 => \N__34955\,
            lcout => data_cntvec_3,
            ltout => OPEN,
            carryin => n13953,
            carryout => n13954,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i4_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37810\,
            in2 => \_gnd_net_\,
            in3 => \N__34952\,
            lcout => data_cntvec_4,
            ltout => OPEN,
            carryin => n13954,
            carryout => n13955,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38333\,
            in2 => \_gnd_net_\,
            in3 => \N__34949\,
            lcout => data_cntvec_5,
            ltout => OPEN,
            carryin => n13955,
            carryout => n13956,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i6_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34946\,
            in2 => \_gnd_net_\,
            in3 => \N__34928\,
            lcout => data_cntvec_6,
            ltout => OPEN,
            carryin => n13956,
            carryout => n13957,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i7_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34920\,
            in2 => \_gnd_net_\,
            in3 => \N__34892\,
            lcout => data_cntvec_7,
            ltout => OPEN,
            carryin => n13957,
            carryout => n13958,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__38048\,
            sr => \N__38006\
        );

    \data_cntvec_i0_i8_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34881\,
            in2 => \_gnd_net_\,
            in3 => \N__34859\,
            lcout => data_cntvec_8,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => n13959,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i9_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34845\,
            in2 => \_gnd_net_\,
            in3 => \N__34823\,
            lcout => data_cntvec_9,
            ltout => OPEN,
            carryin => n13959,
            carryout => n13960,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i10_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34812\,
            in2 => \_gnd_net_\,
            in3 => \N__34790\,
            lcout => data_cntvec_10,
            ltout => OPEN,
            carryin => n13960,
            carryout => n13961,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i11_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34782\,
            in2 => \_gnd_net_\,
            in3 => \N__34763\,
            lcout => data_cntvec_11,
            ltout => OPEN,
            carryin => n13961,
            carryout => n13962,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i12_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35470\,
            in2 => \_gnd_net_\,
            in3 => \N__35456\,
            lcout => data_cntvec_12,
            ltout => OPEN,
            carryin => n13962,
            carryout => n13963,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i13_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35446\,
            in2 => \_gnd_net_\,
            in3 => \N__35432\,
            lcout => data_cntvec_13,
            ltout => OPEN,
            carryin => n13963,
            carryout => n13964,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i14_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35422\,
            in2 => \_gnd_net_\,
            in3 => \N__35408\,
            lcout => data_cntvec_14,
            ltout => OPEN,
            carryin => n13964,
            carryout => n13965,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_cntvec_i0_i15_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35395\,
            in2 => \_gnd_net_\,
            in3 => \N__35405\,
            lcout => data_cntvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__38042\,
            sr => \N__38005\
        );

    \data_count_i0_i0_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35298\,
            in2 => \_gnd_net_\,
            in3 => \N__35276\,
            lcout => data_count_0,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => n13942,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35193\,
            in2 => \_gnd_net_\,
            in3 => \N__35171\,
            lcout => data_count_1,
            ltout => OPEN,
            carryin => n13942,
            carryout => n13943,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i2_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35088\,
            in2 => \_gnd_net_\,
            in3 => \N__35066\,
            lcout => data_count_2,
            ltout => OPEN,
            carryin => n13943,
            carryout => n13944,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i3_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34980\,
            in2 => \_gnd_net_\,
            in3 => \N__34958\,
            lcout => data_count_3,
            ltout => OPEN,
            carryin => n13944,
            carryout => n13945,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i4_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36216\,
            in2 => \_gnd_net_\,
            in3 => \N__36194\,
            lcout => data_count_4,
            ltout => OPEN,
            carryin => n13945,
            carryout => n13946,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i5_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36108\,
            in2 => \_gnd_net_\,
            in3 => \N__36086\,
            lcout => data_count_5,
            ltout => OPEN,
            carryin => n13946,
            carryout => n13947,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i6_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36000\,
            in2 => \_gnd_net_\,
            in3 => \N__35978\,
            lcout => data_count_6,
            ltout => OPEN,
            carryin => n13947,
            carryout => n13948,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i7_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35895\,
            in2 => \_gnd_net_\,
            in3 => \N__35873\,
            lcout => data_count_7,
            ltout => OPEN,
            carryin => n13948,
            carryout => n13949,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__38041\,
            sr => \N__37995\
        );

    \data_count_i0_i8_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35787\,
            in2 => \_gnd_net_\,
            in3 => \N__35870\,
            lcout => data_count_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__38043\,
            sr => \N__37994\
        );

    \CLOCK_DDS.dds_state_i1_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35670\,
            in2 => \_gnd_net_\,
            in3 => \N__48380\,
            lcout => dds_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51124\,
            ce => \N__48299\,
            sr => \N__48538\
        );

    \comm_spi.data_rx_i0_7344_7345_set_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42236\,
            in1 => \N__45818\,
            in2 => \_gnd_net_\,
            in3 => \N__42260\,
            lcout => \comm_spi.n10455\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42371\,
            ce => 'H',
            sr => \N__42203\
        );

    \ADC_VAC2.i1_3_lut_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001100"
        )
    port map (
            in0 => \N__53482\,
            in1 => \N__35539\,
            in2 => \_gnd_net_\,
            in3 => \N__35636\,
            lcout => \ADC_VAC2.n14926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.adc_state_i1_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36485\,
            in2 => \_gnd_net_\,
            in3 => \N__53483\,
            lcout => adc_state_1_adj_1043,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51145\,
            ce => \N__35510\,
            sr => \N__36521\
        );

    \ADC_VAC2.i7600_2_lut_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__36509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36484\,
            lcout => \ADC_VAC2.n10706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i7328_3_lut_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__38465\,
            in1 => \N__37967\,
            in2 => \_gnd_net_\,
            in3 => \N__51335\,
            lcout => \comm_spi.iclk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i2_3_lut_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__36341\,
            in1 => \N__36357\,
            in2 => \_gnd_net_\,
            in3 => \N__36319\,
            lcout => \comm_spi.n12175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.bit_cnt_1603__i3_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__36359\,
            in1 => \N__38419\,
            in2 => \N__36326\,
            in3 => \N__36344\,
            lcout => \comm_spi.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_1603__i3C_net\,
            ce => 'H',
            sr => \N__46584\
        );

    \comm_spi.bit_cnt_1603__i2_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__36343\,
            in1 => \N__36322\,
            in2 => \_gnd_net_\,
            in3 => \N__36358\,
            lcout => \comm_spi.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_1603__i3C_net\,
            ce => 'H',
            sr => \N__46584\
        );

    \comm_spi.bit_cnt_1603__i1_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36342\,
            lcout => \comm_spi.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_1603__i3C_net\,
            ce => 'H',
            sr => \N__46584\
        );

    \comm_spi.bit_cnt_1603__i0_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36320\,
            lcout => \comm_spi.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_1603__i3C_net\,
            ce => 'H',
            sr => \N__46584\
        );

    \i12087_2_lut_3_lut_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__43445\,
            in1 => \N__50501\,
            in2 => \_gnd_net_\,
            in3 => \N__43267\,
            lcout => n15290,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_282_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__43268\,
            in1 => \N__43447\,
            in2 => \_gnd_net_\,
            in3 => \N__50499\,
            lcout => n4_adj_1179,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_175_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__43446\,
            in1 => \N__50500\,
            in2 => \_gnd_net_\,
            in3 => \N__43265\,
            lcout => n15198,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_3_lut_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__43266\,
            in1 => \N__43448\,
            in2 => \_gnd_net_\,
            in3 => \N__50498\,
            lcout => n8530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_378_Mux_1_i8_3_lut_4_lut_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110001101"
        )
    port map (
            in0 => \N__50510\,
            in1 => \N__49774\,
            in2 => \N__39443\,
            in3 => \N__36548\,
            lcout => n8_adj_1201,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12842_2_lut_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50509\,
            in2 => \_gnd_net_\,
            in3 => \N__42706\,
            lcout => OPEN,
            ltout => \n15668_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_1__bdd_4_lut_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__39040\,
            in1 => \N__49773\,
            in2 => \N__36551\,
            in3 => \N__49480\,
            lcout => n16464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i244_2_lut_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__43287\,
            in1 => \_gnd_net_\,
            in2 => \N__43438\,
            in3 => \_gnd_net_\,
            lcout => n1523,
            ltout => \n1523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_378_Mux_1_i2_3_lut_4_lut_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__50511\,
            in1 => \N__43406\,
            in2 => \N__36542\,
            in3 => \N__49775\,
            lcout => OPEN,
            ltout => \n2_adj_1200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n16464_bdd_4_lut_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__49481\,
            in1 => \N__50512\,
            in2 => \N__36539\,
            in3 => \N__36536\,
            lcout => OPEN,
            ltout => \n16467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i1_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51927\,
            in1 => \N__52066\,
            in2 => \N__36530\,
            in3 => \N__36527\,
            lcout => comm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51170\,
            ce => \N__36620\,
            sr => \_gnd_net_\
        );

    \i13037_4_lut_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110111"
        )
    port map (
            in0 => \N__36629\,
            in1 => \N__50508\,
            in2 => \N__52165\,
            in3 => \N__36557\,
            lcout => n14_adj_1189,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_407_i13_2_lut_3_lut_4_lut_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__47509\,
            in1 => \N__45415\,
            in2 => \N__39013\,
            in3 => \N__45224\,
            lcout => n13_adj_1032,
            ltout => \n13_adj_1032_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_249_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43165\,
            in2 => \N__36599\,
            in3 => \N__50502\,
            lcout => n8519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_246_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47048\,
            in2 => \_gnd_net_\,
            in3 => \N__40862\,
            lcout => n12_adj_1027,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_63_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__40863\,
            in1 => \N__47508\,
            in2 => \N__47183\,
            in3 => \N__45454\,
            lcout => n22_adj_1115,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i3_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011101110"
        )
    port map (
            in0 => \N__40965\,
            in1 => \N__41314\,
            in2 => \N__43916\,
            in3 => \N__52302\,
            lcout => buf_dds_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_296_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__40861\,
            in1 => \N__44967\,
            in2 => \N__47184\,
            in3 => \N__43188\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12836_2_lut_3_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__47507\,
            in1 => \N__45414\,
            in2 => \_gnd_net_\,
            in3 => \N__45223\,
            lcout => n15651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12628_3_lut_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__43449\,
            in1 => \N__43289\,
            in2 => \_gnd_net_\,
            in3 => \N__49741\,
            lcout => n15526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12680_4_lut_4_lut_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46908\,
            in1 => \N__40196\,
            in2 => \N__36972\,
            in3 => \N__37687\,
            lcout => n15584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_115_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__40195\,
            in1 => \N__47594\,
            in2 => \N__37016\,
            in3 => \N__46909\,
            lcout => OPEN,
            ltout => \n8058_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_271_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__45279\,
            in1 => \N__46911\,
            in2 => \N__36998\,
            in3 => \N__36973\,
            lcout => OPEN,
            ltout => \n83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12771_4_lut_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__45537\,
            in1 => \N__36896\,
            in2 => \N__36890\,
            in3 => \N__47595\,
            lcout => n15581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i21_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__44404\,
            in1 => \N__49268\,
            in2 => \N__36844\,
            in3 => \N__36877\,
            lcout => buf_adcdata3_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_301_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__45536\,
            in1 => \N__39410\,
            in2 => \N__40224\,
            in3 => \N__40753\,
            lcout => \comm_state_3_N_402_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i15_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44403\,
            in1 => \N__49267\,
            in2 => \N__36806\,
            in3 => \N__36762\,
            lcout => buf_adcdata3_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i129_4_lut_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__36743\,
            in1 => \N__47593\,
            in2 => \N__37169\,
            in3 => \N__45278\,
            lcout => n75_adj_1164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_idxvec_i0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__37049\,
            in1 => \N__51893\,
            in2 => \N__36705\,
            in3 => \N__52301\,
            lcout => data_idxvec_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51223\,
            ce => \N__37556\,
            sr => \_gnd_net_\
        );

    \mux_1494_i1_3_lut_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37060\,
            in1 => \N__47540\,
            in2 => \_gnd_net_\,
            in3 => \N__36653\,
            lcout => OPEN,
            ltout => \n4197_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i1_4_lut_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__47541\,
            in1 => \N__37145\,
            in2 => \N__37127\,
            in3 => \N__45183\,
            lcout => OPEN,
            ltout => \n4234_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i1_3_lut_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37124\,
            in2 => \N__37112\,
            in3 => \N__45436\,
            lcout => OPEN,
            ltout => \n4254_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i1_4_lut_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__37109\,
            in1 => \N__45184\,
            in2 => \N__37091\,
            in3 => \N__46835\,
            lcout => n4264,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i37_4_lut_4_lut_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001001010010"
        )
    port map (
            in0 => \N__45435\,
            in1 => \N__45182\,
            in2 => \N__47670\,
            in3 => \N__46833\,
            lcout => OPEN,
            ltout => \n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12654_4_lut_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__46834\,
            in1 => \N__40754\,
            in2 => \N__37082\,
            in3 => \N__40164\,
            lcout => n15557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_1441_2_lut_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43615\,
            in2 => \N__37064\,
            in3 => \_gnd_net_\,
            lcout => \data_idxvec_15_N_673_0\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => n14040,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_idxvec_i1_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37492\,
            in1 => \N__38242\,
            in2 => \N__52456\,
            in3 => \N__37043\,
            lcout => data_idxvec_1,
            ltout => OPEN,
            carryin => n14040,
            carryout => n14041,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i2_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__40345\,
            in1 => \N__52394\,
            in2 => \N__37040\,
            in3 => \N__37019\,
            lcout => data_idxvec_2,
            ltout => OPEN,
            carryin => n14041,
            carryout => n14042,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i3_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__43909\,
            in1 => \N__42031\,
            in2 => \N__52457\,
            in3 => \N__37403\,
            lcout => data_idxvec_3,
            ltout => OPEN,
            carryin => n14042,
            carryout => n14043,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i4_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37399\,
            in1 => \N__52398\,
            in2 => \N__37829\,
            in3 => \N__37376\,
            lcout => data_idxvec_4,
            ltout => OPEN,
            carryin => n14043,
            carryout => n14044,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i5_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37373\,
            in1 => \N__38347\,
            in2 => \N__52458\,
            in3 => \N__37349\,
            lcout => data_idxvec_5,
            ltout => OPEN,
            carryin => n14044,
            carryout => n14045,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i6_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37945\,
            in1 => \N__52402\,
            in2 => \N__37345\,
            in3 => \N__37325\,
            lcout => data_idxvec_6,
            ltout => OPEN,
            carryin => n14045,
            carryout => n14046,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i7_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37322\,
            in1 => \N__37294\,
            in2 => \N__52459\,
            in3 => \N__37280\,
            lcout => data_idxvec_7,
            ltout => OPEN,
            carryin => n14046,
            carryout => n14047,
            clk => \N__51240\,
            ce => \N__37552\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i8_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37277\,
            in1 => \N__52406\,
            in2 => \N__41003\,
            in3 => \N__37241\,
            lcout => data_idxvec_8,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => n14048,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i9_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37237\,
            in1 => \N__37207\,
            in2 => \N__52460\,
            in3 => \N__37193\,
            lcout => data_idxvec_9,
            ltout => OPEN,
            carryin => n14048,
            carryout => n14049,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i10_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37189\,
            in1 => \N__52410\,
            in2 => \N__37168\,
            in3 => \N__37148\,
            lcout => data_idxvec_10,
            ltout => OPEN,
            carryin => n14049,
            carryout => n14050,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i11_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__43492\,
            in1 => \N__40579\,
            in2 => \N__52461\,
            in3 => \N__37721\,
            lcout => data_idxvec_11,
            ltout => OPEN,
            carryin => n14050,
            carryout => n14051,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i12_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37711\,
            in1 => \N__52414\,
            in2 => \N__37688\,
            in3 => \N__37670\,
            lcout => data_idxvec_12,
            ltout => OPEN,
            carryin => n14051,
            carryout => n14052,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i13_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37667\,
            in1 => \N__37648\,
            in2 => \N__52462\,
            in3 => \N__37634\,
            lcout => data_idxvec_13,
            ltout => OPEN,
            carryin => n14052,
            carryout => n14053,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i14_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37631\,
            in1 => \N__52418\,
            in2 => \N__37606\,
            in3 => \N__37586\,
            lcout => data_idxvec_14,
            ltout => OPEN,
            carryin => n14053,
            carryout => n14054,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i15_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__52419\,
            in1 => \N__37582\,
            in2 => \N__41675\,
            in3 => \N__37559\,
            lcout => data_idxvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51255\,
            ce => \N__37545\,
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i13_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49077\,
            in1 => \N__44398\,
            in2 => \N__41957\,
            in3 => \N__37516\,
            lcout => buf_adcdata3_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i1_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37496\,
            in1 => \N__40462\,
            in2 => \_gnd_net_\,
            in3 => \N__42161\,
            lcout => req_data_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i14_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53115\,
            in1 => \N__37441\,
            in2 => \N__37475\,
            in3 => \N__52794\,
            lcout => buf_adcdata1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i11_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43493\,
            in1 => \N__40461\,
            in2 => \_gnd_net_\,
            in3 => \N__37422\,
            lcout => req_data_cnt_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i22_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__49078\,
            in1 => \N__41574\,
            in2 => \N__41956\,
            in3 => \N__48810\,
            lcout => cmd_rdadctmp_22_adj_1090,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i6_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37949\,
            in1 => \N__40463\,
            in2 => \_gnd_net_\,
            in3 => \N__37917\,
            lcout => req_data_cnt_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i15_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__38923\,
            in1 => \N__41757\,
            in2 => \N__41657\,
            in3 => \N__51896\,
            lcout => \acadc_skipCount_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i6_3_lut_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37727\,
            in1 => \N__45602\,
            in2 => \_gnd_net_\,
            in3 => \N__38300\,
            lcout => OPEN,
            ltout => \n4249_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i6_4_lut_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__45263\,
            in1 => \N__37901\,
            in2 => \N__37889\,
            in3 => \N__47266\,
            lcout => OPEN,
            ltout => \n4259_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i5_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39765\,
            in1 => \_gnd_net_\,
            in2 => \N__37886\,
            in3 => \N__50289\,
            lcout => comm_buf_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51284\,
            ce => \N__44717\,
            sr => \N__44652\
        );

    \mux_1494_i5_3_lut_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37828\,
            in1 => \N__47792\,
            in2 => \_gnd_net_\,
            in3 => \N__37806\,
            lcout => OPEN,
            ltout => \n4193_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i5_4_lut_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__37790\,
            in1 => \N__47798\,
            in2 => \N__37775\,
            in3 => \N__45261\,
            lcout => n4230,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i6_3_lut_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47799\,
            in1 => \N__37767\,
            in2 => \_gnd_net_\,
            in3 => \N__37748\,
            lcout => n4216,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1494_i6_3_lut_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47793\,
            in1 => \N__38348\,
            in2 => \_gnd_net_\,
            in3 => \N__38331\,
            lcout => OPEN,
            ltout => \n4192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i6_4_lut_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__45262\,
            in1 => \N__38315\,
            in2 => \N__38303\,
            in3 => \N__47794\,
            lcout => n4229,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i10_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53752\,
            in1 => \N__38257\,
            in2 => \N__38294\,
            in3 => \N__53493\,
            lcout => buf_adcdata2_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1494_i2_3_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38243\,
            in1 => \N__38223\,
            in2 => \_gnd_net_\,
            in3 => \N__47791\,
            lcout => n4196,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i17_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38200\,
            in1 => \N__49212\,
            in2 => \N__44535\,
            in3 => \N__48809\,
            lcout => cmd_rdadctmp_17_adj_1095,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i4_3_lut_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47928\,
            in1 => \N__38174\,
            in2 => \_gnd_net_\,
            in3 => \N__38150\,
            lcout => n4218,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7374_2_lut_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38131\,
            in2 => \_gnd_net_\,
            in3 => \N__38047\,
            lcout => n10483,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13067_4_lut_3_lut_LC_18_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46560\,
            in1 => \N__51390\,
            in2 => \_gnd_net_\,
            in3 => \N__37960\,
            lcout => \comm_spi.n16887\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_7326_7327_reset_LC_18_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51397\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n10438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51133\,
            ce => 'H',
            sr => \N__38453\
        );

    \comm_spi.i13087_4_lut_3_lut_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46503\,
            in1 => \N__42889\,
            in2 => \_gnd_net_\,
            in3 => \N__38438\,
            lcout => \comm_spi.n16890\,
            ltout => \comm_spi.n16890_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i7346_3_lut_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38432\,
            in2 => \N__38426\,
            in3 => \N__42473\,
            lcout => comm_rx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i7_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38418\,
            in1 => \N__40628\,
            in2 => \_gnd_net_\,
            in3 => \N__38377\,
            lcout => comm_rx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \comm_spi.data_rx_i6_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38376\,
            in1 => \N__39688\,
            in2 => \_gnd_net_\,
            in3 => \N__38417\,
            lcout => comm_rx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \comm_spi.data_rx_i5_LC_18_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38416\,
            in1 => \N__39832\,
            in2 => \_gnd_net_\,
            in3 => \N__38375\,
            lcout => comm_rx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \comm_spi.data_rx_i4_LC_18_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38374\,
            in1 => \N__44807\,
            in2 => \_gnd_net_\,
            in3 => \N__38415\,
            lcout => comm_rx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \comm_spi.data_rx_i3_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38414\,
            in1 => \N__40021\,
            in2 => \_gnd_net_\,
            in3 => \N__38373\,
            lcout => comm_rx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \comm_spi.data_rx_i2_LC_18_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__38372\,
            in1 => \N__44074\,
            in2 => \_gnd_net_\,
            in3 => \N__38413\,
            lcout => comm_rx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \comm_spi.data_rx_i1_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__38412\,
            in1 => \N__38371\,
            in2 => \_gnd_net_\,
            in3 => \N__39118\,
            lcout => comm_rx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42381\,
            ce => 'H',
            sr => \N__46555\
        );

    \i12171_3_lut_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38978\,
            in1 => \N__38927\,
            in2 => \_gnd_net_\,
            in3 => \N__38689\,
            lcout => n15381,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_378_Mux_3_i7_4_lut_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__49735\,
            in1 => \N__39023\,
            in2 => \N__42748\,
            in3 => \N__49550\,
            lcout => OPEN,
            ltout => \n12846_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i3_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011100000101"
        )
    port map (
            in0 => \N__52033\,
            in1 => \N__51923\,
            in2 => \N__38570\,
            in3 => \N__39425\,
            lcout => comm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51171\,
            ce => \N__38477\,
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_65_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__38567\,
            in1 => \N__39065\,
            in2 => \N__42815\,
            in3 => \N__38486\,
            lcout => n15130,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_276_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100000"
        )
    port map (
            in0 => \N__38533\,
            in1 => \N__39082\,
            in2 => \N__43166\,
            in3 => \N__39073\,
            lcout => OPEN,
            ltout => \n4_adj_1184_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_277_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__49734\,
            in1 => \N__43379\,
            in2 => \N__38501\,
            in3 => \N__50621\,
            lcout => n15108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_174_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__52032\,
            in1 => \N__49733\,
            in2 => \_gnd_net_\,
            in3 => \N__49402\,
            lcout => n15241,
            ltout => \n15241_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_285_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__43205\,
            in1 => \N__38498\,
            in2 => \N__38489\,
            in3 => \N__38485\,
            lcout => n15128,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__43460\,
            in1 => \N__39083\,
            in2 => \_gnd_net_\,
            in3 => \N__39074\,
            lcout => n15266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12200_4_lut_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__39041\,
            in1 => \N__39029\,
            in2 => \N__39050\,
            in3 => \N__49438\,
            lcout => OPEN,
            ltout => \n15410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i0_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__51922\,
            in1 => \_gnd_net_\,
            in2 => \N__39059\,
            in3 => \N__52074\,
            lcout => comm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51189\,
            ce => \N__39056\,
            sr => \_gnd_net_\
        );

    \i12198_3_lut_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010101"
        )
    port map (
            in0 => \N__50507\,
            in1 => \N__43391\,
            in2 => \_gnd_net_\,
            in3 => \N__49939\,
            lcout => n15408,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7283_2_lut_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111011"
        )
    port map (
            in0 => \N__43394\,
            in1 => \N__50506\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n10394,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12980_3_lut_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__42727\,
            in1 => \N__49938\,
            in2 => \_gnd_net_\,
            in3 => \N__39254\,
            lcout => n16190,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12728_2_lut_3_lut_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__43392\,
            in1 => \N__42726\,
            in2 => \_gnd_net_\,
            in3 => \N__50558\,
            lcout => n15635,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i22_3_lut_4_lut_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000001010"
        )
    port map (
            in0 => \N__50505\,
            in1 => \N__43393\,
            in2 => \N__50143\,
            in3 => \N__43288\,
            lcout => n7_adj_1190,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9584_3_lut_4_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__44968\,
            in1 => \N__47496\,
            in2 => \N__39017\,
            in3 => \N__40944\,
            lcout => n12622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i31_3_lut_4_lut_3_lut_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__45410\,
            in1 => \N__47491\,
            in2 => \_gnd_net_\,
            in3 => \N__45221\,
            lcout => n14_adj_1152,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_53_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011100000"
        )
    port map (
            in0 => \N__46963\,
            in1 => \N__39552\,
            in2 => \N__40225\,
            in3 => \N__45413\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12103_3_lut_4_lut_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__45412\,
            in1 => \N__47495\,
            in2 => \N__47181\,
            in3 => \N__40860\,
            lcout => OPEN,
            ltout => \n15309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_39_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39452\,
            in1 => \N__39416\,
            in2 => \N__39446\,
            in3 => \N__40793\,
            lcout => \comm_state_3_N_418_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12762_2_lut_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50513\,
            in2 => \_gnd_net_\,
            in3 => \N__39436\,
            lcout => n15637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_119_i13_2_lut_3_lut_4_lut_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__45222\,
            in1 => \N__45411\,
            in2 => \N__47601\,
            in3 => \N__41211\,
            lcout => n13_adj_1040,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__45455\,
            in1 => \N__45041\,
            in2 => \N__47741\,
            in3 => \N__46898\,
            lcout => n22_adj_1078,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i7_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__44035\,
            in1 => \N__43995\,
            in2 => \N__39255\,
            in3 => \N__39307\,
            lcout => comm_cmd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i0_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__47599\,
            in1 => \N__44032\,
            in2 => \N__44002\,
            in3 => \N__39142\,
            lcout => comm_cmd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i2_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__44033\,
            in1 => \N__43994\,
            in2 => \N__45465\,
            in3 => \N__40036\,
            lcout => comm_cmd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_114_i8_2_lut_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45405\,
            in2 => \_gnd_net_\,
            in3 => \N__45040\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i2_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__39998\,
            in1 => \N__43681\,
            in2 => \N__41519\,
            in3 => \N__41378\,
            lcout => buf_dds_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7266_2_lut_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52082\,
            in2 => \_gnd_net_\,
            in3 => \N__49965\,
            lcout => n10363,
            ltout => \n10363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i4_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__44034\,
            in1 => \N__39878\,
            in2 => \N__39812\,
            in3 => \N__40288\,
            lcout => comm_cmd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i3_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__43996\,
            in1 => \N__44039\,
            in2 => \N__44883\,
            in3 => \N__46818\,
            lcout => comm_cmd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i5_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__40303\,
            in1 => \N__43997\,
            in2 => \N__39731\,
            in3 => \N__44041\,
            lcout => comm_cmd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_6__355_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__39665\,
            in1 => \N__41895\,
            in2 => \N__42986\,
            in3 => \N__41126\,
            lcout => buf_control_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__40302\,
            in1 => \N__40284\,
            in2 => \_gnd_net_\,
            in3 => \N__40266\,
            lcout => n8085,
            ltout => \n8085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_251_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47488\,
            in2 => \N__39593\,
            in3 => \N__46817\,
            lcout => n8094,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_2_lut_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__47489\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45058\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i6_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__40267\,
            in1 => \N__40657\,
            in2 => \N__44003\,
            in3 => \N__44040\,
            lcout => comm_cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i129_4_lut_adj_104_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__47490\,
            in1 => \N__40595\,
            in2 => \N__40583\,
            in3 => \N__45059\,
            lcout => n75,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_300_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46819\,
            in2 => \_gnd_net_\,
            in3 => \N__40830\,
            lcout => n12,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2992_3_lut_4_lut_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__50537\,
            in1 => \N__47602\,
            in2 => \N__40550\,
            in3 => \N__40946\,
            lcout => n6301,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9546_2_lut_3_lut_3_lut_3_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110011001"
        )
    port map (
            in0 => \N__47603\,
            in1 => \N__45539\,
            in2 => \_gnd_net_\,
            in3 => \N__45105\,
            lcout => n12702,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i2_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40456\,
            in1 => \N__40349\,
            in2 => \_gnd_net_\,
            in3 => \N__40323\,
            lcout => req_data_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_297_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__40304\,
            in1 => \N__40289\,
            in2 => \_gnd_net_\,
            in3 => \N__40268\,
            lcout => n8043,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__45540\,
            in1 => \N__47604\,
            in2 => \N__45215\,
            in3 => \N__41210\,
            lcout => n7511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i1_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__41368\,
            in1 => \N__41524\,
            in2 => \N__42124\,
            in3 => \N__41097\,
            lcout => buf_dds_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51256\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_84_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__52081\,
            in1 => \N__41180\,
            in2 => \N__51825\,
            in3 => \N__50594\,
            lcout => n8250,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_290_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__45544\,
            in1 => \N__41040\,
            in2 => \N__41002\,
            in3 => \N__45153\,
            lcout => n78_adj_1022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i4_3_lut_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40970\,
            in1 => \N__47636\,
            in2 => \_gnd_net_\,
            in3 => \N__43774\,
            lcout => n4206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12098_3_lut_4_lut_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100101111"
        )
    port map (
            in0 => \N__40945\,
            in1 => \N__41913\,
            in2 => \N__47790\,
            in3 => \N__41200\,
            lcout => n15188,
            ltout => \n15188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__40906\,
            in1 => \N__46931\,
            in2 => \N__40889\,
            in3 => \N__40859\,
            lcout => OPEN,
            ltout => \n6_adj_1171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_4_lut_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011100000"
        )
    port map (
            in0 => \N__45154\,
            in1 => \N__43636\,
            in2 => \N__40796\,
            in3 => \N__45545\,
            lcout => n15190,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i12_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__49220\,
            in1 => \N__44382\,
            in2 => \N__40782\,
            in3 => \N__48598\,
            lcout => buf_adcdata3_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i21_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__41949\,
            in1 => \N__49221\,
            in2 => \N__48599\,
            in3 => \N__48832\,
            lcout => cmd_rdadctmp_21_adj_1091,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9560_2_lut_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45541\,
            in2 => \_gnd_net_\,
            in3 => \N__45151\,
            lcout => n4_adj_1041,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i14_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__41894\,
            in1 => \N__41756\,
            in2 => \N__51930\,
            in3 => \N__41697\,
            lcout => \acadc_skipCount_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12647_4_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__45542\,
            in1 => \N__46946\,
            in2 => \N__41674\,
            in3 => \N__41652\,
            lcout => n15468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i5_3_lut_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41615\,
            in1 => \N__45543\,
            in2 => \_gnd_net_\,
            in3 => \N__41606\,
            lcout => n4250,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i14_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__41550\,
            in1 => \N__41578\,
            in2 => \N__49266\,
            in3 => \N__44399\,
            lcout => buf_adcdata3_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds_i11_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__43562\,
            in1 => \N__41241\,
            in2 => \N__41528\,
            in3 => \N__41379\,
            lcout => buf_dds_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_208_i13_2_lut_3_lut_4_lut_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__45234\,
            in1 => \N__45605\,
            in2 => \N__41222\,
            in3 => \N__47795\,
            lcout => n13_adj_1025,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1502_i2_3_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47797\,
            in1 => \N__42191\,
            in2 => \_gnd_net_\,
            in3 => \N__42160\,
            lcout => OPEN,
            ltout => \n4220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i2_3_lut_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42041\,
            in2 => \N__42143\,
            in3 => \N__45606\,
            lcout => OPEN,
            ltout => \n4253_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i2_4_lut_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__42068\,
            in1 => \N__45235\,
            in2 => \N__42140\,
            in3 => \N__46965\,
            lcout => n4263,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i2_3_lut_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42120\,
            in1 => \N__42088\,
            in2 => \_gnd_net_\,
            in3 => \N__47796\,
            lcout => n4208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i2_4_lut_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__47800\,
            in1 => \N__45236\,
            in2 => \N__42062\,
            in3 => \N__42047\,
            lcout => n4233,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1494_i4_3_lut_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42035\,
            in1 => \N__47802\,
            in2 => \_gnd_net_\,
            in3 => \N__42017\,
            lcout => OPEN,
            ltout => \n4194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1507_i4_4_lut_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__45237\,
            in1 => \N__41996\,
            in2 => \N__41981\,
            in3 => \N__47801\,
            lcout => OPEN,
            ltout => \n4231_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1511_i4_3_lut_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41978\,
            in2 => \N__41972\,
            in3 => \N__45607\,
            lcout => OPEN,
            ltout => \n4251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1513_i4_4_lut_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__45238\,
            in1 => \N__41969\,
            in2 => \N__41960\,
            in3 => \N__46966\,
            lcout => n4261,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1457_i2_4_lut_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__42686\,
            in1 => \N__47803\,
            in2 => \N__42674\,
            in3 => \N__46964\,
            lcout => n4063,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i11_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53810\,
            in1 => \N__53492\,
            in2 => \N__46181\,
            in3 => \N__42616\,
            lcout => buf_adcdata2_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_8_i15_4_lut_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__52183\,
            in1 => \N__42602\,
            in2 => \N__51929\,
            in3 => \N__42581\,
            lcout => \data_index_9_N_258_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_7330_7331_set_LC_19_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45795\,
            lcout => \comm_spi.n10441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51146\,
            ce => 'H',
            sr => \N__42953\
        );

    \comm_spi.data_rx_i0_7344_7345_reset_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42228\,
            in1 => \N__42253\,
            in2 => \_gnd_net_\,
            in3 => \N__45814\,
            lcout => \comm_spi.n10456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42375\,
            ce => 'H',
            sr => \N__42878\
        );

    \comm_spi.i13072_4_lut_3_lut_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45797\,
            in1 => \N__46462\,
            in2 => \_gnd_net_\,
            in3 => \N__42252\,
            lcout => \comm_spi.n16893\,
            ltout => \comm_spi.n16893_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i7332_3_lut_LC_19_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42232\,
            in2 => \N__42209\,
            in3 => \N__45813\,
            lcout => \comm_spi.imosi\,
            ltout => \comm_spi.imosi_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_86_2_lut_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42206\,
            in3 => \N__46464\,
            lcout => \comm_spi.DOUT_7__N_785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_88_2_lut_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46463\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45796\,
            lcout => \comm_spi.imosi_N_791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i1_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53751\,
            in1 => \N__42904\,
            in2 => \N__42944\,
            in3 => \N__53533\,
            lcout => buf_adcdata2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_87_2_lut_LC_19_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46465\,
            in2 => \_gnd_net_\,
            in3 => \N__42890\,
            lcout => \comm_spi.DOUT_7__N_786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_274_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__42849\,
            in1 => \N__42811\,
            in2 => \N__50550\,
            in3 => \N__43614\,
            lcout => n15191,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2727_2_lut_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__50476\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50282\,
            lcout => n10148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_clear_330_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__50283\,
            in1 => \N__50477\,
            in2 => \_gnd_net_\,
            in3 => \N__52073\,
            lcout => comm_clear,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51190\,
            ce => \N__50633\,
            sr => \_gnd_net_\
        );

    \i22_4_lut_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100010"
        )
    port map (
            in0 => \N__49434\,
            in1 => \N__50559\,
            in2 => \N__42731\,
            in3 => \N__43301\,
            lcout => n8_adj_1193,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12879_4_lut_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001001100"
        )
    port map (
            in0 => \N__50560\,
            in1 => \N__49435\,
            in2 => \N__43436\,
            in3 => \N__42707\,
            lcout => OPEN,
            ltout => \n15711_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i2_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__50286\,
            in1 => \N__43398\,
            in2 => \N__42695\,
            in3 => \N__42692\,
            lcout => comm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51207\,
            ce => \N__43469\,
            sr => \N__52424\
        );

    \i1_4_lut_adj_41_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010111100"
        )
    port map (
            in0 => \N__43300\,
            in1 => \N__50285\,
            in2 => \N__43437\,
            in3 => \N__49433\,
            lcout => OPEN,
            ltout => \n26_adj_1192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13040_2_lut_3_lut_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011111"
        )
    port map (
            in0 => \N__50504\,
            in1 => \N__52062\,
            in2 => \N__43472\,
            in3 => \_gnd_net_\,
            lcout => n18_adj_1191,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_229_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__52061\,
            in1 => \N__50284\,
            in2 => \_gnd_net_\,
            in3 => \N__49432\,
            lcout => n15245,
            ltout => \n15245_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111100"
        )
    port map (
            in0 => \N__50503\,
            in1 => \N__43402\,
            in2 => \N__43304\,
            in3 => \N__43299\,
            lcout => n8544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_206_i9_2_lut_3_lut_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__47542\,
            in1 => \N__45437\,
            in2 => \_gnd_net_\,
            in3 => \N__45225\,
            lcout => n9_adj_1028,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_177_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__52185\,
            in1 => \N__50093\,
            in2 => \_gnd_net_\,
            in3 => \N__49403\,
            lcout => n9011,
            ltout => \n9011_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_287_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__49404\,
            in1 => \N__52186\,
            in2 => \N__43142\,
            in3 => \N__45689\,
            lcout => n9215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1469_i4_4_lut_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100000"
        )
    port map (
            in0 => \N__43040\,
            in1 => \N__47543\,
            in2 => \N__47182\,
            in3 => \N__43024\,
            lcout => \comm_buf_3_7_N_501_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i111_4_lut_adj_133_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__43707\,
            in1 => \N__45464\,
            in2 => \N__42985\,
            in3 => \N__46910\,
            lcout => n60,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i0_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__44400\,
            in1 => \N__43800\,
            in2 => \N__43853\,
            in3 => \N__49265\,
            lcout => buf_adcdata3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i11_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49262\,
            in1 => \N__44401\,
            in2 => \N__49286\,
            in3 => \N__43767\,
            lcout => buf_adcdata3_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i22_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__44402\,
            in1 => \N__49263\,
            in2 => \N__43748\,
            in3 => \N__43708\,
            lcout => buf_adcdata3_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_4_lut_adj_272_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__50108\,
            in1 => \N__49469\,
            in2 => \N__52423\,
            in3 => \N__43694\,
            lcout => n8618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1498_i3_3_lut_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43677\,
            in1 => \N__44199\,
            in2 => \_gnd_net_\,
            in3 => \N__47600\,
            lcout => n4207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i19_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__44509\,
            in1 => \N__49281\,
            in2 => \N__48845\,
            in3 => \N__49264\,
            lcout => cmd_rdadctmp_19_adj_1093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51242\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13023_2_lut_3_lut_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__43635\,
            in1 => \N__45409\,
            in2 => \_gnd_net_\,
            in3 => \N__45042\,
            lcout => n729,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i19_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53774\,
            in1 => \N__43576\,
            in2 => \N__43877\,
            in3 => \N__53569\,
            lcout => buf_adcdata2_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9629_2_lut_3_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__50106\,
            in1 => \N__43559\,
            in2 => \_gnd_net_\,
            in3 => \N__49445\,
            lcout => n14_adj_1208,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i2_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53116\,
            in1 => \N__44419\,
            in2 => \N__44471\,
            in3 => \N__52892\,
            lcout => buf_adcdata1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.ADC_DATA_i10_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__44405\,
            in1 => \N__49243\,
            in2 => \N__44206\,
            in3 => \N__44510\,
            lcout => buf_adcdata3_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i1_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__45043\,
            in1 => \N__44139\,
            in2 => \N__44042\,
            in3 => \N__44001\,
            lcout => comm_cmd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51257\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i26_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53534\,
            in1 => \N__43967\,
            in2 => \N__43892\,
            in3 => \N__46115\,
            lcout => cmd_rdadctmp_26_adj_1050,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i18_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__53813\,
            in1 => \N__53536\,
            in2 => \N__43936\,
            in3 => \N__43891\,
            lcout => buf_adcdata2_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9641_2_lut_3_lut_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44764\,
            in1 => \N__50107\,
            in2 => \_gnd_net_\,
            in3 => \N__49446\,
            lcout => n14_adj_1215,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i27_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46116\,
            in1 => \N__53537\,
            in2 => \N__43873\,
            in3 => \N__43890\,
            lcout => cmd_rdadctmp_27_adj_1049,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i28_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__53535\,
            in1 => \N__43869\,
            in2 => \N__45730\,
            in3 => \N__46117\,
            lcout => cmd_rdadctmp_28_adj_1048,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i29_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46118\,
            in1 => \N__45726\,
            in2 => \N__46357\,
            in3 => \N__53538\,
            lcout => cmd_rdadctmp_29_adj_1047,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i30_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__46119\,
            in1 => \N__53539\,
            in2 => \N__48202\,
            in3 => \N__46353\,
            lcout => cmd_rdadctmp_30_adj_1046,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_286_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50092\,
            in2 => \_gnd_net_\,
            in3 => \N__50593\,
            lcout => n4_adj_1250,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i12_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53811\,
            in1 => \N__45676\,
            in2 => \N__46145\,
            in3 => \N__53525\,
            lcout => buf_adcdata2_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51286\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_i9_2_lut_3_lut_LC_19_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__47605\,
            in1 => \N__45500\,
            in2 => \_gnd_net_\,
            in3 => \N__45152\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i3_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44884\,
            in1 => \N__50109\,
            in2 => \_gnd_net_\,
            in3 => \N__44786\,
            lcout => comm_buf_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51297\,
            ce => \N__44716\,
            sr => \N__44657\
        );

    \ADC_VAC1.ADC_DATA_i13_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__52894\,
            in1 => \N__53129\,
            in2 => \N__44567\,
            in3 => \N__44603\,
            lcout => buf_adcdata1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i18_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__49213\,
            in1 => \N__44542\,
            in2 => \N__44508\,
            in3 => \N__48830\,
            lcout => cmd_rdadctmp_18_adj_1094,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i13_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53799\,
            in1 => \N__44485\,
            in2 => \N__45908\,
            in3 => \N__53527\,
            lcout => buf_adcdata2_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i12_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53128\,
            in1 => \N__46252\,
            in2 => \N__46292\,
            in3 => \N__52895\,
            lcout => buf_adcdata1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51304\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i9_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53798\,
            in1 => \N__46195\,
            in2 => \N__46238\,
            in3 => \N__53572\,
            lcout => buf_adcdata2_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i20_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__46177\,
            in1 => \N__46108\,
            in2 => \N__46141\,
            in3 => \N__53573\,
            lcout => cmd_rdadctmp_20_adj_1056,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i21_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__53570\,
            in1 => \N__46137\,
            in2 => \N__46120\,
            in3 => \N__45903\,
            lcout => cmd_rdadctmp_21_adj_1055,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.cmd_rdadctmp_i22_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__53571\,
            in1 => \N__53592\,
            in2 => \N__46121\,
            in3 => \N__45904\,
            lcout => cmd_rdadctmp_22_adj_1054,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1469_i8_4_lut_LC_20_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__45890\,
            in1 => \N__47929\,
            in2 => \N__45877\,
            in3 => \N__47267\,
            lcout => n4101,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_7330_7331_reset_LC_20_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45777\,
            lcout => \comm_spi.n10442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51173\,
            ce => 'H',
            sr => \N__45740\
        );

    \comm_spi.RESET_I_0_89_2_lut_LC_20_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__45794\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46470\,
            lcout => \comm_spi.imosi_N_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i20_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53733\,
            in1 => \N__45703\,
            in2 => \N__45734\,
            in3 => \N__53532\,
            lcout => buf_adcdata2_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i23_LC_20_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__53531\,
            in1 => \N__53734\,
            in2 => \N__48158\,
            in3 => \N__48118\,
            lcout => buf_adcdata2_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_1469_i1_4_lut_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__48104\,
            in1 => \N__47854\,
            in2 => \N__47378\,
            in3 => \N__47094\,
            lcout => n4108,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i2_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53754\,
            in1 => \N__46667\,
            in2 => \N__46706\,
            in3 => \N__53575\,
            lcout => buf_adcdata2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_95_2_lut_LC_20_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__46638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46501\,
            lcout => \comm_spi.data_tx_7__N_808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_90_2_lut_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__51374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46469\,
            lcout => \comm_spi.iclk_N_801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i13102_4_lut_3_lut_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46639\,
            in1 => \N__46502\,
            in2 => \_gnd_net_\,
            in3 => \N__46377\,
            lcout => \comm_spi.n16899\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i21_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53753\,
            in1 => \N__46327\,
            in2 => \N__46361\,
            in3 => \N__53574\,
            lcout => buf_adcdata2_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_response_331_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000011010"
        )
    port map (
            in0 => \N__50141\,
            in1 => \N__49406\,
            in2 => \N__52356\,
            in3 => \N__50554\,
            lcout => \ICE_GPMI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51225\,
            ce => \N__49298\,
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_4_lut_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111000010"
        )
    port map (
            in0 => \N__50552\,
            in1 => \N__52220\,
            in2 => \N__50292\,
            in3 => \N__49436\,
            lcout => n8576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111011"
        )
    port map (
            in0 => \N__50553\,
            in1 => \N__52221\,
            in2 => \N__50293\,
            in3 => \_gnd_net_\,
            lcout => n8117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_226_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__52219\,
            in1 => \N__49405\,
            in2 => \_gnd_net_\,
            in3 => \N__50551\,
            lcout => n6_adj_1175,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_4_lut_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011101111"
        )
    port map (
            in0 => \N__50595\,
            in1 => \N__50142\,
            in2 => \N__52390\,
            in3 => \N__49437\,
            lcout => n8129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC3.cmd_rdadctmp_i20_LC_20_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__49285\,
            in1 => \N__49242\,
            in2 => \N__48589\,
            in3 => \N__48841\,
            lcout => cmd_rdadctmp_20_adj_1092,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51243\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLOCK_DDS.dds_state_i0_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000110011"
        )
    port map (
            in0 => \N__48572\,
            in1 => \N__48334\,
            in2 => \N__48563\,
            in3 => \N__48542\,
            lcout => dds_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51258\,
            ce => \N__48298\,
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i16_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53117\,
            in1 => \N__48226\,
            in2 => \N__48272\,
            in3 => \N__52893\,
            lcout => buf_adcdata1_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i22_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__48201\,
            in1 => \N__53775\,
            in2 => \N__53576\,
            in3 => \N__48172\,
            lcout => buf_adcdata2_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51274\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC2.ADC_DATA_i14_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53812\,
            in1 => \N__53143\,
            in2 => \N__53609\,
            in3 => \N__53526\,
            lcout => buf_adcdata2_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC1.ADC_DATA_i10_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__53114\,
            in1 => \N__52504\,
            in2 => \N__52934\,
            in3 => \N__52896\,
            lcout => buf_adcdata1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_394_Mux_5_i15_4_lut_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__52490\,
            in1 => \N__52455\,
            in2 => \N__51932\,
            in3 => \N__51515\,
            lcout => \data_index_9_N_258_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_7326_7327_set_LC_23_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51375\,
            lcout => \comm_spi.n10437\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__51261\,
            ce => 'H',
            sr => \N__50672\
        );
end \INTERFACE\;
