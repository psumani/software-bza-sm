-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 7 2021 19:29:47

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "zim" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of zim
entity zim is
port (
    VAC_DRDY : in std_logic;
    IAC_FLT1 : out std_logic;
    DDS_SCK : out std_logic;
    ICE_IOR_166 : in std_logic;
    ICE_IOR_119 : in std_logic;
    DDS_MOSI : out std_logic;
    VAC_MISO : in std_logic;
    DDS_MOSI1 : out std_logic;
    ICE_IOR_146 : in std_logic;
    VDC_CLK : out std_logic;
    ICE_IOT_222 : in std_logic;
    IAC_CS : out std_logic;
    ICE_IOL_18B : in std_logic;
    ICE_IOL_13A : in std_logic;
    ICE_IOB_81 : in std_logic;
    VAC_OSR1 : out std_logic;
    IAC_MOSI : out std_logic;
    DDS_CS1 : out std_logic;
    ICE_IOL_4B : in std_logic;
    ICE_IOB_94 : in std_logic;
    VAC_CS : out std_logic;
    VAC_CLK : out std_logic;
    ICE_SPI_CE0 : in std_logic;
    ICE_IOR_167 : in std_logic;
    ICE_IOR_118 : in std_logic;
    RTD_SDO : in std_logic;
    IAC_OSR0 : out std_logic;
    VDC_SCLK : out std_logic;
    VAC_FLT1 : out std_logic;
    ICE_SPI_MOSI : in std_logic;
    ICE_IOR_165 : in std_logic;
    ICE_IOR_147 : in std_logic;
    ICE_IOL_14A : in std_logic;
    ICE_IOL_13B : in std_logic;
    ICE_IOB_91 : in std_logic;
    ICE_GPMO_0 : in std_logic;
    DDS_RNG_0 : out std_logic;
    VDC_RNG0 : out std_logic;
    ICE_SPI_SCLK : in std_logic;
    ICE_IOR_152 : in std_logic;
    ICE_IOL_12A : in std_logic;
    RTD_DRDY : in std_logic;
    ICE_SPI_MISO : out std_logic;
    ICE_IOT_177 : in std_logic;
    ICE_IOR_141 : in std_logic;
    ICE_IOB_80 : in std_logic;
    ICE_IOB_102 : in std_logic;
    ICE_GPMO_2 : in std_logic;
    ICE_GPMI_0 : out std_logic;
    IAC_MISO : in std_logic;
    VAC_OSR0 : out std_logic;
    VAC_MOSI : out std_logic;
    TEST_LED : out std_logic;
    ICE_IOR_148 : in std_logic;
    STAT_COMM : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_IOR_161 : in std_logic;
    ICE_IOB_95 : in std_logic;
    ICE_IOB_82 : in std_logic;
    ICE_IOB_104 : in std_logic;
    IAC_CLK : out std_logic;
    DDS_CS : out std_logic;
    SELIRNG0 : out std_logic;
    RTD_SDI : out std_logic;
    ICE_IOT_221 : in std_logic;
    ICE_IOT_197 : in std_logic;
    DDS_MCLK : out std_logic;
    RTD_SCLK : out std_logic;
    RTD_CS : out std_logic;
    ICE_IOR_137 : in std_logic;
    IAC_OSR1 : out std_logic;
    VAC_FLT0 : out std_logic;
    ICE_IOR_144 : in std_logic;
    ICE_IOR_128 : in std_logic;
    ICE_GPMO_1 : in std_logic;
    IAC_SCLK : out std_logic;
    EIS_SYNCCLK : in std_logic;
    ICE_IOR_139 : in std_logic;
    ICE_IOL_4A : in std_logic;
    VAC_SCLK : out std_logic;
    THERMOSTAT : in std_logic;
    ICE_IOR_164 : in std_logic;
    ICE_IOB_103 : in std_logic;
    AMPV_POW : out std_logic;
    VDC_SDO : in std_logic;
    ICE_IOT_174 : in std_logic;
    ICE_IOR_140 : in std_logic;
    ICE_IOB_96 : in std_logic;
    CONT_SD : out std_logic;
    AC_ADC_SYNC : out std_logic;
    SELIRNG1 : out std_logic;
    ICE_IOL_12B : in std_logic;
    ICE_IOR_160 : in std_logic;
    ICE_IOR_136 : in std_logic;
    DDS_MCLK1 : out std_logic;
    ICE_IOT_198 : in std_logic;
    ICE_IOT_173 : in std_logic;
    IAC_DRDY : in std_logic;
    ICE_IOT_178 : in std_logic;
    ICE_IOR_138 : in std_logic;
    ICE_IOR_120 : in std_logic;
    IAC_FLT0 : out std_logic;
    DDS_SCK1 : out std_logic);
end zim;

-- Architecture of zim
-- View name is \INTERFACE\
architecture \INTERFACE\ of zim is

signal \N__59914\ : std_logic;
signal \N__59913\ : std_logic;
signal \N__59912\ : std_logic;
signal \N__59905\ : std_logic;
signal \N__59904\ : std_logic;
signal \N__59903\ : std_logic;
signal \N__59896\ : std_logic;
signal \N__59895\ : std_logic;
signal \N__59894\ : std_logic;
signal \N__59887\ : std_logic;
signal \N__59886\ : std_logic;
signal \N__59885\ : std_logic;
signal \N__59878\ : std_logic;
signal \N__59877\ : std_logic;
signal \N__59876\ : std_logic;
signal \N__59869\ : std_logic;
signal \N__59868\ : std_logic;
signal \N__59867\ : std_logic;
signal \N__59860\ : std_logic;
signal \N__59859\ : std_logic;
signal \N__59858\ : std_logic;
signal \N__59851\ : std_logic;
signal \N__59850\ : std_logic;
signal \N__59849\ : std_logic;
signal \N__59842\ : std_logic;
signal \N__59841\ : std_logic;
signal \N__59840\ : std_logic;
signal \N__59833\ : std_logic;
signal \N__59832\ : std_logic;
signal \N__59831\ : std_logic;
signal \N__59824\ : std_logic;
signal \N__59823\ : std_logic;
signal \N__59822\ : std_logic;
signal \N__59815\ : std_logic;
signal \N__59814\ : std_logic;
signal \N__59813\ : std_logic;
signal \N__59806\ : std_logic;
signal \N__59805\ : std_logic;
signal \N__59804\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59796\ : std_logic;
signal \N__59795\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59787\ : std_logic;
signal \N__59786\ : std_logic;
signal \N__59779\ : std_logic;
signal \N__59778\ : std_logic;
signal \N__59777\ : std_logic;
signal \N__59770\ : std_logic;
signal \N__59769\ : std_logic;
signal \N__59768\ : std_logic;
signal \N__59761\ : std_logic;
signal \N__59760\ : std_logic;
signal \N__59759\ : std_logic;
signal \N__59752\ : std_logic;
signal \N__59751\ : std_logic;
signal \N__59750\ : std_logic;
signal \N__59743\ : std_logic;
signal \N__59742\ : std_logic;
signal \N__59741\ : std_logic;
signal \N__59734\ : std_logic;
signal \N__59733\ : std_logic;
signal \N__59732\ : std_logic;
signal \N__59725\ : std_logic;
signal \N__59724\ : std_logic;
signal \N__59723\ : std_logic;
signal \N__59716\ : std_logic;
signal \N__59715\ : std_logic;
signal \N__59714\ : std_logic;
signal \N__59707\ : std_logic;
signal \N__59706\ : std_logic;
signal \N__59705\ : std_logic;
signal \N__59698\ : std_logic;
signal \N__59697\ : std_logic;
signal \N__59696\ : std_logic;
signal \N__59689\ : std_logic;
signal \N__59688\ : std_logic;
signal \N__59687\ : std_logic;
signal \N__59680\ : std_logic;
signal \N__59679\ : std_logic;
signal \N__59678\ : std_logic;
signal \N__59671\ : std_logic;
signal \N__59670\ : std_logic;
signal \N__59669\ : std_logic;
signal \N__59662\ : std_logic;
signal \N__59661\ : std_logic;
signal \N__59660\ : std_logic;
signal \N__59653\ : std_logic;
signal \N__59652\ : std_logic;
signal \N__59651\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59643\ : std_logic;
signal \N__59642\ : std_logic;
signal \N__59635\ : std_logic;
signal \N__59634\ : std_logic;
signal \N__59633\ : std_logic;
signal \N__59626\ : std_logic;
signal \N__59625\ : std_logic;
signal \N__59624\ : std_logic;
signal \N__59617\ : std_logic;
signal \N__59616\ : std_logic;
signal \N__59615\ : std_logic;
signal \N__59608\ : std_logic;
signal \N__59607\ : std_logic;
signal \N__59606\ : std_logic;
signal \N__59599\ : std_logic;
signal \N__59598\ : std_logic;
signal \N__59597\ : std_logic;
signal \N__59590\ : std_logic;
signal \N__59589\ : std_logic;
signal \N__59588\ : std_logic;
signal \N__59581\ : std_logic;
signal \N__59580\ : std_logic;
signal \N__59579\ : std_logic;
signal \N__59572\ : std_logic;
signal \N__59571\ : std_logic;
signal \N__59570\ : std_logic;
signal \N__59563\ : std_logic;
signal \N__59562\ : std_logic;
signal \N__59561\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59553\ : std_logic;
signal \N__59552\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59544\ : std_logic;
signal \N__59543\ : std_logic;
signal \N__59536\ : std_logic;
signal \N__59535\ : std_logic;
signal \N__59534\ : std_logic;
signal \N__59527\ : std_logic;
signal \N__59526\ : std_logic;
signal \N__59525\ : std_logic;
signal \N__59518\ : std_logic;
signal \N__59517\ : std_logic;
signal \N__59516\ : std_logic;
signal \N__59509\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59507\ : std_logic;
signal \N__59500\ : std_logic;
signal \N__59499\ : std_logic;
signal \N__59498\ : std_logic;
signal \N__59491\ : std_logic;
signal \N__59490\ : std_logic;
signal \N__59489\ : std_logic;
signal \N__59482\ : std_logic;
signal \N__59481\ : std_logic;
signal \N__59480\ : std_logic;
signal \N__59473\ : std_logic;
signal \N__59472\ : std_logic;
signal \N__59471\ : std_logic;
signal \N__59464\ : std_logic;
signal \N__59463\ : std_logic;
signal \N__59462\ : std_logic;
signal \N__59455\ : std_logic;
signal \N__59454\ : std_logic;
signal \N__59453\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59445\ : std_logic;
signal \N__59444\ : std_logic;
signal \N__59437\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59435\ : std_logic;
signal \N__59428\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59419\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59417\ : std_logic;
signal \N__59410\ : std_logic;
signal \N__59409\ : std_logic;
signal \N__59408\ : std_logic;
signal \N__59401\ : std_logic;
signal \N__59400\ : std_logic;
signal \N__59399\ : std_logic;
signal \N__59392\ : std_logic;
signal \N__59391\ : std_logic;
signal \N__59390\ : std_logic;
signal \N__59383\ : std_logic;
signal \N__59382\ : std_logic;
signal \N__59381\ : std_logic;
signal \N__59374\ : std_logic;
signal \N__59373\ : std_logic;
signal \N__59372\ : std_logic;
signal \N__59365\ : std_logic;
signal \N__59364\ : std_logic;
signal \N__59363\ : std_logic;
signal \N__59356\ : std_logic;
signal \N__59355\ : std_logic;
signal \N__59354\ : std_logic;
signal \N__59347\ : std_logic;
signal \N__59346\ : std_logic;
signal \N__59345\ : std_logic;
signal \N__59338\ : std_logic;
signal \N__59337\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59329\ : std_logic;
signal \N__59328\ : std_logic;
signal \N__59327\ : std_logic;
signal \N__59320\ : std_logic;
signal \N__59319\ : std_logic;
signal \N__59318\ : std_logic;
signal \N__59311\ : std_logic;
signal \N__59310\ : std_logic;
signal \N__59309\ : std_logic;
signal \N__59302\ : std_logic;
signal \N__59301\ : std_logic;
signal \N__59300\ : std_logic;
signal \N__59293\ : std_logic;
signal \N__59292\ : std_logic;
signal \N__59291\ : std_logic;
signal \N__59284\ : std_logic;
signal \N__59283\ : std_logic;
signal \N__59282\ : std_logic;
signal \N__59275\ : std_logic;
signal \N__59274\ : std_logic;
signal \N__59273\ : std_logic;
signal \N__59266\ : std_logic;
signal \N__59265\ : std_logic;
signal \N__59264\ : std_logic;
signal \N__59257\ : std_logic;
signal \N__59256\ : std_logic;
signal \N__59255\ : std_logic;
signal \N__59248\ : std_logic;
signal \N__59247\ : std_logic;
signal \N__59246\ : std_logic;
signal \N__59239\ : std_logic;
signal \N__59238\ : std_logic;
signal \N__59237\ : std_logic;
signal \N__59230\ : std_logic;
signal \N__59229\ : std_logic;
signal \N__59228\ : std_logic;
signal \N__59221\ : std_logic;
signal \N__59220\ : std_logic;
signal \N__59219\ : std_logic;
signal \N__59212\ : std_logic;
signal \N__59211\ : std_logic;
signal \N__59210\ : std_logic;
signal \N__59203\ : std_logic;
signal \N__59202\ : std_logic;
signal \N__59201\ : std_logic;
signal \N__59194\ : std_logic;
signal \N__59193\ : std_logic;
signal \N__59192\ : std_logic;
signal \N__59185\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59183\ : std_logic;
signal \N__59176\ : std_logic;
signal \N__59175\ : std_logic;
signal \N__59174\ : std_logic;
signal \N__59167\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59158\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59156\ : std_logic;
signal \N__59149\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59147\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59139\ : std_logic;
signal \N__59138\ : std_logic;
signal \N__59131\ : std_logic;
signal \N__59130\ : std_logic;
signal \N__59129\ : std_logic;
signal \N__59122\ : std_logic;
signal \N__59121\ : std_logic;
signal \N__59120\ : std_logic;
signal \N__59113\ : std_logic;
signal \N__59112\ : std_logic;
signal \N__59111\ : std_logic;
signal \N__59104\ : std_logic;
signal \N__59103\ : std_logic;
signal \N__59102\ : std_logic;
signal \N__59095\ : std_logic;
signal \N__59094\ : std_logic;
signal \N__59093\ : std_logic;
signal \N__59086\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59084\ : std_logic;
signal \N__59077\ : std_logic;
signal \N__59076\ : std_logic;
signal \N__59075\ : std_logic;
signal \N__59068\ : std_logic;
signal \N__59067\ : std_logic;
signal \N__59066\ : std_logic;
signal \N__59059\ : std_logic;
signal \N__59058\ : std_logic;
signal \N__59057\ : std_logic;
signal \N__59050\ : std_logic;
signal \N__59049\ : std_logic;
signal \N__59048\ : std_logic;
signal \N__59041\ : std_logic;
signal \N__59040\ : std_logic;
signal \N__59039\ : std_logic;
signal \N__59032\ : std_logic;
signal \N__59031\ : std_logic;
signal \N__59030\ : std_logic;
signal \N__59023\ : std_logic;
signal \N__59022\ : std_logic;
signal \N__59021\ : std_logic;
signal \N__59014\ : std_logic;
signal \N__59013\ : std_logic;
signal \N__59012\ : std_logic;
signal \N__59005\ : std_logic;
signal \N__59004\ : std_logic;
signal \N__59003\ : std_logic;
signal \N__58996\ : std_logic;
signal \N__58995\ : std_logic;
signal \N__58994\ : std_logic;
signal \N__58977\ : std_logic;
signal \N__58974\ : std_logic;
signal \N__58973\ : std_logic;
signal \N__58972\ : std_logic;
signal \N__58969\ : std_logic;
signal \N__58968\ : std_logic;
signal \N__58965\ : std_logic;
signal \N__58962\ : std_logic;
signal \N__58959\ : std_logic;
signal \N__58956\ : std_logic;
signal \N__58953\ : std_logic;
signal \N__58950\ : std_logic;
signal \N__58945\ : std_logic;
signal \N__58942\ : std_logic;
signal \N__58939\ : std_logic;
signal \N__58934\ : std_logic;
signal \N__58931\ : std_logic;
signal \N__58926\ : std_logic;
signal \N__58923\ : std_logic;
signal \N__58920\ : std_logic;
signal \N__58917\ : std_logic;
signal \N__58914\ : std_logic;
signal \N__58911\ : std_logic;
signal \N__58910\ : std_logic;
signal \N__58907\ : std_logic;
signal \N__58904\ : std_logic;
signal \N__58899\ : std_logic;
signal \N__58896\ : std_logic;
signal \N__58893\ : std_logic;
signal \N__58892\ : std_logic;
signal \N__58891\ : std_logic;
signal \N__58888\ : std_logic;
signal \N__58885\ : std_logic;
signal \N__58882\ : std_logic;
signal \N__58875\ : std_logic;
signal \N__58874\ : std_logic;
signal \N__58871\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58863\ : std_logic;
signal \N__58860\ : std_logic;
signal \N__58857\ : std_logic;
signal \N__58856\ : std_logic;
signal \N__58853\ : std_logic;
signal \N__58850\ : std_logic;
signal \N__58847\ : std_logic;
signal \N__58844\ : std_logic;
signal \N__58839\ : std_logic;
signal \N__58836\ : std_logic;
signal \N__58833\ : std_logic;
signal \N__58830\ : std_logic;
signal \N__58827\ : std_logic;
signal \N__58824\ : std_logic;
signal \N__58821\ : std_logic;
signal \N__58818\ : std_logic;
signal \N__58817\ : std_logic;
signal \N__58816\ : std_logic;
signal \N__58809\ : std_logic;
signal \N__58806\ : std_logic;
signal \N__58803\ : std_logic;
signal \N__58800\ : std_logic;
signal \N__58797\ : std_logic;
signal \N__58796\ : std_logic;
signal \N__58793\ : std_logic;
signal \N__58790\ : std_logic;
signal \N__58789\ : std_logic;
signal \N__58784\ : std_logic;
signal \N__58781\ : std_logic;
signal \N__58776\ : std_logic;
signal \N__58775\ : std_logic;
signal \N__58774\ : std_logic;
signal \N__58773\ : std_logic;
signal \N__58770\ : std_logic;
signal \N__58767\ : std_logic;
signal \N__58766\ : std_logic;
signal \N__58765\ : std_logic;
signal \N__58764\ : std_logic;
signal \N__58763\ : std_logic;
signal \N__58762\ : std_logic;
signal \N__58759\ : std_logic;
signal \N__58758\ : std_logic;
signal \N__58755\ : std_logic;
signal \N__58754\ : std_logic;
signal \N__58753\ : std_logic;
signal \N__58752\ : std_logic;
signal \N__58751\ : std_logic;
signal \N__58750\ : std_logic;
signal \N__58749\ : std_logic;
signal \N__58748\ : std_logic;
signal \N__58747\ : std_logic;
signal \N__58746\ : std_logic;
signal \N__58745\ : std_logic;
signal \N__58744\ : std_logic;
signal \N__58743\ : std_logic;
signal \N__58738\ : std_logic;
signal \N__58735\ : std_logic;
signal \N__58732\ : std_logic;
signal \N__58729\ : std_logic;
signal \N__58728\ : std_logic;
signal \N__58725\ : std_logic;
signal \N__58722\ : std_logic;
signal \N__58721\ : std_logic;
signal \N__58720\ : std_logic;
signal \N__58719\ : std_logic;
signal \N__58718\ : std_logic;
signal \N__58717\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58715\ : std_logic;
signal \N__58712\ : std_logic;
signal \N__58709\ : std_logic;
signal \N__58708\ : std_logic;
signal \N__58707\ : std_logic;
signal \N__58706\ : std_logic;
signal \N__58705\ : std_logic;
signal \N__58704\ : std_logic;
signal \N__58703\ : std_logic;
signal \N__58702\ : std_logic;
signal \N__58699\ : std_logic;
signal \N__58696\ : std_logic;
signal \N__58695\ : std_logic;
signal \N__58692\ : std_logic;
signal \N__58691\ : std_logic;
signal \N__58688\ : std_logic;
signal \N__58687\ : std_logic;
signal \N__58684\ : std_logic;
signal \N__58683\ : std_logic;
signal \N__58680\ : std_logic;
signal \N__58679\ : std_logic;
signal \N__58676\ : std_logic;
signal \N__58675\ : std_logic;
signal \N__58672\ : std_logic;
signal \N__58671\ : std_logic;
signal \N__58668\ : std_logic;
signal \N__58665\ : std_logic;
signal \N__58664\ : std_logic;
signal \N__58661\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58657\ : std_logic;
signal \N__58656\ : std_logic;
signal \N__58653\ : std_logic;
signal \N__58644\ : std_logic;
signal \N__58641\ : std_logic;
signal \N__58636\ : std_logic;
signal \N__58633\ : std_logic;
signal \N__58630\ : std_logic;
signal \N__58627\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58622\ : std_logic;
signal \N__58619\ : std_logic;
signal \N__58618\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58614\ : std_logic;
signal \N__58611\ : std_logic;
signal \N__58608\ : std_logic;
signal \N__58605\ : std_logic;
signal \N__58598\ : std_logic;
signal \N__58589\ : std_logic;
signal \N__58586\ : std_logic;
signal \N__58571\ : std_logic;
signal \N__58554\ : std_logic;
signal \N__58539\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58508\ : std_logic;
signal \N__58503\ : std_logic;
signal \N__58498\ : std_logic;
signal \N__58495\ : std_logic;
signal \N__58490\ : std_logic;
signal \N__58487\ : std_logic;
signal \N__58486\ : std_logic;
signal \N__58481\ : std_logic;
signal \N__58478\ : std_logic;
signal \N__58475\ : std_logic;
signal \N__58472\ : std_logic;
signal \N__58469\ : std_logic;
signal \N__58466\ : std_logic;
signal \N__58463\ : std_logic;
signal \N__58460\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58450\ : std_logic;
signal \N__58441\ : std_logic;
signal \N__58438\ : std_logic;
signal \N__58431\ : std_logic;
signal \N__58430\ : std_logic;
signal \N__58427\ : std_logic;
signal \N__58424\ : std_logic;
signal \N__58421\ : std_logic;
signal \N__58418\ : std_logic;
signal \N__58413\ : std_logic;
signal \N__58412\ : std_logic;
signal \N__58409\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58407\ : std_logic;
signal \N__58406\ : std_logic;
signal \N__58403\ : std_logic;
signal \N__58402\ : std_logic;
signal \N__58401\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58399\ : std_logic;
signal \N__58396\ : std_logic;
signal \N__58393\ : std_logic;
signal \N__58392\ : std_logic;
signal \N__58391\ : std_logic;
signal \N__58388\ : std_logic;
signal \N__58385\ : std_logic;
signal \N__58384\ : std_logic;
signal \N__58381\ : std_logic;
signal \N__58378\ : std_logic;
signal \N__58375\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58371\ : std_logic;
signal \N__58368\ : std_logic;
signal \N__58367\ : std_logic;
signal \N__58362\ : std_logic;
signal \N__58359\ : std_logic;
signal \N__58358\ : std_logic;
signal \N__58357\ : std_logic;
signal \N__58356\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58352\ : std_logic;
signal \N__58347\ : std_logic;
signal \N__58344\ : std_logic;
signal \N__58341\ : std_logic;
signal \N__58338\ : std_logic;
signal \N__58337\ : std_logic;
signal \N__58332\ : std_logic;
signal \N__58329\ : std_logic;
signal \N__58328\ : std_logic;
signal \N__58325\ : std_logic;
signal \N__58322\ : std_logic;
signal \N__58317\ : std_logic;
signal \N__58314\ : std_logic;
signal \N__58311\ : std_logic;
signal \N__58308\ : std_logic;
signal \N__58307\ : std_logic;
signal \N__58304\ : std_logic;
signal \N__58301\ : std_logic;
signal \N__58298\ : std_logic;
signal \N__58295\ : std_logic;
signal \N__58290\ : std_logic;
signal \N__58287\ : std_logic;
signal \N__58284\ : std_logic;
signal \N__58281\ : std_logic;
signal \N__58278\ : std_logic;
signal \N__58273\ : std_logic;
signal \N__58270\ : std_logic;
signal \N__58267\ : std_logic;
signal \N__58264\ : std_logic;
signal \N__58261\ : std_logic;
signal \N__58258\ : std_logic;
signal \N__58257\ : std_logic;
signal \N__58252\ : std_logic;
signal \N__58243\ : std_logic;
signal \N__58236\ : std_logic;
signal \N__58231\ : std_logic;
signal \N__58222\ : std_logic;
signal \N__58219\ : std_logic;
signal \N__58216\ : std_logic;
signal \N__58211\ : std_logic;
signal \N__58206\ : std_logic;
signal \N__58203\ : std_logic;
signal \N__58194\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58192\ : std_logic;
signal \N__58187\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58178\ : std_logic;
signal \N__58173\ : std_logic;
signal \N__58170\ : std_logic;
signal \N__58167\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58165\ : std_logic;
signal \N__58164\ : std_logic;
signal \N__58163\ : std_logic;
signal \N__58162\ : std_logic;
signal \N__58161\ : std_logic;
signal \N__58160\ : std_logic;
signal \N__58159\ : std_logic;
signal \N__58158\ : std_logic;
signal \N__58157\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58150\ : std_logic;
signal \N__58149\ : std_logic;
signal \N__58146\ : std_logic;
signal \N__58145\ : std_logic;
signal \N__58140\ : std_logic;
signal \N__58139\ : std_logic;
signal \N__58136\ : std_logic;
signal \N__58133\ : std_logic;
signal \N__58132\ : std_logic;
signal \N__58131\ : std_logic;
signal \N__58128\ : std_logic;
signal \N__58127\ : std_logic;
signal \N__58126\ : std_logic;
signal \N__58123\ : std_logic;
signal \N__58122\ : std_logic;
signal \N__58121\ : std_logic;
signal \N__58120\ : std_logic;
signal \N__58117\ : std_logic;
signal \N__58114\ : std_logic;
signal \N__58113\ : std_logic;
signal \N__58110\ : std_logic;
signal \N__58109\ : std_logic;
signal \N__58108\ : std_logic;
signal \N__58101\ : std_logic;
signal \N__58098\ : std_logic;
signal \N__58095\ : std_logic;
signal \N__58092\ : std_logic;
signal \N__58081\ : std_logic;
signal \N__58074\ : std_logic;
signal \N__58071\ : std_logic;
signal \N__58068\ : std_logic;
signal \N__58067\ : std_logic;
signal \N__58066\ : std_logic;
signal \N__58065\ : std_logic;
signal \N__58060\ : std_logic;
signal \N__58059\ : std_logic;
signal \N__58058\ : std_logic;
signal \N__58055\ : std_logic;
signal \N__58054\ : std_logic;
signal \N__58053\ : std_logic;
signal \N__58052\ : std_logic;
signal \N__58051\ : std_logic;
signal \N__58048\ : std_logic;
signal \N__58045\ : std_logic;
signal \N__58038\ : std_logic;
signal \N__58035\ : std_logic;
signal \N__58030\ : std_logic;
signal \N__58023\ : std_logic;
signal \N__58018\ : std_logic;
signal \N__58013\ : std_logic;
signal \N__58010\ : std_logic;
signal \N__58007\ : std_logic;
signal \N__58002\ : std_logic;
signal \N__57999\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57989\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57987\ : std_logic;
signal \N__57982\ : std_logic;
signal \N__57979\ : std_logic;
signal \N__57976\ : std_logic;
signal \N__57973\ : std_logic;
signal \N__57970\ : std_logic;
signal \N__57967\ : std_logic;
signal \N__57960\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57945\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57935\ : std_logic;
signal \N__57932\ : std_logic;
signal \N__57929\ : std_logic;
signal \N__57926\ : std_logic;
signal \N__57919\ : std_logic;
signal \N__57916\ : std_logic;
signal \N__57903\ : std_logic;
signal \N__57900\ : std_logic;
signal \N__57897\ : std_logic;
signal \N__57896\ : std_logic;
signal \N__57893\ : std_logic;
signal \N__57890\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57882\ : std_logic;
signal \N__57879\ : std_logic;
signal \N__57878\ : std_logic;
signal \N__57875\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57866\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57855\ : std_logic;
signal \N__57854\ : std_logic;
signal \N__57851\ : std_logic;
signal \N__57848\ : std_logic;
signal \N__57845\ : std_logic;
signal \N__57840\ : std_logic;
signal \N__57837\ : std_logic;
signal \N__57836\ : std_logic;
signal \N__57833\ : std_logic;
signal \N__57830\ : std_logic;
signal \N__57827\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57819\ : std_logic;
signal \N__57816\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57812\ : std_logic;
signal \N__57809\ : std_logic;
signal \N__57806\ : std_logic;
signal \N__57803\ : std_logic;
signal \N__57798\ : std_logic;
signal \N__57795\ : std_logic;
signal \N__57794\ : std_logic;
signal \N__57791\ : std_logic;
signal \N__57788\ : std_logic;
signal \N__57785\ : std_logic;
signal \N__57782\ : std_logic;
signal \N__57777\ : std_logic;
signal \N__57774\ : std_logic;
signal \N__57773\ : std_logic;
signal \N__57770\ : std_logic;
signal \N__57767\ : std_logic;
signal \N__57764\ : std_logic;
signal \N__57759\ : std_logic;
signal \N__57756\ : std_logic;
signal \N__57753\ : std_logic;
signal \N__57750\ : std_logic;
signal \N__57749\ : std_logic;
signal \N__57746\ : std_logic;
signal \N__57743\ : std_logic;
signal \N__57740\ : std_logic;
signal \N__57735\ : std_logic;
signal \N__57734\ : std_logic;
signal \N__57731\ : std_logic;
signal \N__57728\ : std_logic;
signal \N__57725\ : std_logic;
signal \N__57722\ : std_logic;
signal \N__57719\ : std_logic;
signal \N__57714\ : std_logic;
signal \N__57713\ : std_logic;
signal \N__57710\ : std_logic;
signal \N__57707\ : std_logic;
signal \N__57704\ : std_logic;
signal \N__57699\ : std_logic;
signal \N__57696\ : std_logic;
signal \N__57695\ : std_logic;
signal \N__57692\ : std_logic;
signal \N__57689\ : std_logic;
signal \N__57686\ : std_logic;
signal \N__57681\ : std_logic;
signal \N__57678\ : std_logic;
signal \N__57677\ : std_logic;
signal \N__57674\ : std_logic;
signal \N__57671\ : std_logic;
signal \N__57668\ : std_logic;
signal \N__57665\ : std_logic;
signal \N__57660\ : std_logic;
signal \N__57657\ : std_logic;
signal \N__57654\ : std_logic;
signal \N__57653\ : std_logic;
signal \N__57650\ : std_logic;
signal \N__57647\ : std_logic;
signal \N__57644\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57636\ : std_logic;
signal \N__57635\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57629\ : std_logic;
signal \N__57626\ : std_logic;
signal \N__57623\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57612\ : std_logic;
signal \N__57609\ : std_logic;
signal \N__57606\ : std_logic;
signal \N__57605\ : std_logic;
signal \N__57602\ : std_logic;
signal \N__57599\ : std_logic;
signal \N__57596\ : std_logic;
signal \N__57591\ : std_logic;
signal \N__57588\ : std_logic;
signal \N__57587\ : std_logic;
signal \N__57584\ : std_logic;
signal \N__57581\ : std_logic;
signal \N__57578\ : std_logic;
signal \N__57575\ : std_logic;
signal \N__57570\ : std_logic;
signal \N__57567\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57563\ : std_logic;
signal \N__57560\ : std_logic;
signal \N__57557\ : std_logic;
signal \N__57554\ : std_logic;
signal \N__57549\ : std_logic;
signal \N__57546\ : std_logic;
signal \N__57543\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57536\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57529\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57519\ : std_logic;
signal \N__57516\ : std_logic;
signal \N__57515\ : std_logic;
signal \N__57512\ : std_logic;
signal \N__57509\ : std_logic;
signal \N__57506\ : std_logic;
signal \N__57503\ : std_logic;
signal \N__57500\ : std_logic;
signal \N__57497\ : std_logic;
signal \N__57492\ : std_logic;
signal \N__57491\ : std_logic;
signal \N__57488\ : std_logic;
signal \N__57485\ : std_logic;
signal \N__57482\ : std_logic;
signal \N__57479\ : std_logic;
signal \N__57474\ : std_logic;
signal \N__57471\ : std_logic;
signal \N__57470\ : std_logic;
signal \N__57467\ : std_logic;
signal \N__57464\ : std_logic;
signal \N__57459\ : std_logic;
signal \N__57456\ : std_logic;
signal \N__57453\ : std_logic;
signal \N__57450\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57441\ : std_logic;
signal \N__57438\ : std_logic;
signal \N__57437\ : std_logic;
signal \N__57434\ : std_logic;
signal \N__57431\ : std_logic;
signal \N__57430\ : std_logic;
signal \N__57425\ : std_logic;
signal \N__57422\ : std_logic;
signal \N__57417\ : std_logic;
signal \N__57414\ : std_logic;
signal \N__57413\ : std_logic;
signal \N__57410\ : std_logic;
signal \N__57407\ : std_logic;
signal \N__57402\ : std_logic;
signal \N__57399\ : std_logic;
signal \N__57396\ : std_logic;
signal \N__57395\ : std_logic;
signal \N__57392\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57386\ : std_logic;
signal \N__57383\ : std_logic;
signal \N__57378\ : std_logic;
signal \N__57375\ : std_logic;
signal \N__57372\ : std_logic;
signal \N__57371\ : std_logic;
signal \N__57368\ : std_logic;
signal \N__57365\ : std_logic;
signal \N__57362\ : std_logic;
signal \N__57359\ : std_logic;
signal \N__57354\ : std_logic;
signal \N__57351\ : std_logic;
signal \N__57348\ : std_logic;
signal \N__57345\ : std_logic;
signal \N__57342\ : std_logic;
signal \N__57339\ : std_logic;
signal \N__57336\ : std_logic;
signal \N__57333\ : std_logic;
signal \N__57330\ : std_logic;
signal \N__57327\ : std_logic;
signal \N__57324\ : std_logic;
signal \N__57321\ : std_logic;
signal \N__57318\ : std_logic;
signal \N__57315\ : std_logic;
signal \N__57312\ : std_logic;
signal \N__57309\ : std_logic;
signal \N__57306\ : std_logic;
signal \N__57303\ : std_logic;
signal \N__57300\ : std_logic;
signal \N__57297\ : std_logic;
signal \N__57294\ : std_logic;
signal \N__57291\ : std_logic;
signal \N__57288\ : std_logic;
signal \N__57285\ : std_logic;
signal \N__57282\ : std_logic;
signal \N__57279\ : std_logic;
signal \N__57276\ : std_logic;
signal \N__57273\ : std_logic;
signal \N__57272\ : std_logic;
signal \N__57271\ : std_logic;
signal \N__57270\ : std_logic;
signal \N__57269\ : std_logic;
signal \N__57268\ : std_logic;
signal \N__57267\ : std_logic;
signal \N__57266\ : std_logic;
signal \N__57265\ : std_logic;
signal \N__57264\ : std_logic;
signal \N__57263\ : std_logic;
signal \N__57262\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57260\ : std_logic;
signal \N__57259\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57257\ : std_logic;
signal \N__57254\ : std_logic;
signal \N__57253\ : std_logic;
signal \N__57252\ : std_logic;
signal \N__57251\ : std_logic;
signal \N__57250\ : std_logic;
signal \N__57249\ : std_logic;
signal \N__57246\ : std_logic;
signal \N__57243\ : std_logic;
signal \N__57240\ : std_logic;
signal \N__57239\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57233\ : std_logic;
signal \N__57230\ : std_logic;
signal \N__57227\ : std_logic;
signal \N__57224\ : std_logic;
signal \N__57221\ : std_logic;
signal \N__57218\ : std_logic;
signal \N__57217\ : std_logic;
signal \N__57214\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57212\ : std_logic;
signal \N__57211\ : std_logic;
signal \N__57210\ : std_logic;
signal \N__57209\ : std_logic;
signal \N__57208\ : std_logic;
signal \N__57207\ : std_logic;
signal \N__57206\ : std_logic;
signal \N__57205\ : std_logic;
signal \N__57204\ : std_logic;
signal \N__57203\ : std_logic;
signal \N__57202\ : std_logic;
signal \N__57199\ : std_logic;
signal \N__57198\ : std_logic;
signal \N__57197\ : std_logic;
signal \N__57196\ : std_logic;
signal \N__57195\ : std_logic;
signal \N__57194\ : std_logic;
signal \N__57191\ : std_logic;
signal \N__57188\ : std_logic;
signal \N__57187\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57185\ : std_logic;
signal \N__57184\ : std_logic;
signal \N__57181\ : std_logic;
signal \N__57180\ : std_logic;
signal \N__57179\ : std_logic;
signal \N__57170\ : std_logic;
signal \N__57167\ : std_logic;
signal \N__57164\ : std_logic;
signal \N__57163\ : std_logic;
signal \N__57162\ : std_logic;
signal \N__57159\ : std_logic;
signal \N__57152\ : std_logic;
signal \N__57151\ : std_logic;
signal \N__57150\ : std_logic;
signal \N__57149\ : std_logic;
signal \N__57148\ : std_logic;
signal \N__57147\ : std_logic;
signal \N__57146\ : std_logic;
signal \N__57143\ : std_logic;
signal \N__57140\ : std_logic;
signal \N__57137\ : std_logic;
signal \N__57136\ : std_logic;
signal \N__57135\ : std_logic;
signal \N__57134\ : std_logic;
signal \N__57133\ : std_logic;
signal \N__57132\ : std_logic;
signal \N__57131\ : std_logic;
signal \N__57130\ : std_logic;
signal \N__57129\ : std_logic;
signal \N__57128\ : std_logic;
signal \N__57127\ : std_logic;
signal \N__57122\ : std_logic;
signal \N__57115\ : std_logic;
signal \N__57114\ : std_logic;
signal \N__57113\ : std_logic;
signal \N__57112\ : std_logic;
signal \N__57111\ : std_logic;
signal \N__57110\ : std_logic;
signal \N__57109\ : std_logic;
signal \N__57106\ : std_logic;
signal \N__57105\ : std_logic;
signal \N__57102\ : std_logic;
signal \N__57101\ : std_logic;
signal \N__57100\ : std_logic;
signal \N__57099\ : std_logic;
signal \N__57098\ : std_logic;
signal \N__57097\ : std_logic;
signal \N__57094\ : std_logic;
signal \N__57093\ : std_logic;
signal \N__57092\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57088\ : std_logic;
signal \N__57083\ : std_logic;
signal \N__57080\ : std_logic;
signal \N__57077\ : std_logic;
signal \N__57072\ : std_logic;
signal \N__57067\ : std_logic;
signal \N__57062\ : std_logic;
signal \N__57059\ : std_logic;
signal \N__57052\ : std_logic;
signal \N__57049\ : std_logic;
signal \N__57046\ : std_logic;
signal \N__57043\ : std_logic;
signal \N__57038\ : std_logic;
signal \N__57035\ : std_logic;
signal \N__57032\ : std_logic;
signal \N__57029\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57027\ : std_logic;
signal \N__57026\ : std_logic;
signal \N__57025\ : std_logic;
signal \N__57024\ : std_logic;
signal \N__57023\ : std_logic;
signal \N__57018\ : std_logic;
signal \N__57015\ : std_logic;
signal \N__57012\ : std_logic;
signal \N__57007\ : std_logic;
signal \N__57004\ : std_logic;
signal \N__56999\ : std_logic;
signal \N__56996\ : std_logic;
signal \N__56993\ : std_logic;
signal \N__56986\ : std_logic;
signal \N__56983\ : std_logic;
signal \N__56980\ : std_logic;
signal \N__56975\ : std_logic;
signal \N__56972\ : std_logic;
signal \N__56961\ : std_logic;
signal \N__56960\ : std_logic;
signal \N__56959\ : std_logic;
signal \N__56958\ : std_logic;
signal \N__56957\ : std_logic;
signal \N__56954\ : std_logic;
signal \N__56949\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56943\ : std_logic;
signal \N__56938\ : std_logic;
signal \N__56937\ : std_logic;
signal \N__56934\ : std_logic;
signal \N__56931\ : std_logic;
signal \N__56928\ : std_logic;
signal \N__56925\ : std_logic;
signal \N__56918\ : std_logic;
signal \N__56915\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56913\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56900\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56898\ : std_logic;
signal \N__56895\ : std_logic;
signal \N__56892\ : std_logic;
signal \N__56889\ : std_logic;
signal \N__56884\ : std_logic;
signal \N__56881\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56874\ : std_logic;
signal \N__56873\ : std_logic;
signal \N__56870\ : std_logic;
signal \N__56869\ : std_logic;
signal \N__56868\ : std_logic;
signal \N__56867\ : std_logic;
signal \N__56866\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56856\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56848\ : std_logic;
signal \N__56843\ : std_logic;
signal \N__56836\ : std_logic;
signal \N__56827\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56807\ : std_logic;
signal \N__56802\ : std_logic;
signal \N__56791\ : std_logic;
signal \N__56788\ : std_logic;
signal \N__56787\ : std_logic;
signal \N__56784\ : std_logic;
signal \N__56783\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56767\ : std_logic;
signal \N__56764\ : std_logic;
signal \N__56753\ : std_logic;
signal \N__56752\ : std_logic;
signal \N__56751\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56738\ : std_logic;
signal \N__56731\ : std_logic;
signal \N__56728\ : std_logic;
signal \N__56723\ : std_logic;
signal \N__56720\ : std_logic;
signal \N__56713\ : std_logic;
signal \N__56710\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56704\ : std_logic;
signal \N__56697\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56687\ : std_logic;
signal \N__56680\ : std_logic;
signal \N__56669\ : std_logic;
signal \N__56660\ : std_logic;
signal \N__56655\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56645\ : std_logic;
signal \N__56628\ : std_logic;
signal \N__56601\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56592\ : std_logic;
signal \N__56589\ : std_logic;
signal \N__56586\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56582\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56575\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56573\ : std_logic;
signal \N__56572\ : std_logic;
signal \N__56571\ : std_logic;
signal \N__56568\ : std_logic;
signal \N__56565\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56557\ : std_logic;
signal \N__56552\ : std_logic;
signal \N__56541\ : std_logic;
signal \N__56538\ : std_logic;
signal \N__56537\ : std_logic;
signal \N__56534\ : std_logic;
signal \N__56531\ : std_logic;
signal \N__56526\ : std_logic;
signal \N__56523\ : std_logic;
signal \N__56520\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56514\ : std_logic;
signal \N__56511\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56505\ : std_logic;
signal \N__56504\ : std_logic;
signal \N__56503\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56497\ : std_logic;
signal \N__56494\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56486\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56477\ : std_logic;
signal \N__56474\ : std_logic;
signal \N__56469\ : std_logic;
signal \N__56466\ : std_logic;
signal \N__56463\ : std_logic;
signal \N__56460\ : std_logic;
signal \N__56457\ : std_logic;
signal \N__56454\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56448\ : std_logic;
signal \N__56447\ : std_logic;
signal \N__56446\ : std_logic;
signal \N__56443\ : std_logic;
signal \N__56438\ : std_logic;
signal \N__56435\ : std_logic;
signal \N__56432\ : std_logic;
signal \N__56429\ : std_logic;
signal \N__56426\ : std_logic;
signal \N__56421\ : std_logic;
signal \N__56418\ : std_logic;
signal \N__56415\ : std_logic;
signal \N__56412\ : std_logic;
signal \N__56409\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56402\ : std_logic;
signal \N__56401\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56391\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56385\ : std_logic;
signal \N__56382\ : std_logic;
signal \N__56381\ : std_logic;
signal \N__56378\ : std_logic;
signal \N__56375\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56369\ : std_logic;
signal \N__56366\ : std_logic;
signal \N__56363\ : std_logic;
signal \N__56358\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56351\ : std_logic;
signal \N__56348\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56340\ : std_logic;
signal \N__56339\ : std_logic;
signal \N__56336\ : std_logic;
signal \N__56333\ : std_logic;
signal \N__56328\ : std_logic;
signal \N__56325\ : std_logic;
signal \N__56322\ : std_logic;
signal \N__56319\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56313\ : std_logic;
signal \N__56310\ : std_logic;
signal \N__56307\ : std_logic;
signal \N__56304\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56298\ : std_logic;
signal \N__56297\ : std_logic;
signal \N__56294\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56288\ : std_logic;
signal \N__56285\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56279\ : std_logic;
signal \N__56276\ : std_logic;
signal \N__56273\ : std_logic;
signal \N__56270\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56264\ : std_logic;
signal \N__56261\ : std_logic;
signal \N__56258\ : std_logic;
signal \N__56255\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56249\ : std_logic;
signal \N__56246\ : std_logic;
signal \N__56243\ : std_logic;
signal \N__56238\ : std_logic;
signal \N__56235\ : std_logic;
signal \N__56232\ : std_logic;
signal \N__56231\ : std_logic;
signal \N__56230\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56222\ : std_logic;
signal \N__56217\ : std_logic;
signal \N__56214\ : std_logic;
signal \N__56205\ : std_logic;
signal \N__56202\ : std_logic;
signal \N__56199\ : std_logic;
signal \N__56198\ : std_logic;
signal \N__56195\ : std_logic;
signal \N__56192\ : std_logic;
signal \N__56187\ : std_logic;
signal \N__56184\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56180\ : std_logic;
signal \N__56177\ : std_logic;
signal \N__56174\ : std_logic;
signal \N__56169\ : std_logic;
signal \N__56168\ : std_logic;
signal \N__56165\ : std_logic;
signal \N__56162\ : std_logic;
signal \N__56159\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56151\ : std_logic;
signal \N__56148\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56141\ : std_logic;
signal \N__56140\ : std_logic;
signal \N__56135\ : std_logic;
signal \N__56132\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56126\ : std_logic;
signal \N__56121\ : std_logic;
signal \N__56118\ : std_logic;
signal \N__56115\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56109\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56102\ : std_logic;
signal \N__56101\ : std_logic;
signal \N__56100\ : std_logic;
signal \N__56099\ : std_logic;
signal \N__56098\ : std_logic;
signal \N__56097\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56095\ : std_logic;
signal \N__56094\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56092\ : std_logic;
signal \N__56091\ : std_logic;
signal \N__56090\ : std_logic;
signal \N__56089\ : std_logic;
signal \N__56088\ : std_logic;
signal \N__56087\ : std_logic;
signal \N__56086\ : std_logic;
signal \N__56085\ : std_logic;
signal \N__56084\ : std_logic;
signal \N__56083\ : std_logic;
signal \N__56082\ : std_logic;
signal \N__56081\ : std_logic;
signal \N__56080\ : std_logic;
signal \N__56079\ : std_logic;
signal \N__56078\ : std_logic;
signal \N__56077\ : std_logic;
signal \N__56076\ : std_logic;
signal \N__56075\ : std_logic;
signal \N__56074\ : std_logic;
signal \N__56073\ : std_logic;
signal \N__56072\ : std_logic;
signal \N__56071\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56068\ : std_logic;
signal \N__56067\ : std_logic;
signal \N__56066\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56064\ : std_logic;
signal \N__56063\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56061\ : std_logic;
signal \N__56060\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56058\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56055\ : std_logic;
signal \N__56054\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56052\ : std_logic;
signal \N__56051\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56049\ : std_logic;
signal \N__56048\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56046\ : std_logic;
signal \N__56045\ : std_logic;
signal \N__56044\ : std_logic;
signal \N__56043\ : std_logic;
signal \N__56042\ : std_logic;
signal \N__56041\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56039\ : std_logic;
signal \N__56038\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56036\ : std_logic;
signal \N__56035\ : std_logic;
signal \N__56034\ : std_logic;
signal \N__56033\ : std_logic;
signal \N__56032\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56028\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56026\ : std_logic;
signal \N__56025\ : std_logic;
signal \N__56024\ : std_logic;
signal \N__56023\ : std_logic;
signal \N__56022\ : std_logic;
signal \N__56021\ : std_logic;
signal \N__56020\ : std_logic;
signal \N__56019\ : std_logic;
signal \N__56018\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56016\ : std_logic;
signal \N__56015\ : std_logic;
signal \N__56014\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56012\ : std_logic;
signal \N__56011\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56009\ : std_logic;
signal \N__56008\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56006\ : std_logic;
signal \N__56005\ : std_logic;
signal \N__56004\ : std_logic;
signal \N__56003\ : std_logic;
signal \N__56002\ : std_logic;
signal \N__56001\ : std_logic;
signal \N__56000\ : std_logic;
signal \N__55999\ : std_logic;
signal \N__55998\ : std_logic;
signal \N__55997\ : std_logic;
signal \N__55996\ : std_logic;
signal \N__55995\ : std_logic;
signal \N__55994\ : std_logic;
signal \N__55993\ : std_logic;
signal \N__55992\ : std_logic;
signal \N__55991\ : std_logic;
signal \N__55990\ : std_logic;
signal \N__55989\ : std_logic;
signal \N__55988\ : std_logic;
signal \N__55987\ : std_logic;
signal \N__55986\ : std_logic;
signal \N__55985\ : std_logic;
signal \N__55984\ : std_logic;
signal \N__55983\ : std_logic;
signal \N__55982\ : std_logic;
signal \N__55981\ : std_logic;
signal \N__55980\ : std_logic;
signal \N__55979\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55977\ : std_logic;
signal \N__55976\ : std_logic;
signal \N__55975\ : std_logic;
signal \N__55974\ : std_logic;
signal \N__55973\ : std_logic;
signal \N__55972\ : std_logic;
signal \N__55971\ : std_logic;
signal \N__55970\ : std_logic;
signal \N__55969\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55967\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55963\ : std_logic;
signal \N__55962\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55958\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55955\ : std_logic;
signal \N__55954\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55952\ : std_logic;
signal \N__55951\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55949\ : std_logic;
signal \N__55948\ : std_logic;
signal \N__55947\ : std_logic;
signal \N__55946\ : std_logic;
signal \N__55945\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55942\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55939\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55937\ : std_logic;
signal \N__55602\ : std_logic;
signal \N__55599\ : std_logic;
signal \N__55596\ : std_logic;
signal \N__55593\ : std_logic;
signal \N__55590\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55581\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55574\ : std_logic;
signal \N__55573\ : std_logic;
signal \N__55572\ : std_logic;
signal \N__55571\ : std_logic;
signal \N__55568\ : std_logic;
signal \N__55565\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55562\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55554\ : std_logic;
signal \N__55553\ : std_logic;
signal \N__55548\ : std_logic;
signal \N__55545\ : std_logic;
signal \N__55544\ : std_logic;
signal \N__55541\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55536\ : std_logic;
signal \N__55533\ : std_logic;
signal \N__55530\ : std_logic;
signal \N__55527\ : std_logic;
signal \N__55524\ : std_logic;
signal \N__55521\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55513\ : std_logic;
signal \N__55508\ : std_logic;
signal \N__55503\ : std_logic;
signal \N__55496\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55482\ : std_logic;
signal \N__55479\ : std_logic;
signal \N__55478\ : std_logic;
signal \N__55475\ : std_logic;
signal \N__55474\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55472\ : std_logic;
signal \N__55471\ : std_logic;
signal \N__55470\ : std_logic;
signal \N__55469\ : std_logic;
signal \N__55468\ : std_logic;
signal \N__55467\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55464\ : std_logic;
signal \N__55463\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55461\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55456\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55441\ : std_logic;
signal \N__55440\ : std_logic;
signal \N__55439\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55437\ : std_logic;
signal \N__55436\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55434\ : std_logic;
signal \N__55433\ : std_logic;
signal \N__55432\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55429\ : std_logic;
signal \N__55428\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55424\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55422\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55419\ : std_logic;
signal \N__55418\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55414\ : std_logic;
signal \N__55411\ : std_logic;
signal \N__55410\ : std_logic;
signal \N__55407\ : std_logic;
signal \N__55406\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55402\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55388\ : std_logic;
signal \N__55387\ : std_logic;
signal \N__55384\ : std_logic;
signal \N__55381\ : std_logic;
signal \N__55378\ : std_logic;
signal \N__55373\ : std_logic;
signal \N__55368\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55358\ : std_logic;
signal \N__55355\ : std_logic;
signal \N__55352\ : std_logic;
signal \N__55347\ : std_logic;
signal \N__55346\ : std_logic;
signal \N__55343\ : std_logic;
signal \N__55336\ : std_logic;
signal \N__55325\ : std_logic;
signal \N__55322\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55302\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55298\ : std_logic;
signal \N__55297\ : std_logic;
signal \N__55296\ : std_logic;
signal \N__55295\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55293\ : std_logic;
signal \N__55292\ : std_logic;
signal \N__55289\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55287\ : std_logic;
signal \N__55286\ : std_logic;
signal \N__55285\ : std_logic;
signal \N__55282\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55280\ : std_logic;
signal \N__55279\ : std_logic;
signal \N__55276\ : std_logic;
signal \N__55273\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55271\ : std_logic;
signal \N__55270\ : std_logic;
signal \N__55269\ : std_logic;
signal \N__55268\ : std_logic;
signal \N__55255\ : std_logic;
signal \N__55252\ : std_logic;
signal \N__55251\ : std_logic;
signal \N__55250\ : std_logic;
signal \N__55249\ : std_logic;
signal \N__55248\ : std_logic;
signal \N__55247\ : std_logic;
signal \N__55244\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55238\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55236\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55233\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55227\ : std_logic;
signal \N__55216\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55208\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55204\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55181\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55171\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55144\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55136\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55108\ : std_logic;
signal \N__55105\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55096\ : std_logic;
signal \N__55091\ : std_logic;
signal \N__55088\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55069\ : std_logic;
signal \N__55068\ : std_logic;
signal \N__55067\ : std_logic;
signal \N__55066\ : std_logic;
signal \N__55065\ : std_logic;
signal \N__55062\ : std_logic;
signal \N__55059\ : std_logic;
signal \N__55056\ : std_logic;
signal \N__55051\ : std_logic;
signal \N__55044\ : std_logic;
signal \N__55033\ : std_logic;
signal \N__55030\ : std_logic;
signal \N__55029\ : std_logic;
signal \N__55028\ : std_logic;
signal \N__55027\ : std_logic;
signal \N__55024\ : std_logic;
signal \N__55017\ : std_logic;
signal \N__55014\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55008\ : std_logic;
signal \N__55005\ : std_logic;
signal \N__55002\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54990\ : std_logic;
signal \N__54985\ : std_logic;
signal \N__54980\ : std_logic;
signal \N__54977\ : std_logic;
signal \N__54974\ : std_logic;
signal \N__54965\ : std_logic;
signal \N__54958\ : std_logic;
signal \N__54951\ : std_logic;
signal \N__54946\ : std_logic;
signal \N__54941\ : std_logic;
signal \N__54934\ : std_logic;
signal \N__54931\ : std_logic;
signal \N__54924\ : std_logic;
signal \N__54903\ : std_logic;
signal \N__54900\ : std_logic;
signal \N__54897\ : std_logic;
signal \N__54894\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54892\ : std_logic;
signal \N__54891\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54887\ : std_logic;
signal \N__54886\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54884\ : std_logic;
signal \N__54881\ : std_logic;
signal \N__54876\ : std_logic;
signal \N__54875\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54864\ : std_logic;
signal \N__54863\ : std_logic;
signal \N__54862\ : std_logic;
signal \N__54861\ : std_logic;
signal \N__54860\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54858\ : std_logic;
signal \N__54857\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54853\ : std_logic;
signal \N__54852\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54848\ : std_logic;
signal \N__54847\ : std_logic;
signal \N__54844\ : std_logic;
signal \N__54843\ : std_logic;
signal \N__54842\ : std_logic;
signal \N__54841\ : std_logic;
signal \N__54840\ : std_logic;
signal \N__54839\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54828\ : std_logic;
signal \N__54827\ : std_logic;
signal \N__54826\ : std_logic;
signal \N__54825\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54811\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54804\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54800\ : std_logic;
signal \N__54797\ : std_logic;
signal \N__54796\ : std_logic;
signal \N__54795\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54788\ : std_logic;
signal \N__54787\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54781\ : std_logic;
signal \N__54778\ : std_logic;
signal \N__54777\ : std_logic;
signal \N__54774\ : std_logic;
signal \N__54771\ : std_logic;
signal \N__54766\ : std_logic;
signal \N__54761\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54755\ : std_logic;
signal \N__54754\ : std_logic;
signal \N__54753\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54741\ : std_logic;
signal \N__54740\ : std_logic;
signal \N__54739\ : std_logic;
signal \N__54738\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54734\ : std_logic;
signal \N__54731\ : std_logic;
signal \N__54728\ : std_logic;
signal \N__54725\ : std_logic;
signal \N__54716\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54707\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54696\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54685\ : std_logic;
signal \N__54684\ : std_logic;
signal \N__54683\ : std_logic;
signal \N__54680\ : std_logic;
signal \N__54675\ : std_logic;
signal \N__54670\ : std_logic;
signal \N__54667\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54652\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54646\ : std_logic;
signal \N__54643\ : std_logic;
signal \N__54640\ : std_logic;
signal \N__54633\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54594\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54572\ : std_logic;
signal \N__54571\ : std_logic;
signal \N__54568\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54566\ : std_logic;
signal \N__54563\ : std_logic;
signal \N__54560\ : std_logic;
signal \N__54557\ : std_logic;
signal \N__54556\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54554\ : std_logic;
signal \N__54553\ : std_logic;
signal \N__54552\ : std_logic;
signal \N__54551\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54549\ : std_logic;
signal \N__54548\ : std_logic;
signal \N__54547\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54545\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54542\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54526\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54515\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54503\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54500\ : std_logic;
signal \N__54499\ : std_logic;
signal \N__54498\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54491\ : std_logic;
signal \N__54490\ : std_logic;
signal \N__54489\ : std_logic;
signal \N__54488\ : std_logic;
signal \N__54487\ : std_logic;
signal \N__54486\ : std_logic;
signal \N__54485\ : std_logic;
signal \N__54484\ : std_logic;
signal \N__54467\ : std_logic;
signal \N__54464\ : std_logic;
signal \N__54461\ : std_logic;
signal \N__54458\ : std_logic;
signal \N__54455\ : std_logic;
signal \N__54452\ : std_logic;
signal \N__54449\ : std_logic;
signal \N__54444\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54440\ : std_logic;
signal \N__54439\ : std_logic;
signal \N__54438\ : std_logic;
signal \N__54437\ : std_logic;
signal \N__54436\ : std_logic;
signal \N__54435\ : std_logic;
signal \N__54434\ : std_logic;
signal \N__54433\ : std_logic;
signal \N__54432\ : std_logic;
signal \N__54431\ : std_logic;
signal \N__54430\ : std_logic;
signal \N__54429\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54418\ : std_logic;
signal \N__54417\ : std_logic;
signal \N__54414\ : std_logic;
signal \N__54411\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54409\ : std_logic;
signal \N__54406\ : std_logic;
signal \N__54403\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54401\ : std_logic;
signal \N__54400\ : std_logic;
signal \N__54397\ : std_logic;
signal \N__54390\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54380\ : std_logic;
signal \N__54379\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54375\ : std_logic;
signal \N__54374\ : std_logic;
signal \N__54371\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54366\ : std_logic;
signal \N__54363\ : std_logic;
signal \N__54360\ : std_logic;
signal \N__54357\ : std_logic;
signal \N__54350\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54340\ : std_logic;
signal \N__54339\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54333\ : std_logic;
signal \N__54332\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54326\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54308\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54300\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54276\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__54266\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54256\ : std_logic;
signal \N__54251\ : std_logic;
signal \N__54248\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54242\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54232\ : std_logic;
signal \N__54225\ : std_logic;
signal \N__54222\ : std_logic;
signal \N__54217\ : std_logic;
signal \N__54212\ : std_logic;
signal \N__54201\ : std_logic;
signal \N__54200\ : std_logic;
signal \N__54199\ : std_logic;
signal \N__54198\ : std_logic;
signal \N__54197\ : std_logic;
signal \N__54196\ : std_logic;
signal \N__54195\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54193\ : std_logic;
signal \N__54192\ : std_logic;
signal \N__54191\ : std_logic;
signal \N__54188\ : std_logic;
signal \N__54185\ : std_logic;
signal \N__54184\ : std_logic;
signal \N__54183\ : std_logic;
signal \N__54180\ : std_logic;
signal \N__54179\ : std_logic;
signal \N__54178\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54174\ : std_logic;
signal \N__54173\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54155\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54141\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54129\ : std_logic;
signal \N__54126\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54078\ : std_logic;
signal \N__54075\ : std_logic;
signal \N__54068\ : std_logic;
signal \N__54063\ : std_logic;
signal \N__54054\ : std_logic;
signal \N__54047\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54037\ : std_logic;
signal \N__54032\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54008\ : std_logic;
signal \N__54007\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__54004\ : std_logic;
signal \N__54003\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53989\ : std_logic;
signal \N__53988\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53981\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53965\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53959\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53951\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53946\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53924\ : std_logic;
signal \N__53923\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53921\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53916\ : std_logic;
signal \N__53913\ : std_logic;
signal \N__53910\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53900\ : std_logic;
signal \N__53897\ : std_logic;
signal \N__53894\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53883\ : std_logic;
signal \N__53880\ : std_logic;
signal \N__53877\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53873\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53870\ : std_logic;
signal \N__53869\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53860\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53850\ : std_logic;
signal \N__53845\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53833\ : std_logic;
signal \N__53830\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53820\ : std_logic;
signal \N__53811\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53790\ : std_logic;
signal \N__53775\ : std_logic;
signal \N__53772\ : std_logic;
signal \N__53769\ : std_logic;
signal \N__53766\ : std_logic;
signal \N__53763\ : std_logic;
signal \N__53760\ : std_logic;
signal \N__53757\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53747\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53738\ : std_logic;
signal \N__53735\ : std_logic;
signal \N__53732\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53726\ : std_logic;
signal \N__53723\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53712\ : std_logic;
signal \N__53711\ : std_logic;
signal \N__53708\ : std_logic;
signal \N__53705\ : std_logic;
signal \N__53702\ : std_logic;
signal \N__53697\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53688\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53675\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53671\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53663\ : std_logic;
signal \N__53660\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53652\ : std_logic;
signal \N__53649\ : std_logic;
signal \N__53646\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53644\ : std_logic;
signal \N__53641\ : std_logic;
signal \N__53640\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53636\ : std_logic;
signal \N__53633\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53627\ : std_logic;
signal \N__53624\ : std_logic;
signal \N__53621\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53619\ : std_logic;
signal \N__53612\ : std_logic;
signal \N__53607\ : std_logic;
signal \N__53604\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53600\ : std_logic;
signal \N__53597\ : std_logic;
signal \N__53594\ : std_logic;
signal \N__53591\ : std_logic;
signal \N__53588\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53584\ : std_logic;
signal \N__53581\ : std_logic;
signal \N__53578\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53570\ : std_logic;
signal \N__53567\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53553\ : std_logic;
signal \N__53552\ : std_logic;
signal \N__53549\ : std_logic;
signal \N__53546\ : std_logic;
signal \N__53543\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53535\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53520\ : std_logic;
signal \N__53517\ : std_logic;
signal \N__53514\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53507\ : std_logic;
signal \N__53504\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53499\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53487\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53477\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53471\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53462\ : std_logic;
signal \N__53459\ : std_logic;
signal \N__53458\ : std_logic;
signal \N__53455\ : std_logic;
signal \N__53452\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53435\ : std_logic;
signal \N__53432\ : std_logic;
signal \N__53425\ : std_logic;
signal \N__53424\ : std_logic;
signal \N__53423\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53415\ : std_logic;
signal \N__53412\ : std_logic;
signal \N__53407\ : std_logic;
signal \N__53404\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53398\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53384\ : std_logic;
signal \N__53381\ : std_logic;
signal \N__53378\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53370\ : std_logic;
signal \N__53367\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53355\ : std_logic;
signal \N__53352\ : std_logic;
signal \N__53349\ : std_logic;
signal \N__53346\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53344\ : std_logic;
signal \N__53343\ : std_logic;
signal \N__53342\ : std_logic;
signal \N__53339\ : std_logic;
signal \N__53336\ : std_logic;
signal \N__53333\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53328\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53322\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53313\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53305\ : std_logic;
signal \N__53298\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53292\ : std_logic;
signal \N__53291\ : std_logic;
signal \N__53288\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53280\ : std_logic;
signal \N__53277\ : std_logic;
signal \N__53268\ : std_logic;
signal \N__53267\ : std_logic;
signal \N__53264\ : std_logic;
signal \N__53261\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53235\ : std_logic;
signal \N__53234\ : std_logic;
signal \N__53231\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53227\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53218\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53208\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53202\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53192\ : std_logic;
signal \N__53189\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53177\ : std_logic;
signal \N__53174\ : std_logic;
signal \N__53171\ : std_logic;
signal \N__53166\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53157\ : std_logic;
signal \N__53152\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53141\ : std_logic;
signal \N__53138\ : std_logic;
signal \N__53135\ : std_logic;
signal \N__53132\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53129\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53126\ : std_logic;
signal \N__53123\ : std_logic;
signal \N__53120\ : std_logic;
signal \N__53117\ : std_logic;
signal \N__53114\ : std_logic;
signal \N__53109\ : std_logic;
signal \N__53106\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53084\ : std_logic;
signal \N__53081\ : std_logic;
signal \N__53078\ : std_logic;
signal \N__53073\ : std_logic;
signal \N__53072\ : std_logic;
signal \N__53071\ : std_logic;
signal \N__53070\ : std_logic;
signal \N__53069\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53066\ : std_logic;
signal \N__53065\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53063\ : std_logic;
signal \N__53062\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53051\ : std_logic;
signal \N__53050\ : std_logic;
signal \N__53049\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53047\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53042\ : std_logic;
signal \N__53037\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53033\ : std_logic;
signal \N__53032\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53030\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52992\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52988\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52986\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52980\ : std_logic;
signal \N__52975\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52951\ : std_logic;
signal \N__52948\ : std_logic;
signal \N__52939\ : std_logic;
signal \N__52938\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52920\ : std_logic;
signal \N__52915\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52890\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52884\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52881\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52869\ : std_logic;
signal \N__52864\ : std_logic;
signal \N__52863\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52859\ : std_logic;
signal \N__52858\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52856\ : std_logic;
signal \N__52855\ : std_logic;
signal \N__52852\ : std_logic;
signal \N__52849\ : std_logic;
signal \N__52846\ : std_logic;
signal \N__52839\ : std_logic;
signal \N__52828\ : std_logic;
signal \N__52825\ : std_logic;
signal \N__52820\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52803\ : std_logic;
signal \N__52800\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52798\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52796\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52784\ : std_logic;
signal \N__52783\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52778\ : std_logic;
signal \N__52775\ : std_logic;
signal \N__52772\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52767\ : std_logic;
signal \N__52764\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52756\ : std_logic;
signal \N__52753\ : std_logic;
signal \N__52750\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52724\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52712\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52698\ : std_logic;
signal \N__52695\ : std_logic;
signal \N__52692\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52690\ : std_logic;
signal \N__52685\ : std_logic;
signal \N__52682\ : std_logic;
signal \N__52679\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52661\ : std_logic;
signal \N__52658\ : std_logic;
signal \N__52653\ : std_logic;
signal \N__52650\ : std_logic;
signal \N__52647\ : std_logic;
signal \N__52644\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52628\ : std_logic;
signal \N__52625\ : std_logic;
signal \N__52622\ : std_logic;
signal \N__52619\ : std_logic;
signal \N__52616\ : std_logic;
signal \N__52613\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52607\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52596\ : std_logic;
signal \N__52593\ : std_logic;
signal \N__52590\ : std_logic;
signal \N__52587\ : std_logic;
signal \N__52584\ : std_logic;
signal \N__52581\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52575\ : std_logic;
signal \N__52572\ : std_logic;
signal \N__52569\ : std_logic;
signal \N__52566\ : std_logic;
signal \N__52565\ : std_logic;
signal \N__52564\ : std_logic;
signal \N__52563\ : std_logic;
signal \N__52562\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52560\ : std_logic;
signal \N__52559\ : std_logic;
signal \N__52558\ : std_logic;
signal \N__52557\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52555\ : std_logic;
signal \N__52554\ : std_logic;
signal \N__52553\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52532\ : std_logic;
signal \N__52527\ : std_logic;
signal \N__52524\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52521\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52517\ : std_logic;
signal \N__52514\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52490\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52460\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52448\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52436\ : std_logic;
signal \N__52435\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52433\ : std_logic;
signal \N__52432\ : std_logic;
signal \N__52429\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52423\ : std_logic;
signal \N__52420\ : std_logic;
signal \N__52415\ : std_logic;
signal \N__52412\ : std_logic;
signal \N__52411\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52409\ : std_logic;
signal \N__52406\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52394\ : std_logic;
signal \N__52393\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52382\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52377\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52355\ : std_logic;
signal \N__52350\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52340\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52334\ : std_logic;
signal \N__52325\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52299\ : std_logic;
signal \N__52290\ : std_logic;
signal \N__52287\ : std_logic;
signal \N__52286\ : std_logic;
signal \N__52285\ : std_logic;
signal \N__52282\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52278\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52275\ : std_logic;
signal \N__52272\ : std_logic;
signal \N__52269\ : std_logic;
signal \N__52266\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52260\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52225\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52209\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52197\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52169\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52163\ : std_logic;
signal \N__52160\ : std_logic;
signal \N__52157\ : std_logic;
signal \N__52152\ : std_logic;
signal \N__52151\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52144\ : std_logic;
signal \N__52141\ : std_logic;
signal \N__52138\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52129\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52101\ : std_logic;
signal \N__52098\ : std_logic;
signal \N__52095\ : std_logic;
signal \N__52094\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52075\ : std_logic;
signal \N__52072\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52064\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52056\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52052\ : std_logic;
signal \N__52049\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52041\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52035\ : std_logic;
signal \N__52032\ : std_logic;
signal \N__52029\ : std_logic;
signal \N__52026\ : std_logic;
signal \N__52023\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52014\ : std_logic;
signal \N__52011\ : std_logic;
signal \N__52008\ : std_logic;
signal \N__52005\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__52000\ : std_logic;
signal \N__51997\ : std_logic;
signal \N__51994\ : std_logic;
signal \N__51993\ : std_logic;
signal \N__51990\ : std_logic;
signal \N__51987\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51982\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51959\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51948\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51939\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51918\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51912\ : std_logic;
signal \N__51911\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51909\ : std_logic;
signal \N__51908\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51897\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51889\ : std_logic;
signal \N__51886\ : std_logic;
signal \N__51883\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51880\ : std_logic;
signal \N__51877\ : std_logic;
signal \N__51874\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51864\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51858\ : std_logic;
signal \N__51857\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51833\ : std_logic;
signal \N__51828\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51820\ : std_logic;
signal \N__51817\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51811\ : std_logic;
signal \N__51806\ : std_logic;
signal \N__51803\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51789\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51762\ : std_logic;
signal \N__51761\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51759\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51754\ : std_logic;
signal \N__51753\ : std_logic;
signal \N__51750\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51746\ : std_logic;
signal \N__51745\ : std_logic;
signal \N__51744\ : std_logic;
signal \N__51741\ : std_logic;
signal \N__51738\ : std_logic;
signal \N__51735\ : std_logic;
signal \N__51732\ : std_logic;
signal \N__51729\ : std_logic;
signal \N__51726\ : std_logic;
signal \N__51723\ : std_logic;
signal \N__51722\ : std_logic;
signal \N__51721\ : std_logic;
signal \N__51720\ : std_logic;
signal \N__51717\ : std_logic;
signal \N__51714\ : std_logic;
signal \N__51713\ : std_logic;
signal \N__51712\ : std_logic;
signal \N__51711\ : std_logic;
signal \N__51710\ : std_logic;
signal \N__51709\ : std_logic;
signal \N__51708\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51706\ : std_logic;
signal \N__51705\ : std_logic;
signal \N__51704\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51701\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51699\ : std_logic;
signal \N__51698\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51696\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51690\ : std_logic;
signal \N__51687\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51661\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51648\ : std_logic;
signal \N__51645\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51641\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51636\ : std_logic;
signal \N__51635\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51625\ : std_logic;
signal \N__51616\ : std_logic;
signal \N__51609\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51603\ : std_logic;
signal \N__51602\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51600\ : std_logic;
signal \N__51599\ : std_logic;
signal \N__51596\ : std_logic;
signal \N__51593\ : std_logic;
signal \N__51590\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51575\ : std_logic;
signal \N__51560\ : std_logic;
signal \N__51557\ : std_logic;
signal \N__51550\ : std_logic;
signal \N__51539\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51521\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51501\ : std_logic;
signal \N__51500\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51497\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51494\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51491\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51489\ : std_logic;
signal \N__51488\ : std_logic;
signal \N__51485\ : std_logic;
signal \N__51484\ : std_logic;
signal \N__51483\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51481\ : std_logic;
signal \N__51480\ : std_logic;
signal \N__51479\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51475\ : std_logic;
signal \N__51474\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51456\ : std_logic;
signal \N__51455\ : std_logic;
signal \N__51452\ : std_logic;
signal \N__51449\ : std_logic;
signal \N__51446\ : std_logic;
signal \N__51443\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51437\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51416\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51413\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51385\ : std_logic;
signal \N__51380\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51371\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51363\ : std_logic;
signal \N__51362\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51357\ : std_logic;
signal \N__51356\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51345\ : std_logic;
signal \N__51344\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51332\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51329\ : std_logic;
signal \N__51328\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51295\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51281\ : std_logic;
signal \N__51278\ : std_logic;
signal \N__51275\ : std_logic;
signal \N__51272\ : std_logic;
signal \N__51269\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51257\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51246\ : std_logic;
signal \N__51237\ : std_logic;
signal \N__51216\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51212\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51209\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51188\ : std_logic;
signal \N__51185\ : std_logic;
signal \N__51184\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51179\ : std_logic;
signal \N__51176\ : std_logic;
signal \N__51175\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51158\ : std_logic;
signal \N__51155\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51152\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51149\ : std_logic;
signal \N__51146\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51133\ : std_logic;
signal \N__51130\ : std_logic;
signal \N__51125\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51072\ : std_logic;
signal \N__51069\ : std_logic;
signal \N__51066\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51060\ : std_logic;
signal \N__51057\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51051\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51030\ : std_logic;
signal \N__51027\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51021\ : std_logic;
signal \N__51020\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51012\ : std_logic;
signal \N__51009\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51005\ : std_logic;
signal \N__51002\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50991\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50982\ : std_logic;
signal \N__50981\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50972\ : std_logic;
signal \N__50969\ : std_logic;
signal \N__50966\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50941\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50928\ : std_logic;
signal \N__50925\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50905\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50892\ : std_logic;
signal \N__50891\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50879\ : std_logic;
signal \N__50876\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50870\ : std_logic;
signal \N__50869\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50863\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50846\ : std_logic;
signal \N__50843\ : std_logic;
signal \N__50840\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50832\ : std_logic;
signal \N__50829\ : std_logic;
signal \N__50826\ : std_logic;
signal \N__50823\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50807\ : std_logic;
signal \N__50804\ : std_logic;
signal \N__50803\ : std_logic;
signal \N__50800\ : std_logic;
signal \N__50799\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50796\ : std_logic;
signal \N__50795\ : std_logic;
signal \N__50794\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50792\ : std_logic;
signal \N__50791\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50789\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50786\ : std_logic;
signal \N__50785\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50783\ : std_logic;
signal \N__50782\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50729\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50720\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50691\ : std_logic;
signal \N__50688\ : std_logic;
signal \N__50685\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50679\ : std_logic;
signal \N__50676\ : std_logic;
signal \N__50673\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50664\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50654\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50644\ : std_logic;
signal \N__50641\ : std_logic;
signal \N__50638\ : std_logic;
signal \N__50635\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50607\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50600\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50583\ : std_logic;
signal \N__50580\ : std_logic;
signal \N__50577\ : std_logic;
signal \N__50574\ : std_logic;
signal \N__50571\ : std_logic;
signal \N__50568\ : std_logic;
signal \N__50567\ : std_logic;
signal \N__50564\ : std_logic;
signal \N__50561\ : std_logic;
signal \N__50556\ : std_logic;
signal \N__50553\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50549\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50535\ : std_logic;
signal \N__50534\ : std_logic;
signal \N__50531\ : std_logic;
signal \N__50528\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50505\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50447\ : std_logic;
signal \N__50442\ : std_logic;
signal \N__50439\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50433\ : std_logic;
signal \N__50430\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50423\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50414\ : std_logic;
signal \N__50411\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50385\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50364\ : std_logic;
signal \N__50361\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50343\ : std_logic;
signal \N__50342\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50333\ : std_logic;
signal \N__50330\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50321\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50305\ : std_logic;
signal \N__50302\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50291\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50261\ : std_logic;
signal \N__50258\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50250\ : std_logic;
signal \N__50247\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50243\ : std_logic;
signal \N__50240\ : std_logic;
signal \N__50237\ : std_logic;
signal \N__50232\ : std_logic;
signal \N__50231\ : std_logic;
signal \N__50228\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50216\ : std_logic;
signal \N__50213\ : std_logic;
signal \N__50210\ : std_logic;
signal \N__50207\ : std_logic;
signal \N__50204\ : std_logic;
signal \N__50201\ : std_logic;
signal \N__50198\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50156\ : std_logic;
signal \N__50153\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50125\ : std_logic;
signal \N__50122\ : std_logic;
signal \N__50119\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50108\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50085\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50072\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50066\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50034\ : std_logic;
signal \N__50031\ : std_logic;
signal \N__50028\ : std_logic;
signal \N__50025\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49993\ : std_logic;
signal \N__49988\ : std_logic;
signal \N__49985\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49970\ : std_logic;
signal \N__49967\ : std_logic;
signal \N__49964\ : std_logic;
signal \N__49959\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49749\ : std_logic;
signal \N__49746\ : std_logic;
signal \N__49745\ : std_logic;
signal \N__49742\ : std_logic;
signal \N__49739\ : std_logic;
signal \N__49736\ : std_logic;
signal \N__49733\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49724\ : std_logic;
signal \N__49723\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49721\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49717\ : std_logic;
signal \N__49714\ : std_logic;
signal \N__49711\ : std_logic;
signal \N__49708\ : std_logic;
signal \N__49705\ : std_logic;
signal \N__49704\ : std_logic;
signal \N__49701\ : std_logic;
signal \N__49698\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49679\ : std_logic;
signal \N__49678\ : std_logic;
signal \N__49675\ : std_logic;
signal \N__49672\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49659\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49649\ : std_logic;
signal \N__49644\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49623\ : std_logic;
signal \N__49620\ : std_logic;
signal \N__49617\ : std_logic;
signal \N__49614\ : std_logic;
signal \N__49611\ : std_logic;
signal \N__49608\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49586\ : std_logic;
signal \N__49585\ : std_logic;
signal \N__49582\ : std_logic;
signal \N__49579\ : std_logic;
signal \N__49576\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49568\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49541\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49505\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49496\ : std_logic;
signal \N__49495\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49491\ : std_logic;
signal \N__49488\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49483\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49465\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49376\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49310\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__49284\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49273\ : std_logic;
signal \N__49272\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49258\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49235\ : std_logic;
signal \N__49234\ : std_logic;
signal \N__49231\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49214\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49204\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49151\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49133\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49127\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49112\ : std_logic;
signal \N__49109\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49062\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49043\ : std_logic;
signal \N__49030\ : std_logic;
signal \N__49021\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48992\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48956\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48946\ : std_logic;
signal \N__48943\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48876\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48697\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48690\ : std_logic;
signal \N__48687\ : std_logic;
signal \N__48684\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48676\ : std_logic;
signal \N__48673\ : std_logic;
signal \N__48668\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48650\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48615\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48606\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48598\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48595\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48589\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48579\ : std_logic;
signal \N__48576\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48560\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48543\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48444\ : std_logic;
signal \N__48441\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48423\ : std_logic;
signal \N__48420\ : std_logic;
signal \N__48417\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48407\ : std_logic;
signal \N__48404\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48398\ : std_logic;
signal \N__48395\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48363\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48273\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48072\ : std_logic;
signal \N__48069\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48063\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48054\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48030\ : std_logic;
signal \N__48027\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48015\ : std_logic;
signal \N__48012\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__48000\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47976\ : std_logic;
signal \N__47973\ : std_logic;
signal \N__47970\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47946\ : std_logic;
signal \N__47943\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47923\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47920\ : std_logic;
signal \N__47917\ : std_logic;
signal \N__47916\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47910\ : std_logic;
signal \N__47909\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47906\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47896\ : std_logic;
signal \N__47893\ : std_logic;
signal \N__47890\ : std_logic;
signal \N__47887\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47760\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47723\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47712\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47709\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47692\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47679\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47675\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47672\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47668\ : std_logic;
signal \N__47667\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47663\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47625\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47560\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47397\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47270\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47251\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47227\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47215\ : std_logic;
signal \N__47212\ : std_logic;
signal \N__47209\ : std_logic;
signal \N__47204\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47194\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47191\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47133\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47131\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46954\ : std_logic;
signal \N__46951\ : std_logic;
signal \N__46948\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46931\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46925\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46906\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46894\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46890\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46886\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46873\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46859\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46847\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46836\ : std_logic;
signal \N__46833\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46801\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46784\ : std_logic;
signal \N__46781\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46766\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46755\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46745\ : std_logic;
signal \N__46742\ : std_logic;
signal \N__46739\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46729\ : std_logic;
signal \N__46726\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46673\ : std_logic;
signal \N__46670\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46617\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46571\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46551\ : std_logic;
signal \N__46548\ : std_logic;
signal \N__46545\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46505\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46478\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46472\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46445\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46403\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46397\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46324\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46291\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46244\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46197\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46178\ : std_logic;
signal \N__46175\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46072\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46036\ : std_logic;
signal \N__46033\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46024\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45936\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45918\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45878\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45821\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45806\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45791\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45729\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45690\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45420\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45399\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45363\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45348\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45339\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45335\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45290\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45269\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45237\ : std_logic;
signal \N__45234\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45171\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45151\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45145\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45063\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45017\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45008\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44986\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44970\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44959\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44904\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44856\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44841\ : std_logic;
signal \N__44838\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44816\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44810\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44791\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44775\ : std_logic;
signal \N__44772\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44753\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44708\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44702\ : std_logic;
signal \N__44699\ : std_logic;
signal \N__44696\ : std_logic;
signal \N__44693\ : std_logic;
signal \N__44690\ : std_logic;
signal \N__44687\ : std_logic;
signal \N__44684\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44668\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44645\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44633\ : std_logic;
signal \N__44630\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44627\ : std_logic;
signal \N__44626\ : std_logic;
signal \N__44623\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44579\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44512\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44504\ : std_logic;
signal \N__44503\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44456\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44453\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44450\ : std_logic;
signal \N__44449\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44444\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44385\ : std_logic;
signal \N__44380\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44324\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44312\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44280\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44078\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44051\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44037\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44002\ : std_logic;
signal \N__44001\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43992\ : std_logic;
signal \N__43989\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43926\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43900\ : std_logic;
signal \N__43897\ : std_logic;
signal \N__43894\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43862\ : std_logic;
signal \N__43859\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43812\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43785\ : std_logic;
signal \N__43782\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43745\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43741\ : std_logic;
signal \N__43738\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43697\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43636\ : std_logic;
signal \N__43633\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43617\ : std_logic;
signal \N__43614\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43610\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43602\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43595\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43538\ : std_logic;
signal \N__43535\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43482\ : std_logic;
signal \N__43479\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43433\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43318\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43309\ : std_logic;
signal \N__43306\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43286\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43271\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43106\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43100\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43072\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43064\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43025\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43015\ : std_logic;
signal \N__43012\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43002\ : std_logic;
signal \N__42999\ : std_logic;
signal \N__42996\ : std_logic;
signal \N__42995\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42938\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42891\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42887\ : std_logic;
signal \N__42884\ : std_logic;
signal \N__42881\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42877\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42871\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42857\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42847\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42775\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42744\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42683\ : std_logic;
signal \N__42680\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42639\ : std_logic;
signal \N__42636\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42627\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42542\ : std_logic;
signal \N__42539\ : std_logic;
signal \N__42536\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42517\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42480\ : std_logic;
signal \N__42477\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42443\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42430\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42425\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42410\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42403\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42395\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42383\ : std_logic;
signal \N__42380\ : std_logic;
signal \N__42377\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42365\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42335\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42320\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42302\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42286\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42276\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42218\ : std_logic;
signal \N__42215\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42131\ : std_logic;
signal \N__42128\ : std_logic;
signal \N__42125\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42083\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42032\ : std_logic;
signal \N__42029\ : std_logic;
signal \N__42026\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41974\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41963\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41900\ : std_logic;
signal \N__41897\ : std_logic;
signal \N__41894\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41843\ : std_logic;
signal \N__41840\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41831\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41810\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41804\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41780\ : std_logic;
signal \N__41777\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41742\ : std_logic;
signal \N__41739\ : std_logic;
signal \N__41736\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41701\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41683\ : std_logic;
signal \N__41680\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41666\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41663\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41644\ : std_logic;
signal \N__41641\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41599\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41568\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41530\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41508\ : std_logic;
signal \N__41505\ : std_logic;
signal \N__41502\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41498\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41455\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41435\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41411\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41373\ : std_logic;
signal \N__41370\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41297\ : std_logic;
signal \N__41296\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41237\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41219\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41049\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41019\ : std_logic;
signal \N__41016\ : std_logic;
signal \N__41013\ : std_logic;
signal \N__41010\ : std_logic;
signal \N__41007\ : std_logic;
signal \N__41004\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40897\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40812\ : std_logic;
signal \N__40809\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40719\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40707\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40688\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40550\ : std_logic;
signal \N__40547\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40516\ : std_logic;
signal \N__40505\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40427\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40379\ : std_logic;
signal \N__40376\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40343\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40328\ : std_logic;
signal \N__40327\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40322\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40307\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40172\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40148\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40124\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40103\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40055\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40046\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39998\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39938\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39854\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39839\ : std_logic;
signal \N__39836\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39731\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39722\ : std_logic;
signal \N__39719\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39641\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39586\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39515\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39503\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39435\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39266\ : std_logic;
signal \N__39263\ : std_logic;
signal \N__39260\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39242\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39230\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39188\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39170\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39136\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39127\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39118\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39100\ : std_logic;
signal \N__39097\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39070\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38972\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38944\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38847\ : std_logic;
signal \N__38844\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38745\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38579\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38563\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38552\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38507\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38447\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38415\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38404\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38401\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38398\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38150\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38096\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38045\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38033\ : std_logic;
signal \N__38030\ : std_logic;
signal \N__38027\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37856\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37850\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37821\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37802\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37667\ : std_logic;
signal \N__37664\ : std_logic;
signal \N__37661\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37572\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37295\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37276\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37079\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37043\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36998\ : std_logic;
signal \N__36995\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36740\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36726\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36533\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36522\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36482\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36374\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36331\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35981\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35800\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35728\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35703\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35463\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35156\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35030\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35000\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34874\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34714\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34187\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34172\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34039\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33842\ : std_logic;
signal \N__33839\ : std_logic;
signal \N__33836\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33816\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33800\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33791\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33464\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33275\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33247\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33167\ : std_logic;
signal \N__33164\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33104\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32601\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32522\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31562\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31151\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30407\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29899\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29501\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28283\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28132\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25430\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23215\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \ICE_GPMO_2\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\ : std_logic;
signal \ICE_SYSCLK\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\ : std_logic;
signal \RTD.n18092\ : std_logic;
signal \RTD_SCLK\ : std_logic;
signal \CLK_DDS.n16974\ : std_logic;
signal bit_cnt_0_adj_1498 : std_logic;
signal bit_cnt_3 : std_logic;
signal bit_cnt_2 : std_logic;
signal bit_cnt_1 : std_logic;
signal \n8_adj_1680_cascade_\ : std_logic;
signal n21625 : std_logic;
signal \RTD.n18043_cascade_\ : std_logic;
signal \RTD.n21494\ : std_logic;
signal \RTD.n21492_cascade_\ : std_logic;
signal \RTD.n7_adj_1435\ : std_logic;
signal \RTD.bit_cnt_2\ : std_logic;
signal \RTD.bit_cnt_1\ : std_logic;
signal \RTD.bit_cnt_0\ : std_logic;
signal \RTD_SDI\ : std_logic;
signal \RTD.n21471_cascade_\ : std_logic;
signal \RTD.n19032\ : std_logic;
signal \RTD.n4_cascade_\ : std_logic;
signal \RTD.n21387\ : std_logic;
signal \RTD.n21199_cascade_\ : std_logic;
signal \RTD.adc_state_3_N_1114_1\ : std_logic;
signal \RTD.n7_cascade_\ : std_logic;
signal \RTD.n11868\ : std_logic;
signal \RTD.n11860\ : std_logic;
signal \RTD.n8\ : std_logic;
signal adress_1 : std_logic;
signal adress_2 : std_logic;
signal adress_3 : std_logic;
signal adress_4 : std_logic;
signal adress_5 : std_logic;
signal \RTD_SDO\ : std_logic;
signal \RTD.n11915\ : std_logic;
signal n14692 : std_logic;
signal \RTD.n15280\ : std_logic;
signal read_buf_10 : std_logic;
signal \n13212_cascade_\ : std_logic;
signal read_buf_15 : std_logic;
signal \n11856_cascade_\ : std_logic;
signal read_buf_14 : std_logic;
signal \RTD.n12_adj_1445\ : std_logic;
signal \RTD.mode\ : std_logic;
signal read_buf_4 : std_logic;
signal read_buf_11 : std_logic;
signal read_buf_5 : std_logic;
signal read_buf_3 : std_logic;
signal \n19_adj_1600_cascade_\ : std_logic;
signal \n19_adj_1597_cascade_\ : std_logic;
signal buf_adcdata_vac_7 : std_logic;
signal cmd_rdadctmp_7_adj_1485 : std_logic;
signal \VAC_MISO\ : std_logic;
signal cmd_rdadctmp_0_adj_1492 : std_logic;
signal cmd_rdadctmp_1_adj_1491 : std_logic;
signal cmd_rdadctmp_2_adj_1490 : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \ADC_VAC.n19835\ : std_logic;
signal \ADC_VAC.n19836\ : std_logic;
signal \ADC_VAC.n19837\ : std_logic;
signal \ADC_VAC.n19838\ : std_logic;
signal \ADC_VAC.n19839\ : std_logic;
signal \ADC_VAC.n19840\ : std_logic;
signal \ADC_VAC.n19841\ : std_logic;
signal \ADC_VAC.bit_cnt_4\ : std_logic;
signal \ADC_VAC.bit_cnt_3\ : std_logic;
signal \ADC_VAC.bit_cnt_1\ : std_logic;
signal \ADC_VAC.bit_cnt_2\ : std_logic;
signal \ADC_VAC.bit_cnt_6\ : std_logic;
signal \ADC_VAC.bit_cnt_0\ : std_logic;
signal \ADC_VAC.n21224_cascade_\ : std_logic;
signal \ADC_VAC.bit_cnt_7\ : std_logic;
signal \ADC_VAC.bit_cnt_5\ : std_logic;
signal \ADC_VAC.n21234_cascade_\ : std_logic;
signal \ADC_VAC.n12803\ : std_logic;
signal \ADC_VAC.n15052\ : std_logic;
signal \ADC_VAC.n21157_cascade_\ : std_logic;
signal \ADC_VAC.n21468\ : std_logic;
signal \ADC_VAC.n21158\ : std_logic;
signal \RTD.n16766\ : std_logic;
signal \RTD_CS\ : std_logic;
signal \RTD.n14\ : std_logic;
signal \RTD.n21181_cascade_\ : std_logic;
signal \RTD.n13137_cascade_\ : std_logic;
signal \RTD.n7889\ : std_logic;
signal \RTD.bit_cnt_3\ : std_logic;
signal \RTD.n18043\ : std_logic;
signal \RTD.n19026\ : std_logic;
signal adress_6 : std_logic;
signal \RTD.n9_cascade_\ : std_logic;
signal \RTD.adress_7_N_1086_7_cascade_\ : std_logic;
signal \RTD_DRDY\ : std_logic;
signal \RTD.n11_cascade_\ : std_logic;
signal \RTD.n19_cascade_\ : std_logic;
signal \RTD.adress_7\ : std_logic;
signal \RTD.adress_7_N_1086_7\ : std_logic;
signal adress_0 : std_logic;
signal n13054 : std_logic;
signal \RTD.n20370\ : std_logic;
signal \RTD.cfg_buf_6\ : std_logic;
signal read_buf_9 : std_logic;
signal \RTD.adc_state_1\ : std_logic;
signal \RTD.n11829\ : std_logic;
signal read_buf_8 : std_logic;
signal read_buf_0 : std_logic;
signal read_buf_2 : std_logic;
signal n11856 : std_logic;
signal read_buf_1 : std_logic;
signal read_buf_12 : std_logic;
signal read_buf_13 : std_logic;
signal n13212 : std_logic;
signal n1_adj_1592 : std_logic;
signal read_buf_6 : std_logic;
signal read_buf_7 : std_logic;
signal buf_adcdata_iac_6 : std_logic;
signal buf_adcdata_vac_4 : std_logic;
signal \n19_adj_1606_cascade_\ : std_logic;
signal buf_data_iac_4 : std_logic;
signal \n22_adj_1607_cascade_\ : std_logic;
signal cmd_rdadctmp_31_adj_1461 : std_logic;
signal buf_adcdata_iac_7 : std_logic;
signal cmd_rdadctmp_8_adj_1484 : std_logic;
signal buf_data_iac_7 : std_logic;
signal n22_adj_1598 : std_logic;
signal cmd_rdadctmp_12_adj_1480 : std_logic;
signal buf_adcdata_iac_4 : std_logic;
signal \ADC_VAC.n17\ : std_logic;
signal \VAC_SCLK\ : std_logic;
signal cmd_rdadctmp_26_adj_1466 : std_logic;
signal cmd_rdadctmp_3_adj_1489 : std_logic;
signal \ADC_VAC.n12\ : std_logic;
signal n21050 : std_logic;
signal \VAC_DRDY\ : std_logic;
signal \n21050_cascade_\ : std_logic;
signal \VAC_CS\ : std_logic;
signal n14_adj_1657 : std_logic;
signal \DTRIG_N_958_adj_1493\ : std_logic;
signal adc_state_1_adj_1459 : std_logic;
signal cmd_rdadctmp_14 : std_logic;
signal \ADC_IAC.n21458_cascade_\ : std_logic;
signal \ADC_IAC.n16\ : std_logic;
signal \ADC_IAC.bit_cnt_0\ : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal \ADC_IAC.bit_cnt_1\ : std_logic;
signal \ADC_IAC.n19828\ : std_logic;
signal \ADC_IAC.bit_cnt_2\ : std_logic;
signal \ADC_IAC.n19829\ : std_logic;
signal \ADC_IAC.bit_cnt_3\ : std_logic;
signal \ADC_IAC.n19830\ : std_logic;
signal \ADC_IAC.bit_cnt_4\ : std_logic;
signal \ADC_IAC.n19831\ : std_logic;
signal \ADC_IAC.bit_cnt_5\ : std_logic;
signal \ADC_IAC.n19832\ : std_logic;
signal \ADC_IAC.bit_cnt_6\ : std_logic;
signal \ADC_IAC.n19833\ : std_logic;
signal \ADC_IAC.n19834\ : std_logic;
signal \ADC_IAC.bit_cnt_7\ : std_logic;
signal \ADC_IAC.n12698\ : std_logic;
signal \ADC_IAC.n12698_cascade_\ : std_logic;
signal \ADC_IAC.n15014\ : std_logic;
signal \AC_ADC_SYNC\ : std_logic;
signal \n14_adj_1662_cascade_\ : std_logic;
signal \IAC_CS\ : std_logic;
signal \DDS_CS1\ : std_logic;
signal \RTD.cfg_tmp_1\ : std_logic;
signal \RTD.cfg_tmp_2\ : std_logic;
signal \RTD.cfg_tmp_3\ : std_logic;
signal \RTD.cfg_tmp_4\ : std_logic;
signal \RTD.cfg_tmp_5\ : std_logic;
signal \RTD.cfg_tmp_6\ : std_logic;
signal \RTD.adc_state_0\ : std_logic;
signal \RTD.cfg_tmp_7\ : std_logic;
signal adc_state_2 : std_logic;
signal \RTD.cfg_tmp_0\ : std_logic;
signal \RTD.n13137\ : std_logic;
signal \RTD.n15115\ : std_logic;
signal \RTD.cfg_buf_5\ : std_logic;
signal \RTD.n11_adj_1444\ : std_logic;
signal \RTD.cfg_buf_3\ : std_logic;
signal \RTD.cfg_buf_4\ : std_logic;
signal \RTD.cfg_buf_2\ : std_logic;
signal \RTD.n10\ : std_logic;
signal \RTD.n11\ : std_logic;
signal \RTD.adc_state_3\ : std_logic;
signal \RTD.n21036\ : std_logic;
signal \RTD.n21199\ : std_logic;
signal \RTD.n13090_cascade_\ : std_logic;
signal \RTD.cfg_buf_1\ : std_logic;
signal \RTD.n12\ : std_logic;
signal \RTD.cfg_buf_7\ : std_logic;
signal \RTD.n13090\ : std_logic;
signal \RTD.n21061\ : std_logic;
signal \RTD.cfg_buf_0\ : std_logic;
signal \buf_readRTD_9\ : std_logic;
signal buf_adcdata_vdc_3 : std_logic;
signal buf_adcdata_iac_3 : std_logic;
signal \n19_adj_1609_cascade_\ : std_logic;
signal \buf_readRTD_14\ : std_logic;
signal cmd_rdadctmp_10_adj_1482 : std_logic;
signal \DDS_MOSI1\ : std_logic;
signal n20_adj_1693 : std_logic;
signal n22407 : std_logic;
signal buf_adcdata_vac_2 : std_logic;
signal \n19_adj_1612_cascade_\ : std_logic;
signal buf_adcdata_vac_6 : std_logic;
signal buf_adcdata_vac_22 : std_logic;
signal n22629 : std_logic;
signal cmd_rdadctmp_14_adj_1478 : std_logic;
signal cmd_rdadctmp_15_adj_1477 : std_logic;
signal buf_data_iac_6 : std_logic;
signal n22_adj_1601 : std_logic;
signal buf_data_iac_2 : std_logic;
signal n22_adj_1613 : std_logic;
signal \buf_readRTD_10\ : std_logic;
signal \buf_cfgRTD_2\ : std_logic;
signal cmd_rdadctmp_11_adj_1481 : std_logic;
signal buf_adcdata_vac_3 : std_logic;
signal cmd_rdadctmp_13_adj_1479 : std_logic;
signal cmd_rdadctmp_30_adj_1462 : std_logic;
signal buf_adcdata_vac_9 : std_logic;
signal cmd_rdadctmp_11 : std_logic;
signal cmd_rdadctmp_12 : std_logic;
signal cmd_rdadctmp_8 : std_logic;
signal cmd_rdadctmp_17_adj_1475 : std_logic;
signal cmd_rdadctmp_29_adj_1463 : std_logic;
signal cmd_rdadctmp_9_adj_1483 : std_logic;
signal \CLK_DDS.tmp_buf_10\ : std_logic;
signal \CLK_DDS.tmp_buf_11\ : std_logic;
signal \CLK_DDS.tmp_buf_12\ : std_logic;
signal \CLK_DDS.tmp_buf_13\ : std_logic;
signal \CLK_DDS.tmp_buf_14\ : std_logic;
signal \CLK_DDS.tmp_buf_9\ : std_logic;
signal \CLK_DDS.tmp_buf_8\ : std_logic;
signal \buf_readRTD_7\ : std_logic;
signal n16_adj_1690 : std_logic;
signal n17_adj_1691 : std_logic;
signal \ADC_IAC.n12\ : std_logic;
signal \ADC_IAC.n21457\ : std_logic;
signal cmd_rdadctmp_7 : std_logic;
signal cmd_rdadctmp_6 : std_logic;
signal n21082 : std_logic;
signal \n21082_cascade_\ : std_logic;
signal cmd_rdadctmp_3 : std_logic;
signal \n12771_cascade_\ : std_logic;
signal cmd_rdadctmp_4 : std_logic;
signal cmd_rdadctmp_5 : std_logic;
signal \ADC_IAC.n17\ : std_logic;
signal \DDS_MCLK1\ : std_logic;
signal cmd_rdadctmp_0_adj_1523 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_0\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_1\ : std_logic;
signal \ADC_VDC.n19842\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_2\ : std_logic;
signal \ADC_VDC.n19843\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_3\ : std_logic;
signal \ADC_VDC.n19844\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_4\ : std_logic;
signal \ADC_VDC.n19845\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_5\ : std_logic;
signal \ADC_VDC.n19846\ : std_logic;
signal cmd_rdadctmp_6_adj_1517 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_6\ : std_logic;
signal \ADC_VDC.n19847\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_7\ : std_logic;
signal \ADC_VDC.n19848\ : std_logic;
signal \ADC_VDC.n19849\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_8\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_9\ : std_logic;
signal \ADC_VDC.n19850\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_10\ : std_logic;
signal \ADC_VDC.n19851\ : std_logic;
signal \ADC_VDC.n19852\ : std_logic;
signal \ADC_VDC.n19853\ : std_logic;
signal \ADC_VDC.n19854\ : std_logic;
signal cmd_rdadcbuf_14 : std_logic;
signal \ADC_VDC.n19855\ : std_logic;
signal \ADC_VDC.n19856\ : std_logic;
signal \ADC_VDC.n19857\ : std_logic;
signal cmd_rdadctmp_16_adj_1507 : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal cmd_rdadctmp_17_adj_1506 : std_logic;
signal \ADC_VDC.n19858\ : std_logic;
signal cmd_rdadctmp_18_adj_1505 : std_logic;
signal \ADC_VDC.n19859\ : std_logic;
signal \ADC_VDC.n19860\ : std_logic;
signal \ADC_VDC.n19861\ : std_logic;
signal \ADC_VDC.n19862\ : std_logic;
signal \ADC_VDC.n19863\ : std_logic;
signal \ADC_VDC.n19864\ : std_logic;
signal \ADC_VDC.n19865\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \ADC_VDC.n19866\ : std_logic;
signal \ADC_VDC.n19867\ : std_logic;
signal \ADC_VDC.n19868\ : std_logic;
signal \ADC_VDC.n19869\ : std_logic;
signal cmd_rdadcbuf_29 : std_logic;
signal \ADC_VDC.n19870\ : std_logic;
signal \ADC_VDC.n19871\ : std_logic;
signal \ADC_VDC.n19872\ : std_logic;
signal \ADC_VDC.n19873\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \ADC_VDC.n19874\ : std_logic;
signal \ADC_VDC.n19875\ : std_logic;
signal buf_adcdata_vdc_18 : std_logic;
signal buf_adcdata_vac_18 : std_logic;
signal n19_adj_1692 : std_logic;
signal cmd_rdadctmp_13 : std_logic;
signal cmd_rdadctmp_10 : std_logic;
signal buf_adcdata_iac_2 : std_logic;
signal buf_adcdata_vac_5 : std_logic;
signal buf_adcdata_iac_5 : std_logic;
signal \n19_adj_1603_cascade_\ : std_logic;
signal \n22377_cascade_\ : std_logic;
signal n21237 : std_logic;
signal cmd_rdadctmp_28_adj_1464 : std_logic;
signal tmp_buf_15_adj_1497 : std_logic;
signal \CLK_DDS.tmp_buf_0\ : std_logic;
signal \CLK_DDS.tmp_buf_1\ : std_logic;
signal \CLK_DDS.tmp_buf_2\ : std_logic;
signal \CLK_DDS.tmp_buf_3\ : std_logic;
signal \CLK_DDS.tmp_buf_4\ : std_logic;
signal \CLK_DDS.tmp_buf_5\ : std_logic;
signal \CLK_DDS.tmp_buf_6\ : std_logic;
signal \CLK_DDS.tmp_buf_7\ : std_logic;
signal buf_adcdata_vac_17 : std_logic;
signal \SIG_DDS.bit_cnt_1\ : std_logic;
signal \SIG_DDS.bit_cnt_2\ : std_logic;
signal \SIG_DDS.n10\ : std_logic;
signal bit_cnt_0 : std_logic;
signal cmd_rdadctmp_4_adj_1488 : std_logic;
signal cmd_rdadctmp_5_adj_1487 : std_logic;
signal cmd_rdadctmp_6_adj_1486 : std_logic;
signal cmd_rdadctmp_22 : std_logic;
signal n15092 : std_logic;
signal \IAC_DRDY\ : std_logic;
signal \ADC_IAC.n21159_cascade_\ : std_logic;
signal \ADC_IAC.n21160\ : std_logic;
signal cmd_rdadctmp_1 : std_logic;
signal cmd_rdadctmp_2 : std_logic;
signal \IAC_MISO\ : std_logic;
signal cmd_rdadctmp_0 : std_logic;
signal \DTRIG_N_958\ : std_logic;
signal adc_state_1 : std_logic;
signal \IAC_SCLK\ : std_logic;
signal buf_adcdata_iac_17 : std_logic;
signal cmd_rdadcbuf_27 : std_logic;
signal \ADC_VDC.n10309_cascade_\ : std_logic;
signal \ADC_VDC.n13276\ : std_logic;
signal cmd_rdadctmp_1_adj_1522 : std_logic;
signal cmd_rdadctmp_2_adj_1521 : std_logic;
signal cmd_rdadctmp_3_adj_1520 : std_logic;
signal cmd_rdadctmp_4_adj_1519 : std_logic;
signal cmd_rdadctmp_5_adj_1518 : std_logic;
signal cmd_rdadctmp_7_adj_1516 : std_logic;
signal cmd_rdadctmp_19_adj_1504 : std_logic;
signal cmd_rdadctmp_8_adj_1515 : std_logic;
signal cmd_rdadctmp_9_adj_1514 : std_logic;
signal cmd_rdadctmp_10_adj_1513 : std_logic;
signal cmd_rdadctmp_11_adj_1512 : std_logic;
signal cmd_rdadctmp_12_adj_1511 : std_logic;
signal cmd_rdadctmp_13_adj_1510 : std_logic;
signal cmd_rdadctmp_14_adj_1509 : std_logic;
signal cmd_rdadctmp_15_adj_1508 : std_logic;
signal cmd_rdadcbuf_20 : std_logic;
signal buf_adcdata_vdc_9 : std_logic;
signal cmd_rdadcbuf_17 : std_logic;
signal buf_adcdata_vdc_6 : std_logic;
signal cmd_rdadcbuf_11 : std_logic;
signal buf_dds1_5 : std_logic;
signal cmd_rdadcbuf_21 : std_logic;
signal cmd_rdadcbuf_33 : std_logic;
signal buf_adcdata_vdc_22 : std_logic;
signal cmd_rdadcbuf_13 : std_logic;
signal buf_adcdata_vdc_2 : std_logic;
signal cmd_rdadcbuf_15 : std_logic;
signal buf_adcdata_vdc_4 : std_logic;
signal cmd_rdadcbuf_16 : std_logic;
signal buf_adcdata_vdc_5 : std_logic;
signal cmd_rdadctmp_20_adj_1503 : std_logic;
signal cmd_rdadctmp_21_adj_1502 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_35_N_1296_34\ : std_logic;
signal \ADC_VDC.n19\ : std_logic;
signal \ADC_VDC.n21_cascade_\ : std_logic;
signal cmd_rdadcbuf_34 : std_logic;
signal \ADC_VDC.n18780_cascade_\ : std_logic;
signal \ADC_VDC.n4_adj_1451\ : std_logic;
signal \ADC_VDC.n13503\ : std_logic;
signal \buf_readRTD_8\ : std_logic;
signal buf_adcdata_vdc_16 : std_logic;
signal buf_adcdata_vac_16 : std_logic;
signal \n22575_cascade_\ : std_logic;
signal \buf_cfgRTD_0\ : std_logic;
signal \n10902_cascade_\ : std_logic;
signal \n12624_cascade_\ : std_logic;
signal \buf_cfgRTD_3\ : std_logic;
signal \buf_readRTD_11\ : std_logic;
signal n22473 : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal n19813 : std_logic;
signal n19814 : std_logic;
signal n19815 : std_logic;
signal n19816 : std_logic;
signal n19817 : std_logic;
signal n19818 : std_logic;
signal n19819 : std_logic;
signal n19820 : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal n19821 : std_logic;
signal n19822 : std_logic;
signal n19823 : std_logic;
signal n19824 : std_logic;
signal n19825 : std_logic;
signal n19826 : std_logic;
signal n19827 : std_logic;
signal cmd_rdadctmp_27_adj_1465 : std_logic;
signal buf_adcdata_vac_19 : std_logic;
signal n12493 : std_logic;
signal n21705 : std_logic;
signal cmd_rdadctmp_18_adj_1474 : std_logic;
signal \IAC_OSR1\ : std_logic;
signal data_idxvec_11 : std_logic;
signal \n26_adj_1678_cascade_\ : std_logic;
signal n22509 : std_logic;
signal buf_dds1_2 : std_logic;
signal n22476 : std_logic;
signal cmd_rdadctmp_16_adj_1476 : std_logic;
signal cmd_rdadctmp_25_adj_1467 : std_logic;
signal cmd_rdadctmp_24_adj_1468 : std_logic;
signal cmd_rdadctmp_22_adj_1470 : std_logic;
signal cmd_rdadctmp_23_adj_1469 : std_logic;
signal n69 : std_logic;
signal cmd_rdadctmp_15 : std_logic;
signal \IAC_FLT1\ : std_logic;
signal buf_adcdata_iac_19 : std_logic;
signal \n22605_cascade_\ : std_logic;
signal buf_dds1_11 : std_logic;
signal n22608 : std_logic;
signal cmd_rdadctmp_27 : std_logic;
signal cmd_rdadctmp_19 : std_logic;
signal cmd_rdadctmp_24 : std_logic;
signal cmd_rdadctmp_30 : std_logic;
signal \ADC_VDC.n18780\ : std_logic;
signal \ADC_VDC.n18783_cascade_\ : std_logic;
signal \ADC_VDC.n16_adj_1450\ : std_logic;
signal \ADC_VDC.n18\ : std_logic;
signal \ADC_VDC.n18_cascade_\ : std_logic;
signal \THERMOSTAT\ : std_logic;
signal \ADC_VDC.avg_cnt_0\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \ADC_VDC.avg_cnt_1\ : std_logic;
signal \ADC_VDC.n19877\ : std_logic;
signal \ADC_VDC.avg_cnt_2\ : std_logic;
signal \ADC_VDC.n19878\ : std_logic;
signal \ADC_VDC.n19879\ : std_logic;
signal \ADC_VDC.avg_cnt_4\ : std_logic;
signal \ADC_VDC.n19880\ : std_logic;
signal \ADC_VDC.avg_cnt_5\ : std_logic;
signal \ADC_VDC.n19881\ : std_logic;
signal \ADC_VDC.n19882\ : std_logic;
signal \ADC_VDC.avg_cnt_7\ : std_logic;
signal \ADC_VDC.n19883\ : std_logic;
signal \ADC_VDC.n19884\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \ADC_VDC.n19885\ : std_logic;
signal \ADC_VDC.avg_cnt_10\ : std_logic;
signal \ADC_VDC.n19886\ : std_logic;
signal \ADC_VDC.n19887\ : std_logic;
signal \ADC_VDC.avg_cnt_11\ : std_logic;
signal \ADC_VDC.n13463\ : std_logic;
signal \ADC_VDC.n15175\ : std_logic;
signal cmd_rdadcbuf_23 : std_logic;
signal cmd_rdadcbuf_18 : std_logic;
signal buf_adcdata_vdc_7 : std_logic;
signal \n11891_cascade_\ : std_logic;
signal cmd_rdadcbuf_26 : std_logic;
signal cmd_rdadcbuf_25 : std_logic;
signal cmd_rdadcbuf_22 : std_logic;
signal buf_control_7 : std_logic;
signal \DDS_SCK1\ : std_logic;
signal \buf_readRTD_15\ : std_logic;
signal buf_adcdata_vdc_23 : std_logic;
signal \n22593_cascade_\ : std_logic;
signal buf_adcdata_vac_23 : std_logic;
signal \buf_cfgRTD_6\ : std_logic;
signal \buf_cfgRTD_7\ : std_logic;
signal n30_adj_1499 : std_logic;
signal cmd_rdadctmp_19_adj_1473 : std_logic;
signal buf_adcdata_vac_21 : std_logic;
signal \VAC_OSR1\ : std_logic;
signal buf_adcdata_vdc_10 : std_logic;
signal buf_adcdata_vac_10 : std_logic;
signal buf_adcdata_vdc_0 : std_logic;
signal buf_adcdata_vac_0 : std_logic;
signal buf_adcdata_iac_0 : std_logic;
signal \n19_adj_1534_cascade_\ : std_logic;
signal n19_adj_1652 : std_logic;
signal \buf_readRTD_1\ : std_logic;
signal buf_adcdata_vac_13 : std_logic;
signal \buf_readRTD_5\ : std_logic;
signal \n19_adj_1629_cascade_\ : std_logic;
signal n12850 : std_logic;
signal cmd_rdadctmp_21_adj_1471 : std_logic;
signal n8 : std_logic;
signal n10695 : std_logic;
signal buf_adcdata_vdc_12 : std_logic;
signal n21076 : std_logic;
signal adc_state_0_adj_1460 : std_logic;
signal cmd_rdadctmp_20_adj_1472 : std_logic;
signal buf_adcdata_vac_12 : std_logic;
signal \iac_raw_buf_N_774\ : std_logic;
signal n21334 : std_logic;
signal n22512 : std_logic;
signal data_idxvec_15 : std_logic;
signal buf_data_iac_23 : std_logic;
signal \n26_adj_1659_cascade_\ : std_logic;
signal \n21324_cascade_\ : std_logic;
signal buf_adcdata_vac_15 : std_logic;
signal buf_adcdata_vdc_15 : std_logic;
signal n19_adj_1621 : std_logic;
signal n23_adj_1658 : std_logic;
signal n21323 : std_logic;
signal n22371 : std_logic;
signal \n12_adj_1454_cascade_\ : std_logic;
signal acadc_trig : std_logic;
signal n21053 : std_logic;
signal \n21042_cascade_\ : std_logic;
signal \n21030_cascade_\ : std_logic;
signal eis_end : std_logic;
signal \INVacadc_trig_300C_net\ : std_logic;
signal n17728 : std_logic;
signal \n11_cascade_\ : std_logic;
signal acadc_dtrig_v : std_logic;
signal acadc_dtrig_i : std_logic;
signal \eis_state_2_N_392_1\ : std_logic;
signal \eis_state_2_N_392_1_cascade_\ : std_logic;
signal \n2_adj_1696_cascade_\ : std_logic;
signal n22437 : std_logic;
signal \INVeis_state_i1C_net\ : std_logic;
signal cmd_rdadctmp_23 : std_logic;
signal \VAC_FLT1\ : std_logic;
signal cmd_rdadctmp_29 : std_logic;
signal buf_adcdata_iac_21 : std_logic;
signal cmd_rdadctmp_28 : std_logic;
signal cmd_rdadctmp_25 : std_logic;
signal cmd_rdadctmp_20 : std_logic;
signal n12771 : std_logic;
signal cmd_rdadctmp_31 : std_logic;
signal buf_adcdata_iac_23 : std_logic;
signal \ADC_VDC.n16\ : std_logic;
signal \ADC_VDC.n21593_cascade_\ : std_logic;
signal \ADC_VDC.n21590_cascade_\ : std_logic;
signal \ADC_VDC.n22590\ : std_logic;
signal n13324 : std_logic;
signal \ADC_VDC.n7_cascade_\ : std_logic;
signal \ADC_VDC.n21193\ : std_logic;
signal cmd_rdadcbuf_19 : std_logic;
signal cmd_rdadcbuf_24 : std_logic;
signal buf_adcdata_vdc_13 : std_logic;
signal cmd_rdadcbuf_30 : std_logic;
signal buf_adcdata_vdc_19 : std_logic;
signal cmd_rdadcbuf_28 : std_logic;
signal buf_adcdata_vdc_17 : std_logic;
signal cmd_rdadcbuf_32 : std_logic;
signal buf_adcdata_vdc_21 : std_logic;
signal cmd_rdadcbuf_31 : std_logic;
signal buf_dds1_4 : std_logic;
signal \ADC_VDC.n22587\ : std_logic;
signal \ADC_VDC.n10708\ : std_logic;
signal cmd_rdadctmp_22_adj_1501 : std_logic;
signal \ADC_VDC.n10708_cascade_\ : std_logic;
signal \ADC_VDC.cmd_rdadctmp_23\ : std_logic;
signal \ADC_VDC.n5\ : std_logic;
signal \ADC_VDC.avg_cnt_9\ : std_logic;
signal \ADC_VDC.avg_cnt_8\ : std_logic;
signal \ADC_VDC.avg_cnt_6\ : std_logic;
signal \ADC_VDC.avg_cnt_3\ : std_logic;
signal \ADC_VDC.n20\ : std_logic;
signal \CLK_DDS.n13005\ : std_logic;
signal \CLK_DDS.n9_adj_1433\ : std_logic;
signal dds_state_2_adj_1494 : std_logic;
signal dds_state_0_adj_1496 : std_logic;
signal dds_state_1_adj_1495 : std_logic;
signal \CLK_DDS.n9\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal n19956 : std_logic;
signal n19957 : std_logic;
signal n19958 : std_logic;
signal n19959 : std_logic;
signal n19960 : std_logic;
signal n19961 : std_logic;
signal n19962 : std_logic;
signal n19963 : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal n19964 : std_logic;
signal n19965 : std_logic;
signal n19966 : std_logic;
signal n19967 : std_logic;
signal n19968 : std_logic;
signal n19969 : std_logic;
signal n19970 : std_logic;
signal n19971 : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal n19972 : std_logic;
signal n19973 : std_logic;
signal n19974 : std_logic;
signal n19975 : std_logic;
signal n19976 : std_logic;
signal n19977 : std_logic;
signal secclk_cnt_21 : std_logic;
signal secclk_cnt_19 : std_logic;
signal secclk_cnt_12 : std_logic;
signal secclk_cnt_22 : std_logic;
signal n14_adj_1571 : std_logic;
signal n21329 : std_logic;
signal \IAC_FLT0\ : std_logic;
signal n22374 : std_logic;
signal n21240 : std_logic;
signal n22401 : std_logic;
signal n21122 : std_logic;
signal \n21122_cascade_\ : std_logic;
signal \n12610_cascade_\ : std_logic;
signal buf_data_iac_5 : std_logic;
signal n22_adj_1604 : std_logic;
signal data_idxvec_4 : std_logic;
signal \n26_adj_1635_cascade_\ : std_logic;
signal \n22443_cascade_\ : std_logic;
signal \n22446_cascade_\ : std_logic;
signal \n30_adj_1636_cascade_\ : std_logic;
signal n19_adj_1634 : std_logic;
signal \buf_readRTD_4\ : std_logic;
signal buf_adcdata_iac_12 : std_logic;
signal \n22467_cascade_\ : std_logic;
signal n16_adj_1633 : std_logic;
signal n22470 : std_logic;
signal \n22395_cascade_\ : std_logic;
signal req_data_cnt_8 : std_logic;
signal \VAC_FLT0\ : std_logic;
signal buf_adcdata_iac_22 : std_logic;
signal \n22635_cascade_\ : std_logic;
signal n21236 : std_logic;
signal n14_adj_1578 : std_logic;
signal \n2_cascade_\ : std_logic;
signal \n21501_cascade_\ : std_logic;
signal \eis_state_2_N_392_0\ : std_logic;
signal n22479 : std_logic;
signal eis_start : std_logic;
signal \n11_adj_1632_cascade_\ : std_logic;
signal \INVeis_state_i0C_net\ : std_logic;
signal n11908 : std_logic;
signal eis_state_0 : std_logic;
signal n21041 : std_logic;
signal buf_dds1_15 : std_logic;
signal buf_dds1_10 : std_logic;
signal \acadc_skipCount_15\ : std_logic;
signal n11570 : std_logic;
signal \EIS_SYNCCLK\ : std_logic;
signal \IAC_CLK\ : std_logic;
signal buf_dds0_10 : std_logic;
signal \SIG_DDS.tmp_buf_10\ : std_logic;
signal buf_dds0_11 : std_logic;
signal \SIG_DDS.tmp_buf_11\ : std_logic;
signal \SIG_DDS.tmp_buf_12\ : std_logic;
signal \SIG_DDS.tmp_buf_13\ : std_logic;
signal buf_dds0_14 : std_logic;
signal buf_dds0_15 : std_logic;
signal \SIG_DDS.tmp_buf_14\ : std_logic;
signal buf_dds0_9 : std_logic;
signal \SIG_DDS.tmp_buf_9\ : std_logic;
signal \SIG_DDS.tmp_buf_8\ : std_logic;
signal \SIG_DDS.tmp_buf_0\ : std_logic;
signal buf_dds0_1 : std_logic;
signal \SIG_DDS.tmp_buf_1\ : std_logic;
signal buf_dds0_2 : std_logic;
signal \SIG_DDS.tmp_buf_2\ : std_logic;
signal \SIG_DDS.tmp_buf_3\ : std_logic;
signal \SIG_DDS.tmp_buf_4\ : std_logic;
signal \SIG_DDS.tmp_buf_5\ : std_logic;
signal \ADC_VDC.n21007\ : std_logic;
signal \ADC_VDC.n21007_cascade_\ : std_logic;
signal \ADC_VDC.n4\ : std_logic;
signal \ADC_VDC.n11\ : std_logic;
signal \ADC_VDC.n65\ : std_logic;
signal \ADC_VDC.n21133\ : std_logic;
signal \ADC_VDC.n42_adj_1452\ : std_logic;
signal \ADC_VDC.n20998\ : std_logic;
signal \ADC_VDC.n11494\ : std_logic;
signal \ADC_VDC.n11494_cascade_\ : std_logic;
signal \ADC_VDC.n15\ : std_logic;
signal \ADC_VDC.n15_cascade_\ : std_logic;
signal \ADC_VDC.n21185\ : std_logic;
signal n11891 : std_logic;
signal cmd_rdadcbuf_12 : std_logic;
signal \ADC_VDC.n21203\ : std_logic;
signal \ADC_VDC.n21211\ : std_logic;
signal \ADC_VDC.n13368\ : std_logic;
signal secclk_cnt_20 : std_logic;
signal \n20048_cascade_\ : std_logic;
signal n14 : std_logic;
signal buf_adcdata_vdc_20 : std_logic;
signal buf_adcdata_vac_20 : std_logic;
signal secclk_cnt_6 : std_logic;
signal secclk_cnt_14 : std_logic;
signal secclk_cnt_10 : std_logic;
signal secclk_cnt_3 : std_logic;
signal n27 : std_logic;
signal secclk_cnt_2 : std_logic;
signal secclk_cnt_13 : std_logic;
signal secclk_cnt_7 : std_logic;
signal secclk_cnt_16 : std_logic;
signal n26_adj_1656 : std_logic;
signal n14_adj_1552 : std_logic;
signal n30 : std_logic;
signal n14_adj_1574 : std_logic;
signal buf_data_iac_3 : std_logic;
signal n22_adj_1610 : std_logic;
signal req_data_cnt_14 : std_logic;
signal req_data_cnt_11 : std_logic;
signal n23 : std_logic;
signal n14_adj_1551 : std_logic;
signal buf_dds0_4 : std_logic;
signal n23_adj_1661 : std_logic;
signal \acadc_skipCount_14\ : std_logic;
signal buf_adcdata_vdc_1 : std_logic;
signal buf_adcdata_vac_1 : std_logic;
signal buf_adcdata_iac_20 : std_logic;
signal \VAC_OSR0\ : std_logic;
signal comm_cmd_4 : std_logic;
signal \n16818_cascade_\ : std_logic;
signal n16_adj_1628 : std_logic;
signal n22365 : std_logic;
signal data_idxvec_5 : std_logic;
signal \n26_adj_1630_cascade_\ : std_logic;
signal \n22449_cascade_\ : std_logic;
signal req_data_cnt_5 : std_logic;
signal n22368 : std_logic;
signal \n22452_cascade_\ : std_logic;
signal \n30_adj_1631_cascade_\ : std_logic;
signal n9 : std_logic;
signal buf_data_iac_22 : std_logic;
signal data_idxvec_14 : std_logic;
signal n21330 : std_logic;
signal \acadc_skipCount_11\ : std_logic;
signal n23_adj_1677 : std_logic;
signal buf_dds1_9 : std_logic;
signal buf_adcdata_vdc_14 : std_logic;
signal buf_adcdata_vac_14 : std_logic;
signal n20 : std_logic;
signal \n17_cascade_\ : std_logic;
signal n19_adj_1526 : std_logic;
signal n29 : std_logic;
signal data_idxvec_13 : std_logic;
signal buf_dds1_3 : std_logic;
signal \acadc_skipCount_4\ : std_logic;
signal n8_adj_1560 : std_logic;
signal \n8_adj_1560_cascade_\ : std_logic;
signal \data_index_9_N_212_7\ : std_logic;
signal n24_adj_1593 : std_logic;
signal n23_adj_1591 : std_logic;
signal \n22_adj_1590_cascade_\ : std_logic;
signal n18 : std_logic;
signal \n30_adj_1543_cascade_\ : std_logic;
signal n31_adj_1537 : std_logic;
signal cmd_rdadctmp_26 : std_logic;
signal buf_adcdata_iac_18 : std_logic;
signal \acadc_skipCount_8\ : std_logic;
signal \n14_adj_1538_cascade_\ : std_logic;
signal n26_adj_1525 : std_logic;
signal cmd_rdadctmp_21 : std_logic;
signal buf_adcdata_iac_13 : std_logic;
signal \acadc_skipCount_13\ : std_logic;
signal buf_dds0_5 : std_logic;
signal buf_dds0_3 : std_logic;
signal \acadc_skipCount_5\ : std_logic;
signal n20_adj_1670 : std_logic;
signal cmd_rdadctmp_16 : std_logic;
signal cmd_rdadctmp_17 : std_logic;
signal data_count_0 : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal data_count_1 : std_logic;
signal n19765 : std_logic;
signal data_count_2 : std_logic;
signal n19766 : std_logic;
signal data_count_3 : std_logic;
signal n19767 : std_logic;
signal data_count_4 : std_logic;
signal n19768 : std_logic;
signal data_count_5 : std_logic;
signal n19769 : std_logic;
signal data_count_6 : std_logic;
signal n19770 : std_logic;
signal data_count_7 : std_logic;
signal n19771 : std_logic;
signal n19772 : std_logic;
signal \INVdata_count_i0_i0C_net\ : std_logic;
signal data_count_8 : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal n19773 : std_logic;
signal data_count_9 : std_logic;
signal \INVdata_count_i0_i8C_net\ : std_logic;
signal \comm_spi.n23089\ : std_logic;
signal \comm_spi.n14822\ : std_logic;
signal \comm_spi.n23089_cascade_\ : std_logic;
signal \comm_spi.n14823\ : std_logic;
signal \ADC_VDC.bit_cnt_0\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \ADC_VDC.bit_cnt_1\ : std_logic;
signal \ADC_VDC.n19918\ : std_logic;
signal \ADC_VDC.bit_cnt_2\ : std_logic;
signal \ADC_VDC.n19919\ : std_logic;
signal \ADC_VDC.bit_cnt_3\ : std_logic;
signal \ADC_VDC.n19920\ : std_logic;
signal \ADC_VDC.bit_cnt_4\ : std_logic;
signal \ADC_VDC.n19921\ : std_logic;
signal \ADC_VDC.bit_cnt_5\ : std_logic;
signal \ADC_VDC.n19922\ : std_logic;
signal \ADC_VDC.bit_cnt_6\ : std_logic;
signal \ADC_VDC.n19923\ : std_logic;
signal \ADC_VDC.n19924\ : std_logic;
signal \ADC_VDC.bit_cnt_7\ : std_logic;
signal \ADC_VDC.n15273\ : std_logic;
signal n21_adj_1594 : std_logic;
signal n14899 : std_logic;
signal \TEST_LED\ : std_logic;
signal secclk_cnt_15 : std_logic;
signal secclk_cnt_8 : std_logic;
signal secclk_cnt_1 : std_logic;
signal secclk_cnt_5 : std_logic;
signal n25 : std_logic;
signal secclk_cnt_18 : std_logic;
signal secclk_cnt_0 : std_logic;
signal secclk_cnt_11 : std_logic;
signal secclk_cnt_4 : std_logic;
signal n28_adj_1554 : std_logic;
signal req_data_cnt_15 : std_logic;
signal n24 : std_logic;
signal req_data_cnt_12 : std_logic;
signal n22 : std_logic;
signal n14_adj_1548 : std_logic;
signal \comm_spi.n23095\ : std_logic;
signal \comm_spi.data_tx_7__N_807\ : std_logic;
signal req_data_cnt_13 : std_logic;
signal secclk_cnt_9 : std_logic;
signal secclk_cnt_17 : std_logic;
signal n10 : std_logic;
signal n19_adj_1683 : std_logic;
signal n20_adj_1684 : std_logic;
signal buf_adcdata_vdc_11 : std_logic;
signal buf_adcdata_vac_11 : std_logic;
signal \buf_readRTD_12\ : std_logic;
signal \buf_cfgRTD_4\ : std_logic;
signal buf_dds1_13 : std_logic;
signal \buf_cfgRTD_5\ : std_logic;
signal \buf_readRTD_13\ : std_logic;
signal n9269 : std_logic;
signal \n12082_cascade_\ : std_logic;
signal n14_adj_1573 : std_logic;
signal \comm_spi.data_tx_7__N_817\ : std_logic;
signal req_data_cnt_10 : std_logic;
signal n19_adj_1646 : std_logic;
signal \buf_readRTD_2\ : std_logic;
signal n16_adj_1645 : std_logic;
signal \n22641_cascade_\ : std_logic;
signal data_idxvec_2 : std_logic;
signal \n26_adj_1647_cascade_\ : std_logic;
signal \acadc_skipCount_2\ : std_logic;
signal \n22383_cascade_\ : std_logic;
signal req_data_cnt_2 : std_logic;
signal n22644 : std_logic;
signal \n22386_cascade_\ : std_logic;
signal \n30_adj_1648_cascade_\ : std_logic;
signal req_data_cnt_4 : std_logic;
signal n18_adj_1644 : std_logic;
signal buf_dds0_13 : std_logic;
signal n66 : std_logic;
signal buf_dds1_14 : std_logic;
signal buf_dds1_1 : std_logic;
signal n12662 : std_logic;
signal n5_adj_1536 : std_logic;
signal \n7_adj_1650_cascade_\ : std_logic;
signal n12 : std_logic;
signal \SELIRNG1\ : std_logic;
signal n14_adj_1546 : std_logic;
signal n14_adj_1549 : std_logic;
signal n8_adj_1562 : std_logic;
signal \data_index_9_N_212_6\ : std_logic;
signal n17_adj_1553 : std_logic;
signal \AMPV_POW\ : std_logic;
signal \data_index_9_N_212_3\ : std_logic;
signal eis_state_1 : std_logic;
signal eis_state_2 : std_logic;
signal acadc_rst : std_logic;
signal n20011 : std_logic;
signal n19_adj_1616 : std_logic;
signal n14_adj_1547 : std_logic;
signal \n8_adj_1564_cascade_\ : std_logic;
signal \data_index_9_N_212_4\ : std_logic;
signal cmd_rdadctmp_9 : std_logic;
signal buf_adcdata_iac_1 : std_logic;
signal buf_dds1_12 : std_logic;
signal buf_dds0_12 : std_logic;
signal n8_adj_1566 : std_logic;
signal \n8_adj_1566_cascade_\ : std_logic;
signal \SIG_DDS.tmp_buf_6\ : std_logic;
signal \SIG_DDS.tmp_buf_7\ : std_logic;
signal \SIG_DDS.bit_cnt_3\ : std_logic;
signal \SIG_DDS.n21744\ : std_logic;
signal buf_dds1_7 : std_logic;
signal acadc_skipcnt_0 : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \INVacadc_skipcnt_i0_i0C_net\ : std_logic;
signal n21226 : std_logic;
signal n19789 : std_logic;
signal \n19789_THRU_CRY_0_THRU_CO\ : std_logic;
signal \n19789_THRU_CRY_1_THRU_CO\ : std_logic;
signal \n19789_THRU_CRY_2_THRU_CO\ : std_logic;
signal \n19789_THRU_CRY_3_THRU_CO\ : std_logic;
signal \n19789_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n19789_THRU_CRY_5_THRU_CO\ : std_logic;
signal \n19789_THRU_CRY_6_THRU_CO\ : std_logic;
signal acadc_skipcnt_1 : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal acadc_skipcnt_2 : std_logic;
signal n19790 : std_logic;
signal acadc_skipcnt_3 : std_logic;
signal n19791 : std_logic;
signal acadc_skipcnt_4 : std_logic;
signal n19792 : std_logic;
signal acadc_skipcnt_5 : std_logic;
signal n19793 : std_logic;
signal acadc_skipcnt_6 : std_logic;
signal n19794 : std_logic;
signal acadc_skipcnt_7 : std_logic;
signal n19795 : std_logic;
signal acadc_skipcnt_8 : std_logic;
signal n19796 : std_logic;
signal n19797 : std_logic;
signal \INVacadc_skipcnt_i0_i1C_net\ : std_logic;
signal acadc_skipcnt_9 : std_logic;
signal \bfn_13_20_0_\ : std_logic;
signal n19798 : std_logic;
signal acadc_skipcnt_11 : std_logic;
signal n19799 : std_logic;
signal n19800 : std_logic;
signal acadc_skipcnt_13 : std_logic;
signal n19801 : std_logic;
signal acadc_skipcnt_14 : std_logic;
signal n19802 : std_logic;
signal n19803 : std_logic;
signal acadc_skipcnt_15 : std_logic;
signal \INVacadc_skipcnt_i0_i9C_net\ : std_logic;
signal n11989 : std_logic;
signal n14915 : std_logic;
signal \INVcomm_spi.imiso_83_12297_12298_resetC_net\ : std_logic;
signal \comm_spi.n23083\ : std_logic;
signal \comm_spi.n14846\ : std_logic;
signal \comm_spi.n14847\ : std_logic;
signal \INVADC_VDC.genclk.t_clk_24C_net\ : std_logic;
signal \comm_spi.n14808\ : std_logic;
signal \comm_spi.n14809\ : std_logic;
signal \comm_spi.imosi_cascade_\ : std_logic;
signal \comm_spi.DOUT_7__N_786\ : std_logic;
signal \comm_spi.imosi_N_792\ : std_logic;
signal \n12_adj_1542_cascade_\ : std_logic;
signal \n19986_cascade_\ : std_logic;
signal n30_adj_1530 : std_logic;
signal n33 : std_logic;
signal \n34_cascade_\ : std_logic;
signal n31 : std_logic;
signal \n49_cascade_\ : std_logic;
signal n32 : std_logic;
signal \INVcomm_spi.bit_cnt_3767__i3C_net\ : std_logic;
signal n19_adj_1673 : std_logic;
signal n20_adj_1674 : std_logic;
signal \comm_spi.bit_cnt_1\ : std_logic;
signal \comm_spi.bit_cnt_2\ : std_logic;
signal \comm_spi.bit_cnt_0\ : std_logic;
signal n14_adj_1579 : std_logic;
signal n14_adj_1572 : std_logic;
signal n4_adj_1637 : std_logic;
signal n14_adj_1544 : std_logic;
signal n14_adj_1575 : std_logic;
signal n19_adj_1666 : std_logic;
signal n20_adj_1667 : std_logic;
signal n16_adj_1664 : std_logic;
signal n17_adj_1665 : std_logic;
signal \n22413_cascade_\ : std_logic;
signal n21671 : std_logic;
signal n23_adj_1668 : std_logic;
signal \n22569_cascade_\ : std_logic;
signal n21702 : std_logic;
signal n22416 : std_logic;
signal \n22572_cascade_\ : std_logic;
signal \n30_adj_1669_cascade_\ : std_logic;
signal n22404 : std_logic;
signal n22380 : std_logic;
signal n30_adj_1679 : std_logic;
signal \n8_adj_1689_cascade_\ : std_logic;
signal \n26_adj_1595_cascade_\ : std_logic;
signal n18_adj_1615 : std_logic;
signal n16818 : std_logic;
signal n21714 : std_logic;
signal \n7_cascade_\ : std_logic;
signal n12107 : std_logic;
signal \iac_raw_buf_N_776\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal n19774 : std_logic;
signal data_cntvec_2 : std_logic;
signal n19775 : std_logic;
signal n19776 : std_logic;
signal data_cntvec_4 : std_logic;
signal n19777 : std_logic;
signal data_cntvec_5 : std_logic;
signal n19778 : std_logic;
signal n19779 : std_logic;
signal n19780 : std_logic;
signal n19781 : std_logic;
signal \INVdata_cntvec_i0_i0C_net\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal n19782 : std_logic;
signal n19783 : std_logic;
signal data_cntvec_11 : std_logic;
signal n19784 : std_logic;
signal data_cntvec_12 : std_logic;
signal n19785 : std_logic;
signal data_cntvec_13 : std_logic;
signal n19786 : std_logic;
signal data_cntvec_14 : std_logic;
signal n19787 : std_logic;
signal n19788 : std_logic;
signal data_cntvec_15 : std_logic;
signal \INVdata_cntvec_i0_i8C_net\ : std_logic;
signal n11933 : std_logic;
signal n14907 : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal n19804 : std_logic;
signal n19805 : std_logic;
signal data_index_3 : std_logic;
signal n7_adj_1565 : std_logic;
signal n19806 : std_logic;
signal n19807 : std_logic;
signal n19808 : std_logic;
signal data_index_6 : std_logic;
signal n7_adj_1561 : std_logic;
signal n19809 : std_logic;
signal data_index_7 : std_logic;
signal n7_adj_1559 : std_logic;
signal n19810 : std_logic;
signal n19811 : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal n10756 : std_logic;
signal n19812 : std_logic;
signal buf_data_iac_1 : std_logic;
signal n22_adj_1617 : std_logic;
signal trig_dds1 : std_logic;
signal buf_dds0_7 : std_logic;
signal n21079 : std_logic;
signal adc_state_0 : std_logic;
signal cmd_rdadctmp_18 : std_logic;
signal buf_adcdata_iac_10 : std_logic;
signal n8_adj_1564 : std_logic;
signal n7_adj_1563 : std_logic;
signal data_index_4 : std_logic;
signal n11611 : std_logic;
signal buf_adcdata_iac_16 : std_logic;
signal buf_dds1_8 : std_logic;
signal \n22389_cascade_\ : std_logic;
signal buf_dds0_8 : std_logic;
signal data_index_5 : std_logic;
signal \DDS_SCK\ : std_logic;
signal tmp_buf_15 : std_logic;
signal \DDS_MOSI\ : std_logic;
signal data_index_9 : std_logic;
signal n12624 : std_logic;
signal \buf_cfgRTD_1\ : std_logic;
signal n12610 : std_logic;
signal \IAC_OSR0\ : std_logic;
signal \data_index_9_N_212_8\ : std_logic;
signal data_index_1 : std_logic;
signal n8_adj_1570 : std_logic;
signal \n8_adj_1570_cascade_\ : std_logic;
signal n7_adj_1569 : std_logic;
signal \data_index_9_N_212_1\ : std_logic;
signal data_index_2 : std_logic;
signal n8_adj_1558 : std_logic;
signal n7_adj_1557 : std_logic;
signal data_index_8 : std_logic;
signal n8_adj_1568 : std_logic;
signal n7_adj_1567 : std_logic;
signal \data_index_9_N_212_2\ : std_logic;
signal \comm_spi.n14815\ : std_logic;
signal \comm_spi.n14816\ : std_logic;
signal \INVcomm_spi.imiso_83_12297_12298_setC_net\ : std_logic;
signal \comm_spi.imosi\ : std_logic;
signal \comm_spi.DOUT_7__N_787\ : std_logic;
signal wdtick_cnt_0 : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal wdtick_cnt_1 : std_logic;
signal n19932 : std_logic;
signal wdtick_cnt_2 : std_logic;
signal n19933 : std_logic;
signal wdtick_cnt_3 : std_logic;
signal n19934 : std_logic;
signal wdtick_cnt_4 : std_logic;
signal n19935 : std_logic;
signal wdtick_cnt_5 : std_logic;
signal n19936 : std_logic;
signal wdtick_cnt_6 : std_logic;
signal n19937 : std_logic;
signal wdtick_cnt_7 : std_logic;
signal n19938 : std_logic;
signal n19939 : std_logic;
signal wdtick_cnt_8 : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal wdtick_cnt_9 : std_logic;
signal n19940 : std_logic;
signal wdtick_cnt_10 : std_logic;
signal n19941 : std_logic;
signal wdtick_cnt_11 : std_logic;
signal n19942 : std_logic;
signal wdtick_cnt_12 : std_logic;
signal n19943 : std_logic;
signal wdtick_cnt_13 : std_logic;
signal n19944 : std_logic;
signal wdtick_cnt_14 : std_logic;
signal n19945 : std_logic;
signal wdtick_cnt_15 : std_logic;
signal n19946 : std_logic;
signal n19947 : std_logic;
signal wdtick_cnt_16 : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal wdtick_cnt_17 : std_logic;
signal n19948 : std_logic;
signal wdtick_cnt_18 : std_logic;
signal n19949 : std_logic;
signal wdtick_cnt_19 : std_logic;
signal n19950 : std_logic;
signal wdtick_cnt_20 : std_logic;
signal n19951 : std_logic;
signal wdtick_cnt_21 : std_logic;
signal n19952 : std_logic;
signal wdtick_cnt_22 : std_logic;
signal n19953 : std_logic;
signal wdtick_cnt_23 : std_logic;
signal n19954 : std_logic;
signal n19955 : std_logic;
signal n49 : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal wdtick_cnt_24 : std_logic;
signal \clk_RTD\ : std_logic;
signal n14_adj_1550 : std_logic;
signal n17_adj_1672 : std_logic;
signal n22461 : std_logic;
signal n16_adj_1671 : std_logic;
signal data_idxvec_12 : std_logic;
signal \n21556_cascade_\ : std_logic;
signal n21703 : std_logic;
signal n22521 : std_logic;
signal n22464 : std_logic;
signal \n22524_cascade_\ : std_logic;
signal \n30_adj_1676_cascade_\ : std_logic;
signal n17_adj_1682 : std_logic;
signal n16_adj_1681 : std_logic;
signal n22485 : std_logic;
signal data_idxvec_10 : std_logic;
signal data_cntvec_10 : std_logic;
signal \n26_adj_1687_cascade_\ : std_logic;
signal \n22455_cascade_\ : std_logic;
signal n24_adj_1686 : std_logic;
signal n22488 : std_logic;
signal \n22458_cascade_\ : std_logic;
signal \n30_adj_1688_cascade_\ : std_logic;
signal data_idxvec_8 : std_logic;
signal data_cntvec_8 : std_logic;
signal buf_data_iac_16 : std_logic;
signal \n26_adj_1533_cascade_\ : std_logic;
signal n22398 : std_logic;
signal \n21246_cascade_\ : std_logic;
signal n22392 : std_logic;
signal n22578 : std_logic;
signal \n22581_cascade_\ : std_logic;
signal \n22584_cascade_\ : std_logic;
signal \buf_readRTD_3\ : std_logic;
signal n19_adj_1641 : std_logic;
signal buf_adcdata_iac_11 : std_logic;
signal n16_adj_1640 : std_logic;
signal \n22623_cascade_\ : std_logic;
signal \n22626_cascade_\ : std_logic;
signal n30_adj_1643 : std_logic;
signal data_idxvec_3 : std_logic;
signal data_cntvec_3 : std_logic;
signal \n26_adj_1642_cascade_\ : std_logic;
signal req_data_cnt_3 : std_logic;
signal \n22425_cascade_\ : std_logic;
signal \acadc_skipCount_3\ : std_logic;
signal n22428 : std_logic;
signal data_index_0 : std_logic;
signal n8841 : std_logic;
signal n8_adj_1540 : std_logic;
signal n7_adj_1539 : std_logic;
signal \n8_adj_1540_cascade_\ : std_logic;
signal \data_index_9_N_212_0\ : std_logic;
signal buf_dds1_0 : std_logic;
signal \n16_cascade_\ : std_logic;
signal buf_adcdata_iac_8 : std_logic;
signal n12596 : std_logic;
signal buf_dds0_0 : std_logic;
signal \VDC_RNG0\ : std_logic;
signal n23_adj_1675 : std_logic;
signal buf_dds0_6 : std_logic;
signal n17705 : std_logic;
signal \n9342_cascade_\ : std_logic;
signal n17703 : std_logic;
signal \data_index_9_N_212_5\ : std_logic;
signal buf_adcdata_iac_15 : std_logic;
signal n16_adj_1620 : std_logic;
signal n12144 : std_logic;
signal \DDS_CS\ : std_logic;
signal \SIG_DDS.n9_adj_1434\ : std_logic;
signal n8_adj_1556 : std_logic;
signal n7_adj_1555 : std_logic;
signal \data_index_9_N_212_9\ : std_logic;
signal \INVcomm_spi.MISO_48_12291_12292_resetC_net\ : std_logic;
signal \comm_spi.n14818\ : std_logic;
signal \comm_spi.n14819\ : std_logic;
signal \INVcomm_spi.MISO_48_12291_12292_setC_net\ : std_logic;
signal buf_data_iac_21 : std_logic;
signal n21672 : std_logic;
signal \ADC_VDC.n22124_cascade_\ : std_logic;
signal \VDC_SCLK\ : std_logic;
signal \VDC_CLK\ : std_logic;
signal buf_data_iac_20 : std_logic;
signal n21557 : std_logic;
signal flagcntwd : std_logic;
signal \n21187_cascade_\ : std_logic;
signal n11605 : std_logic;
signal n20578 : std_logic;
signal \n11576_cascade_\ : std_logic;
signal n12148 : std_logic;
signal n11910 : std_logic;
signal buf_data_iac_10 : std_logic;
signal n21385 : std_logic;
signal comm_buf_0_7 : std_logic;
signal n21276 : std_logic;
signal \n22542_cascade_\ : std_logic;
signal n4_adj_1580 : std_logic;
signal \comm_spi.data_tx_7__N_814\ : std_logic;
signal comm_tx_buf_7 : std_logic;
signal \comm_spi.data_tx_7__N_806\ : std_logic;
signal \comm_spi.bit_cnt_3\ : std_logic;
signal \comm_spi.n17254\ : std_logic;
signal \INVcomm_spi.data_valid_85C_net\ : std_logic;
signal \n22551_cascade_\ : std_logic;
signal comm_buf_1_4 : std_logic;
signal \n4_adj_1582_cascade_\ : std_logic;
signal \n21285_cascade_\ : std_logic;
signal n22554 : std_logic;
signal \n21474_cascade_\ : std_logic;
signal \n12_adj_1596_cascade_\ : std_logic;
signal data_idxvec_9 : std_logic;
signal data_cntvec_9 : std_logic;
signal buf_data_iac_17 : std_logic;
signal \n26_adj_1694_cascade_\ : std_logic;
signal eis_stop : std_logic;
signal req_data_cnt_9 : std_logic;
signal \acadc_skipCount_9\ : std_logic;
signal \DDS_RNG_0\ : std_logic;
signal \n22617_cascade_\ : std_logic;
signal \n22620_cascade_\ : std_logic;
signal n21360 : std_logic;
signal n22410 : std_logic;
signal \n21361_cascade_\ : std_logic;
signal \n30_adj_1695_cascade_\ : std_logic;
signal n12184 : std_logic;
signal n14958 : std_logic;
signal n22539 : std_logic;
signal n14_adj_1541 : std_logic;
signal buf_data_iac_0 : std_logic;
signal n22_adj_1532 : std_logic;
signal n21586 : std_logic;
signal comm_buf_6_7 : std_logic;
signal \acadc_skipCount_6\ : std_logic;
signal req_data_cnt_6 : std_logic;
signal n19_adj_1625 : std_logic;
signal \buf_readRTD_6\ : std_logic;
signal data_idxvec_6 : std_logic;
signal data_cntvec_6 : std_logic;
signal \n26_adj_1626_cascade_\ : std_logic;
signal n22515 : std_logic;
signal n16_adj_1624 : std_logic;
signal buf_adcdata_iac_14 : std_logic;
signal n22527 : std_logic;
signal \n22530_cascade_\ : std_logic;
signal n22518 : std_logic;
signal \n30_adj_1627_cascade_\ : std_logic;
signal data_idxvec_0 : std_logic;
signal data_cntvec_0 : std_logic;
signal buf_data_iac_8 : std_logic;
signal \n26_cascade_\ : std_logic;
signal \n21261_cascade_\ : std_logic;
signal \n22563_cascade_\ : std_logic;
signal n21257 : std_logic;
signal \n22566_cascade_\ : std_logic;
signal buf_adcdata_vdc_8 : std_logic;
signal buf_adcdata_vac_8 : std_logic;
signal \buf_readRTD_0\ : std_logic;
signal \n19_cascade_\ : std_logic;
signal n21258 : std_logic;
signal \acadc_skipCount_0\ : std_logic;
signal req_data_cnt_0 : std_logic;
signal n21260 : std_logic;
signal buf_adcdata_iac_9 : std_logic;
signal n16_adj_1651 : std_logic;
signal n22431 : std_logic;
signal data_idxvec_1 : std_logic;
signal data_cntvec_1 : std_logic;
signal \n26_adj_1653_cascade_\ : std_logic;
signal \acadc_skipCount_1\ : std_logic;
signal \n22497_cascade_\ : std_logic;
signal req_data_cnt_1 : std_logic;
signal n22434 : std_logic;
signal \n22500_cascade_\ : std_logic;
signal \n30_adj_1654_cascade_\ : std_logic;
signal n28 : std_logic;
signal comm_buf_1_7 : std_logic;
signal n14965 : std_logic;
signal trig_dds0 : std_logic;
signal \SIG_DDS.n12895\ : std_logic;
signal wdtick_flag : std_logic;
signal buf_control_0 : std_logic;
signal \CONT_SD\ : std_logic;
signal dds_state_0 : std_logic;
signal dds_state_2 : std_logic;
signal \SIG_DDS.n9\ : std_logic;
signal dds_state_1 : std_logic;
signal \comm_spi.n14813\ : std_logic;
signal \comm_spi.n14812\ : std_logic;
signal \comm_spi.n14811\ : std_logic;
signal \ICE_SPI_MISO\ : std_logic;
signal \ADC_VDC.n11895\ : std_logic;
signal \comm_spi.n23086\ : std_logic;
signal \comm_spi.n23086_cascade_\ : std_logic;
signal \comm_spi.n14804\ : std_logic;
signal n80 : std_logic;
signal n5 : std_logic;
signal \comm_spi.n23092\ : std_logic;
signal clk_cnt_1 : std_logic;
signal clk_cnt_0 : std_logic;
signal n17773 : std_logic;
signal buf_data_vac_8 : std_logic;
signal buf_data_vac_15 : std_logic;
signal comm_buf_4_7 : std_logic;
signal buf_data_vac_14 : std_logic;
signal buf_data_vac_13 : std_logic;
signal buf_data_vac_12 : std_logic;
signal comm_buf_4_4 : std_logic;
signal buf_data_vac_11 : std_logic;
signal buf_data_vac_10 : std_logic;
signal buf_data_vac_9 : std_logic;
signal n14986 : std_logic;
signal \n21268_cascade_\ : std_logic;
signal n22094 : std_logic;
signal n21266 : std_logic;
signal n12407 : std_logic;
signal \n21085_cascade_\ : std_logic;
signal n19188 : std_logic;
signal \n19188_cascade_\ : std_logic;
signal comm_buf_0_3 : std_logic;
signal \n22557_cascade_\ : std_logic;
signal comm_buf_1_3 : std_logic;
signal comm_buf_4_3 : std_logic;
signal \n4_adj_1583_cascade_\ : std_logic;
signal n22560 : std_logic;
signal \n21288_cascade_\ : std_logic;
signal n21479 : std_logic;
signal \n21477_cascade_\ : std_logic;
signal \n44_cascade_\ : std_logic;
signal n12260 : std_logic;
signal comm_buf_1_2 : std_logic;
signal \n1_cascade_\ : std_logic;
signal n2_adj_1584 : std_logic;
signal comm_buf_4_2 : std_logic;
signal n21528 : std_logic;
signal \n4_adj_1585_cascade_\ : std_logic;
signal n22491 : std_logic;
signal n21143 : std_logic;
signal \n19193_cascade_\ : std_logic;
signal n21273 : std_logic;
signal comm_buf_1_0 : std_logic;
signal \n22533_cascade_\ : std_logic;
signal comm_buf_0_0 : std_logic;
signal n22536 : std_logic;
signal n24_adj_1639 : std_logic;
signal \n21497_cascade_\ : std_logic;
signal \n34_adj_1649_cascade_\ : std_logic;
signal n30_adj_1531 : std_logic;
signal comm_buf_2_0 : std_logic;
signal n30_adj_1599 : std_logic;
signal comm_buf_2_7 : std_logic;
signal n30_adj_1602 : std_logic;
signal n30_adj_1605 : std_logic;
signal n30_adj_1608 : std_logic;
signal comm_buf_2_4 : std_logic;
signal n30_adj_1611 : std_logic;
signal comm_buf_2_3 : std_logic;
signal n30_adj_1614 : std_logic;
signal comm_buf_2_2 : std_logic;
signal n30_adj_1618 : std_logic;
signal n12314 : std_logic;
signal n14972 : std_logic;
signal comm_buf_0_2 : std_logic;
signal buf_data_iac_19 : std_logic;
signal n21543 : std_logic;
signal \SELIRNG0\ : std_logic;
signal n23_adj_1685 : std_logic;
signal comm_buf_6_0 : std_logic;
signal comm_buf_6_3 : std_logic;
signal \acadc_skipCount_7\ : std_logic;
signal req_data_cnt_7 : std_logic;
signal data_idxvec_7 : std_logic;
signal data_cntvec_7 : std_logic;
signal buf_data_iac_15 : std_logic;
signal \n26_adj_1622_cascade_\ : std_logic;
signal comm_cmd_1 : std_logic;
signal n16824 : std_logic;
signal comm_length_1 : std_logic;
signal n5_adj_1524 : std_logic;
signal n12654 : std_logic;
signal comm_buf_0_4 : std_logic;
signal comm_cmd_2 : std_logic;
signal n21368 : std_logic;
signal n21369 : std_logic;
signal n21362 : std_logic;
signal n21363 : std_logic;
signal \n22599_cascade_\ : std_logic;
signal comm_cmd_3 : std_logic;
signal n22602 : std_logic;
signal buf_dds1_6 : std_logic;
signal n68 : std_logic;
signal n12048 : std_logic;
signal \n12048_cascade_\ : std_logic;
signal n16971 : std_logic;
signal \comm_spi.n14805\ : std_logic;
signal \comm_spi.iclk_N_802\ : std_logic;
signal \ICE_SPI_SCLK\ : std_logic;
signal \comm_spi.iclk_N_803\ : std_logic;
signal buf_data_vac_0 : std_logic;
signal buf_data_vac_7 : std_logic;
signal comm_buf_5_7 : std_logic;
signal buf_data_vac_6 : std_logic;
signal buf_data_vac_5 : std_logic;
signal buf_data_vac_4 : std_logic;
signal comm_buf_5_4 : std_logic;
signal buf_data_vac_3 : std_logic;
signal comm_buf_5_3 : std_logic;
signal buf_data_vac_2 : std_logic;
signal comm_buf_5_2 : std_logic;
signal buf_data_vac_1 : std_logic;
signal n12431 : std_logic;
signal n14993 : std_logic;
signal n11652 : std_logic;
signal \n2_adj_1576_cascade_\ : std_logic;
signal n22611 : std_logic;
signal \comm_state_3_N_460_3\ : std_logic;
signal \n1348_cascade_\ : std_logic;
signal \n21139_cascade_\ : std_logic;
signal n1348 : std_logic;
signal n8_adj_1577 : std_logic;
signal n22614 : std_logic;
signal n4 : std_logic;
signal \n21013_cascade_\ : std_logic;
signal n21035 : std_logic;
signal comm_length_0 : std_logic;
signal n4_adj_1623 : std_logic;
signal n3 : std_logic;
signal n21110 : std_logic;
signal \n3_cascade_\ : std_logic;
signal n12442 : std_logic;
signal n4_adj_1589 : std_logic;
signal \n20095_cascade_\ : std_logic;
signal n21013 : std_logic;
signal n11619 : std_logic;
signal n21588 : std_logic;
signal n9342 : std_logic;
signal n18070 : std_logic;
signal n21033 : std_logic;
signal n7_adj_1650 : std_logic;
signal comm_cmd_6 : std_logic;
signal comm_cmd_5 : std_logic;
signal n4_adj_1455 : std_logic;
signal n21147 : std_logic;
signal \n21219_cascade_\ : std_logic;
signal n21089 : std_logic;
signal n21043 : std_logic;
signal buf_data_vac_16 : std_logic;
signal comm_rx_buf_0 : std_logic;
signal comm_buf_3_0 : std_logic;
signal buf_data_vac_23 : std_logic;
signal comm_rx_buf_7 : std_logic;
signal comm_buf_3_7 : std_logic;
signal buf_data_vac_22 : std_logic;
signal buf_data_vac_21 : std_logic;
signal buf_data_vac_20 : std_logic;
signal comm_buf_3_4 : std_logic;
signal comm_rx_buf_3 : std_logic;
signal buf_data_vac_19 : std_logic;
signal comm_buf_3_3 : std_logic;
signal buf_data_vac_18 : std_logic;
signal comm_buf_3_2 : std_logic;
signal comm_rx_buf_1 : std_logic;
signal buf_data_vac_17 : std_logic;
signal comm_buf_5_6 : std_logic;
signal comm_buf_4_6 : std_logic;
signal comm_buf_2_6 : std_logic;
signal comm_buf_3_6 : std_logic;
signal comm_buf_0_6 : std_logic;
signal \n22545_cascade_\ : std_logic;
signal comm_buf_1_6 : std_logic;
signal n12353 : std_logic;
signal n14979 : std_logic;
signal comm_rx_buf_2 : std_logic;
signal comm_buf_6_2 : std_logic;
signal comm_buf_5_0 : std_logic;
signal comm_buf_4_0 : std_logic;
signal n4_adj_1457 : std_logic;
signal comm_buf_5_1 : std_logic;
signal comm_buf_4_1 : std_logic;
signal comm_cmd_7 : std_logic;
signal comm_buf_6_1 : std_logic;
signal n4_adj_1588 : std_logic;
signal \n21433_cascade_\ : std_logic;
signal \n22419_cascade_\ : std_logic;
signal n21085 : std_logic;
signal \n7_adj_1458_cascade_\ : std_logic;
signal n4_adj_1581 : std_logic;
signal \n21282_cascade_\ : std_logic;
signal n22548 : std_logic;
signal comm_tx_buf_6 : std_logic;
signal comm_buf_5_5 : std_logic;
signal comm_buf_1_5 : std_logic;
signal comm_buf_3_5 : std_logic;
signal \n17698_cascade_\ : std_logic;
signal \n21270_cascade_\ : std_logic;
signal n12541 : std_logic;
signal n15007 : std_logic;
signal \n20996_cascade_\ : std_logic;
signal n12_adj_1663 : std_logic;
signal n20996 : std_logic;
signal \INVdds0_mclk_294C_net\ : std_logic;
signal \clk_16MHz\ : std_logic;
signal dds0_mclk : std_logic;
signal buf_control_6 : std_logic;
signal \DDS_MCLK\ : std_logic;
signal acadc_skipcnt_10 : std_logic;
signal \acadc_skipCount_12\ : std_logic;
signal acadc_skipcnt_12 : std_logic;
signal \acadc_skipCount_10\ : std_logic;
signal n21 : std_logic;
signal n11590 : std_logic;
signal dds0_mclkcnt_0 : std_logic;
signal \bfn_18_16_0_\ : std_logic;
signal dds0_mclkcnt_1 : std_logic;
signal n19925 : std_logic;
signal dds0_mclkcnt_2 : std_logic;
signal n19926 : std_logic;
signal dds0_mclkcnt_3 : std_logic;
signal n19927 : std_logic;
signal dds0_mclkcnt_4 : std_logic;
signal n19928 : std_logic;
signal dds0_mclkcnt_5 : std_logic;
signal n19929 : std_logic;
signal n10_adj_1528 : std_logic;
signal dds0_mclkcnt_6 : std_logic;
signal n19930 : std_logic;
signal n19931 : std_logic;
signal dds0_mclkcnt_7 : std_logic;
signal \INVdds0_mclkcnt_i7_3772__i0C_net\ : std_logic;
signal n14716 : std_logic;
signal \ICE_SPI_MOSI\ : std_logic;
signal \comm_spi.imosi_N_793\ : std_logic;
signal \comm_spi.data_tx_7__N_810\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i1C_net\ : std_logic;
signal \VDC_SDO\ : std_logic;
signal \ADC_VDC.adc_state_0\ : std_logic;
signal adc_state_3 : std_logic;
signal adc_state_2_adj_1500 : std_logic;
signal \ADC_VDC.n52_cascade_\ : std_logic;
signal \ADC_VDC.adc_state_1\ : std_logic;
signal \ADC_VDC.n11905\ : std_logic;
signal \bfn_19_7_0_\ : std_logic;
signal \ADC_VDC.genclk.n19888\ : std_logic;
signal \ADC_VDC.genclk.n19889\ : std_logic;
signal \ADC_VDC.genclk.n19890\ : std_logic;
signal \ADC_VDC.genclk.n19891\ : std_logic;
signal \ADC_VDC.genclk.n19892\ : std_logic;
signal \ADC_VDC.genclk.n19893\ : std_logic;
signal \ADC_VDC.genclk.n19894\ : std_logic;
signal \ADC_VDC.genclk.n19895\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i0C_net\ : std_logic;
signal \bfn_19_8_0_\ : std_logic;
signal \ADC_VDC.genclk.n19896\ : std_logic;
signal \ADC_VDC.genclk.n19897\ : std_logic;
signal \ADC_VDC.genclk.n19898\ : std_logic;
signal \ADC_VDC.genclk.n19899\ : std_logic;
signal \ADC_VDC.genclk.n19900\ : std_logic;
signal \ADC_VDC.genclk.n19901\ : std_logic;
signal \ADC_VDC.genclk.n19902\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.n11900\ : std_logic;
signal n14350 : std_logic;
signal n21453 : std_logic;
signal \n21454_cascade_\ : std_logic;
signal n14_adj_1638 : std_logic;
signal n21481 : std_logic;
signal n12089 : std_logic;
signal comm_length_2 : std_logic;
signal n6541 : std_logic;
signal n21154 : std_logic;
signal comm_data_vld : std_logic;
signal \ICE_SPI_CE0\ : std_logic;
signal n6401 : std_logic;
signal n16821 : std_logic;
signal \comm_spi.n14842\ : std_logic;
signal buf_data_iac_18 : std_logic;
signal n21460 : std_logic;
signal comm_buf_2_5 : std_logic;
signal comm_index_2 : std_logic;
signal comm_index_1 : std_logic;
signal comm_buf_0_5 : std_logic;
signal \n22503_cascade_\ : std_logic;
signal comm_buf_4_5 : std_logic;
signal n22506 : std_logic;
signal comm_tx_buf_5 : std_logic;
signal \comm_spi.data_tx_7__N_808\ : std_logic;
signal comm_rx_buf_4 : std_logic;
signal comm_buf_6_4 : std_logic;
signal comm_buf_3_1 : std_logic;
signal comm_buf_2_1 : std_logic;
signal n2_adj_1587 : std_logic;
signal comm_buf_1_1 : std_logic;
signal comm_buf_0_1 : std_logic;
signal n1_adj_1586 : std_logic;
signal comm_rx_buf_5 : std_logic;
signal comm_buf_6_5 : std_logic;
signal buf_data_iac_14 : std_logic;
signal n21547 : std_logic;
signal comm_rx_buf_6 : std_logic;
signal n12477 : std_logic;
signal comm_buf_6_6 : std_logic;
signal comm_index_0 : std_logic;
signal n8_adj_1456 : std_logic;
signal comm_tx_buf_3 : std_logic;
signal \ICE_GPMI_0\ : std_logic;
signal \clk_32MHz\ : std_logic;
signal n11600 : std_logic;
signal n12433 : std_logic;
signal \n10_adj_1619_cascade_\ : std_logic;
signal comm_state_3 : std_logic;
signal n12079 : std_logic;
signal comm_state_2 : std_logic;
signal comm_state_1 : std_logic;
signal comm_state_0 : std_logic;
signal n10804 : std_logic;
signal \ADC_VDC.genclk.t0off_12\ : std_logic;
signal \ADC_VDC.genclk.t0off_2\ : std_logic;
signal \ADC_VDC.genclk.t0off_7\ : std_logic;
signal \ADC_VDC.genclk.t0off_10\ : std_logic;
signal \ADC_VDC.genclk.n27_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n21598_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n6\ : std_logic;
signal \ADC_VDC.genclk.t0off_6\ : std_logic;
signal \ADC_VDC.genclk.t0off_1\ : std_logic;
signal \ADC_VDC.genclk.t0off_4\ : std_logic;
signal \ADC_VDC.genclk.t0off_0\ : std_logic;
signal \ADC_VDC.genclk.n21600\ : std_logic;
signal \ADC_VDC.genclk.n27_adj_1449_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n21597\ : std_logic;
signal \ADC_VDC.genclk.n21598\ : std_logic;
signal \ADC_VDC.genclk.n21597_cascade_\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.n21603\ : std_logic;
signal \ADC_VDC.genclk.t0off_13\ : std_logic;
signal \ADC_VDC.genclk.t0off_3\ : std_logic;
signal \ADC_VDC.genclk.t0off_5\ : std_logic;
signal \ADC_VDC.genclk.t0off_8\ : std_logic;
signal \ADC_VDC.genclk.n26\ : std_logic;
signal \ADC_VDC.genclk.div_state_0\ : std_logic;
signal \ADC_VDC.genclk.n28_adj_1447\ : std_logic;
signal \ADC_VDC.genclk.t0off_14\ : std_logic;
signal \ADC_VDC.genclk.t0off_9\ : std_logic;
signal \ADC_VDC.genclk.t0off_15\ : std_logic;
signal \ADC_VDC.genclk.t0off_11\ : std_logic;
signal \ADC_VDC.genclk.n28\ : std_logic;
signal \ADC_VDC.genclk.n26_adj_1448\ : std_logic;
signal \comm_spi.n23101\ : std_logic;
signal \comm_spi.n14834\ : std_logic;
signal \comm_spi.data_tx_7__N_823\ : std_logic;
signal \comm_spi.data_tx_7__N_811\ : std_logic;
signal comm_tx_buf_4 : std_logic;
signal \comm_spi.data_tx_7__N_809\ : std_logic;
signal comm_tx_buf_2 : std_logic;
signal \comm_spi.data_tx_7__N_829\ : std_logic;
signal \comm_spi.n23098\ : std_logic;
signal \comm_spi.n14838\ : std_logic;
signal \comm_spi.n14839\ : std_logic;
signal \comm_spi.n14843\ : std_logic;
signal \comm_spi.data_tx_7__N_820\ : std_logic;
signal \comm_spi.n23104\ : std_logic;
signal \comm_spi.n14830\ : std_logic;
signal \comm_spi.n14831\ : std_logic;
signal \comm_spi.n14835\ : std_logic;
signal \comm_spi.data_tx_7__N_826\ : std_logic;
signal buf_data_iac_13 : std_logic;
signal n21456 : std_logic;
signal buf_data_iac_12 : std_logic;
signal n21447 : std_logic;
signal buf_data_iac_9 : std_logic;
signal n21512 : std_logic;
signal buf_data_iac_11 : std_logic;
signal comm_cmd_0 : std_logic;
signal n21434 : std_logic;
signal \ADC_VDC.genclk.div_state_1\ : std_logic;
signal \ADC_VDC.genclk.t0on_0\ : std_logic;
signal \bfn_22_7_0_\ : std_logic;
signal \ADC_VDC.genclk.t0on_1\ : std_logic;
signal \ADC_VDC.genclk.n19903\ : std_logic;
signal \ADC_VDC.genclk.t0on_2\ : std_logic;
signal \ADC_VDC.genclk.n19904\ : std_logic;
signal \ADC_VDC.genclk.t0on_3\ : std_logic;
signal \ADC_VDC.genclk.n19905\ : std_logic;
signal \ADC_VDC.genclk.t0on_4\ : std_logic;
signal \ADC_VDC.genclk.n19906\ : std_logic;
signal \ADC_VDC.genclk.t0on_5\ : std_logic;
signal \ADC_VDC.genclk.n19907\ : std_logic;
signal \ADC_VDC.genclk.t0on_6\ : std_logic;
signal \ADC_VDC.genclk.n19908\ : std_logic;
signal \ADC_VDC.genclk.t0on_7\ : std_logic;
signal \ADC_VDC.genclk.n19909\ : std_logic;
signal \ADC_VDC.genclk.n19910\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.t0on_8\ : std_logic;
signal \bfn_22_8_0_\ : std_logic;
signal \ADC_VDC.genclk.t0on_9\ : std_logic;
signal \ADC_VDC.genclk.n19911\ : std_logic;
signal \ADC_VDC.genclk.t0on_10\ : std_logic;
signal \ADC_VDC.genclk.n19912\ : std_logic;
signal \ADC_VDC.genclk.t0on_11\ : std_logic;
signal \ADC_VDC.genclk.n19913\ : std_logic;
signal \ADC_VDC.genclk.t0on_12\ : std_logic;
signal \ADC_VDC.genclk.n19914\ : std_logic;
signal \ADC_VDC.genclk.t0on_13\ : std_logic;
signal \ADC_VDC.genclk.n19915\ : std_logic;
signal \ADC_VDC.genclk.t0on_14\ : std_logic;
signal \ADC_VDC.genclk.n19916\ : std_logic;
signal \ADC_VDC.genclk.n19917\ : std_logic;
signal \ADC_VDC.genclk.t0on_15\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.div_state_1__N_1432\ : std_logic;
signal \ADC_VDC.genclk.n14894\ : std_logic;
signal \comm_spi.data_tx_7__N_835\ : std_logic;
signal \comm_spi.n14827\ : std_logic;
signal \comm_spi.n23110\ : std_logic;
signal \comm_spi.n14801\ : std_logic;
signal \comm_spi.n14826\ : std_logic;
signal \comm_spi.data_tx_7__N_812\ : std_logic;
signal \comm_spi.data_tx_7__N_832\ : std_logic;
signal comm_tx_buf_1 : std_logic;
signal \comm_spi.n23107\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \comm_spi.n14800\ : std_logic;
signal \comm_spi.iclk\ : std_logic;
signal comm_tx_buf_0 : std_logic;
signal comm_clear : std_logic;
signal \comm_spi.data_tx_7__N_813\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VAC_DRDY_wire\ : std_logic;
signal \IAC_FLT1_wire\ : std_logic;
signal \DDS_SCK_wire\ : std_logic;
signal \ICE_IOR_166_wire\ : std_logic;
signal \ICE_IOR_119_wire\ : std_logic;
signal \DDS_MOSI_wire\ : std_logic;
signal \VAC_MISO_wire\ : std_logic;
signal \DDS_MOSI1_wire\ : std_logic;
signal \ICE_IOR_146_wire\ : std_logic;
signal \VDC_CLK_wire\ : std_logic;
signal \ICE_IOT_222_wire\ : std_logic;
signal \IAC_CS_wire\ : std_logic;
signal \ICE_IOL_18B_wire\ : std_logic;
signal \ICE_IOL_13A_wire\ : std_logic;
signal \ICE_IOB_81_wire\ : std_logic;
signal \VAC_OSR1_wire\ : std_logic;
signal \IAC_MOSI_wire\ : std_logic;
signal \DDS_CS1_wire\ : std_logic;
signal \ICE_IOL_4B_wire\ : std_logic;
signal \ICE_IOB_94_wire\ : std_logic;
signal \VAC_CS_wire\ : std_logic;
signal \VAC_CLK_wire\ : std_logic;
signal \ICE_SPI_CE0_wire\ : std_logic;
signal \ICE_IOR_167_wire\ : std_logic;
signal \ICE_IOR_118_wire\ : std_logic;
signal \RTD_SDO_wire\ : std_logic;
signal \IAC_OSR0_wire\ : std_logic;
signal \VDC_SCLK_wire\ : std_logic;
signal \VAC_FLT1_wire\ : std_logic;
signal \ICE_SPI_MOSI_wire\ : std_logic;
signal \ICE_IOR_165_wire\ : std_logic;
signal \ICE_IOR_147_wire\ : std_logic;
signal \ICE_IOL_14A_wire\ : std_logic;
signal \ICE_IOL_13B_wire\ : std_logic;
signal \ICE_IOB_91_wire\ : std_logic;
signal \ICE_GPMO_0_wire\ : std_logic;
signal \DDS_RNG_0_wire\ : std_logic;
signal \VDC_RNG0_wire\ : std_logic;
signal \ICE_SPI_SCLK_wire\ : std_logic;
signal \ICE_IOR_152_wire\ : std_logic;
signal \ICE_IOL_12A_wire\ : std_logic;
signal \RTD_DRDY_wire\ : std_logic;
signal \ICE_SPI_MISO_wire\ : std_logic;
signal \ICE_IOT_177_wire\ : std_logic;
signal \ICE_IOR_141_wire\ : std_logic;
signal \ICE_IOB_80_wire\ : std_logic;
signal \ICE_IOB_102_wire\ : std_logic;
signal \ICE_GPMO_2_wire\ : std_logic;
signal \ICE_GPMI_0_wire\ : std_logic;
signal \IAC_MISO_wire\ : std_logic;
signal \VAC_OSR0_wire\ : std_logic;
signal \VAC_MOSI_wire\ : std_logic;
signal \TEST_LED_wire\ : std_logic;
signal \ICE_IOR_148_wire\ : std_logic;
signal \STAT_COMM_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \ICE_IOR_161_wire\ : std_logic;
signal \ICE_IOB_95_wire\ : std_logic;
signal \ICE_IOB_82_wire\ : std_logic;
signal \ICE_IOB_104_wire\ : std_logic;
signal \IAC_CLK_wire\ : std_logic;
signal \DDS_CS_wire\ : std_logic;
signal \SELIRNG0_wire\ : std_logic;
signal \RTD_SDI_wire\ : std_logic;
signal \ICE_IOT_221_wire\ : std_logic;
signal \ICE_IOT_197_wire\ : std_logic;
signal \DDS_MCLK_wire\ : std_logic;
signal \RTD_SCLK_wire\ : std_logic;
signal \RTD_CS_wire\ : std_logic;
signal \ICE_IOR_137_wire\ : std_logic;
signal \IAC_OSR1_wire\ : std_logic;
signal \VAC_FLT0_wire\ : std_logic;
signal \ICE_IOR_144_wire\ : std_logic;
signal \ICE_IOR_128_wire\ : std_logic;
signal \ICE_GPMO_1_wire\ : std_logic;
signal \IAC_SCLK_wire\ : std_logic;
signal \EIS_SYNCCLK_wire\ : std_logic;
signal \ICE_IOR_139_wire\ : std_logic;
signal \ICE_IOL_4A_wire\ : std_logic;
signal \VAC_SCLK_wire\ : std_logic;
signal \THERMOSTAT_wire\ : std_logic;
signal \ICE_IOR_164_wire\ : std_logic;
signal \ICE_IOB_103_wire\ : std_logic;
signal \AMPV_POW_wire\ : std_logic;
signal \VDC_SDO_wire\ : std_logic;
signal \ICE_IOT_174_wire\ : std_logic;
signal \ICE_IOR_140_wire\ : std_logic;
signal \ICE_IOB_96_wire\ : std_logic;
signal \CONT_SD_wire\ : std_logic;
signal \AC_ADC_SYNC_wire\ : std_logic;
signal \SELIRNG1_wire\ : std_logic;
signal \ICE_IOL_12B_wire\ : std_logic;
signal \ICE_IOR_160_wire\ : std_logic;
signal \ICE_IOR_136_wire\ : std_logic;
signal \DDS_MCLK1_wire\ : std_logic;
signal \ICE_IOT_198_wire\ : std_logic;
signal \ICE_IOT_173_wire\ : std_logic;
signal \IAC_DRDY_wire\ : std_logic;
signal \ICE_IOT_178_wire\ : std_logic;
signal \ICE_IOR_138_wire\ : std_logic;
signal \ICE_IOR_120_wire\ : std_logic;
signal \IAC_FLT0_wire\ : std_logic;
signal \DDS_SCK1_wire\ : std_logic;
signal \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \VAC_DRDY_wire\ <= VAC_DRDY;
    IAC_FLT1 <= \IAC_FLT1_wire\;
    DDS_SCK <= \DDS_SCK_wire\;
    \ICE_IOR_166_wire\ <= ICE_IOR_166;
    \ICE_IOR_119_wire\ <= ICE_IOR_119;
    DDS_MOSI <= \DDS_MOSI_wire\;
    \VAC_MISO_wire\ <= VAC_MISO;
    DDS_MOSI1 <= \DDS_MOSI1_wire\;
    \ICE_IOR_146_wire\ <= ICE_IOR_146;
    VDC_CLK <= \VDC_CLK_wire\;
    \ICE_IOT_222_wire\ <= ICE_IOT_222;
    IAC_CS <= \IAC_CS_wire\;
    \ICE_IOL_18B_wire\ <= ICE_IOL_18B;
    \ICE_IOL_13A_wire\ <= ICE_IOL_13A;
    \ICE_IOB_81_wire\ <= ICE_IOB_81;
    VAC_OSR1 <= \VAC_OSR1_wire\;
    IAC_MOSI <= \IAC_MOSI_wire\;
    DDS_CS1 <= \DDS_CS1_wire\;
    \ICE_IOL_4B_wire\ <= ICE_IOL_4B;
    \ICE_IOB_94_wire\ <= ICE_IOB_94;
    VAC_CS <= \VAC_CS_wire\;
    VAC_CLK <= \VAC_CLK_wire\;
    \ICE_SPI_CE0_wire\ <= ICE_SPI_CE0;
    \ICE_IOR_167_wire\ <= ICE_IOR_167;
    \ICE_IOR_118_wire\ <= ICE_IOR_118;
    \RTD_SDO_wire\ <= RTD_SDO;
    IAC_OSR0 <= \IAC_OSR0_wire\;
    VDC_SCLK <= \VDC_SCLK_wire\;
    VAC_FLT1 <= \VAC_FLT1_wire\;
    \ICE_SPI_MOSI_wire\ <= ICE_SPI_MOSI;
    \ICE_IOR_165_wire\ <= ICE_IOR_165;
    \ICE_IOR_147_wire\ <= ICE_IOR_147;
    \ICE_IOL_14A_wire\ <= ICE_IOL_14A;
    \ICE_IOL_13B_wire\ <= ICE_IOL_13B;
    \ICE_IOB_91_wire\ <= ICE_IOB_91;
    \ICE_GPMO_0_wire\ <= ICE_GPMO_0;
    DDS_RNG_0 <= \DDS_RNG_0_wire\;
    VDC_RNG0 <= \VDC_RNG0_wire\;
    \ICE_SPI_SCLK_wire\ <= ICE_SPI_SCLK;
    \ICE_IOR_152_wire\ <= ICE_IOR_152;
    \ICE_IOL_12A_wire\ <= ICE_IOL_12A;
    \RTD_DRDY_wire\ <= RTD_DRDY;
    ICE_SPI_MISO <= \ICE_SPI_MISO_wire\;
    \ICE_IOT_177_wire\ <= ICE_IOT_177;
    \ICE_IOR_141_wire\ <= ICE_IOR_141;
    \ICE_IOB_80_wire\ <= ICE_IOB_80;
    \ICE_IOB_102_wire\ <= ICE_IOB_102;
    \ICE_GPMO_2_wire\ <= ICE_GPMO_2;
    ICE_GPMI_0 <= \ICE_GPMI_0_wire\;
    \IAC_MISO_wire\ <= IAC_MISO;
    VAC_OSR0 <= \VAC_OSR0_wire\;
    VAC_MOSI <= \VAC_MOSI_wire\;
    TEST_LED <= \TEST_LED_wire\;
    \ICE_IOR_148_wire\ <= ICE_IOR_148;
    STAT_COMM <= \STAT_COMM_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    \ICE_IOR_161_wire\ <= ICE_IOR_161;
    \ICE_IOB_95_wire\ <= ICE_IOB_95;
    \ICE_IOB_82_wire\ <= ICE_IOB_82;
    \ICE_IOB_104_wire\ <= ICE_IOB_104;
    IAC_CLK <= \IAC_CLK_wire\;
    DDS_CS <= \DDS_CS_wire\;
    SELIRNG0 <= \SELIRNG0_wire\;
    RTD_SDI <= \RTD_SDI_wire\;
    \ICE_IOT_221_wire\ <= ICE_IOT_221;
    \ICE_IOT_197_wire\ <= ICE_IOT_197;
    DDS_MCLK <= \DDS_MCLK_wire\;
    RTD_SCLK <= \RTD_SCLK_wire\;
    RTD_CS <= \RTD_CS_wire\;
    \ICE_IOR_137_wire\ <= ICE_IOR_137;
    IAC_OSR1 <= \IAC_OSR1_wire\;
    VAC_FLT0 <= \VAC_FLT0_wire\;
    \ICE_IOR_144_wire\ <= ICE_IOR_144;
    \ICE_IOR_128_wire\ <= ICE_IOR_128;
    \ICE_GPMO_1_wire\ <= ICE_GPMO_1;
    IAC_SCLK <= \IAC_SCLK_wire\;
    \EIS_SYNCCLK_wire\ <= EIS_SYNCCLK;
    \ICE_IOR_139_wire\ <= ICE_IOR_139;
    \ICE_IOL_4A_wire\ <= ICE_IOL_4A;
    VAC_SCLK <= \VAC_SCLK_wire\;
    \THERMOSTAT_wire\ <= THERMOSTAT;
    \ICE_IOR_164_wire\ <= ICE_IOR_164;
    \ICE_IOB_103_wire\ <= ICE_IOB_103;
    AMPV_POW <= \AMPV_POW_wire\;
    \VDC_SDO_wire\ <= VDC_SDO;
    \ICE_IOT_174_wire\ <= ICE_IOT_174;
    \ICE_IOR_140_wire\ <= ICE_IOR_140;
    \ICE_IOB_96_wire\ <= ICE_IOB_96;
    CONT_SD <= \CONT_SD_wire\;
    AC_ADC_SYNC <= \AC_ADC_SYNC_wire\;
    SELIRNG1 <= \SELIRNG1_wire\;
    \ICE_IOL_12B_wire\ <= ICE_IOL_12B;
    \ICE_IOR_160_wire\ <= ICE_IOR_160;
    \ICE_IOR_136_wire\ <= ICE_IOR_136;
    DDS_MCLK1 <= \DDS_MCLK1_wire\;
    \ICE_IOT_198_wire\ <= ICE_IOT_198;
    \ICE_IOT_173_wire\ <= ICE_IOT_173;
    \IAC_DRDY_wire\ <= IAC_DRDY;
    \ICE_IOT_178_wire\ <= ICE_IOT_178;
    \ICE_IOR_138_wire\ <= ICE_IOR_138;
    \ICE_IOR_120_wire\ <= ICE_IOR_120;
    IAC_FLT0 <= \IAC_FLT0_wire\;
    DDS_SCK1 <= \DDS_SCK1_wire\;
    \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    buf_data_iac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(13);
    buf_data_vac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(9);
    buf_data_iac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(5);
    buf_data_vac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ <= '0'&\N__41862\&\N__39420\&\N__32922\&\N__36093\&\N__41382\&\N__36414\&\N__35943\&\N__39879\&\N__39288\&\N__41010\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ <= '0'&\N__33885\&\N__33996\&\N__34104\&\N__34212\&\N__33198\&\N__33300\&\N__33411\&\N__33522\&\N__33630\&\N__33732\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ <= '0'&'0'&\N__26472\&'0'&'0'&'0'&\N__25980\&'0'&'0'&'0'&\N__32763\&'0'&'0'&'0'&\N__24138\&'0';
    buf_data_iac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(13);
    buf_data_vac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(9);
    buf_data_iac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(5);
    buf_data_vac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ <= '0'&\N__41822\&\N__39380\&\N__32885\&\N__36047\&\N__41336\&\N__36377\&\N__35906\&\N__39836\&\N__39245\&\N__40967\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ <= '0'&\N__33848\&\N__33956\&\N__34058\&\N__34172\&\N__33155\&\N__33266\&\N__33374\&\N__33485\&\N__33590\&\N__33692\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ <= '0'&'0'&\N__43620\&'0'&'0'&'0'&\N__23568\&'0'&'0'&'0'&\N__41706\&'0'&'0'&'0'&\N__43758\&'0';
    buf_data_iac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(13);
    buf_data_vac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(9);
    buf_data_iac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(5);
    buf_data_vac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ <= '0'&\N__41880\&\N__39438\&\N__32940\&\N__36111\&\N__41400\&\N__36432\&\N__35961\&\N__39897\&\N__39306\&\N__41028\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ <= '0'&\N__33903\&\N__34014\&\N__34122\&\N__34230\&\N__33216\&\N__33318\&\N__33429\&\N__33540\&\N__33648\&\N__33750\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ <= '0'&'0'&\N__28947\&'0'&'0'&'0'&\N__27429\&'0'&'0'&'0'&\N__32148\&'0'&'0'&'0'&\N__31884\&'0';
    buf_data_iac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(13);
    buf_data_vac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(9);
    buf_data_iac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(5);
    buf_data_vac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ <= '0'&\N__41834\&\N__39392\&\N__32897\&\N__36059\&\N__41348\&\N__36389\&\N__35918\&\N__39848\&\N__39257\&\N__40979\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ <= '0'&\N__33860\&\N__33968\&\N__34070\&\N__34184\&\N__33167\&\N__33276\&\N__33386\&\N__33497\&\N__33602\&\N__33704\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ <= '0'&'0'&\N__41303\&'0'&'0'&'0'&\N__35052\&'0'&'0'&'0'&\N__38237\&'0'&'0'&'0'&\N__27333\&'0';
    buf_data_iac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(13);
    buf_data_vac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(9);
    buf_data_iac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(5);
    buf_data_vac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ <= '0'&\N__41886\&\N__39444\&\N__32946\&\N__36117\&\N__41406\&\N__36438\&\N__35967\&\N__39903\&\N__39312\&\N__41034\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ <= '0'&\N__33909\&\N__34020\&\N__34128\&\N__34236\&\N__33222\&\N__33324\&\N__33435\&\N__33546\&\N__33654\&\N__33756\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ <= '0'&'0'&\N__29201\&'0'&'0'&'0'&\N__27120\&'0'&'0'&'0'&\N__30779\&'0'&'0'&'0'&\N__23109\&'0';
    buf_data_iac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(13);
    buf_data_vac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(9);
    buf_data_iac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(5);
    buf_data_vac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ <= '0'&\N__41844\&\N__39402\&\N__32904\&\N__36071\&\N__41360\&\N__36396\&\N__35925\&\N__39860\&\N__39269\&\N__40991\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ <= '0'&\N__33867\&\N__33978\&\N__34082\&\N__34194\&\N__33179\&\N__33282\&\N__33393\&\N__33504\&\N__33612\&\N__33714\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ <= '0'&'0'&\N__33079\&'0'&'0'&'0'&\N__28320\&'0'&'0'&'0'&\N__30609\&'0'&'0'&'0'&\N__27486\&'0';
    buf_data_iac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(13);
    buf_data_vac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(9);
    buf_data_iac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(5);
    buf_data_vac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ <= '0'&\N__41831\&\N__39389\&\N__32888\&\N__36068\&\N__41357\&\N__36380\&\N__35909\&\N__39851\&\N__39260\&\N__40982\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ <= '0'&\N__33851\&\N__33965\&\N__34079\&\N__34181\&\N__33170\&\N__33263\&\N__33377\&\N__33488\&\N__33599\&\N__33701\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ <= '0'&'0'&\N__24237\&'0'&'0'&'0'&\N__24264\&'0'&'0'&'0'&\N__21315\&'0'&'0'&'0'&\N__21288\&'0';
    buf_data_iac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(13);
    buf_data_vac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(9);
    buf_data_iac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(5);
    buf_data_vac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ <= '0'&\N__41850\&\N__39408\&\N__32910\&\N__36081\&\N__41370\&\N__36402\&\N__35931\&\N__39867\&\N__39276\&\N__40998\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ <= '0'&\N__33873\&\N__33984\&\N__34092\&\N__34200\&\N__33186\&\N__33288\&\N__33399\&\N__33510\&\N__33618\&\N__33720\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ <= '0'&'0'&\N__42054\&'0'&'0'&'0'&\N__28440\&'0'&'0'&'0'&\N__43392\&'0'&'0'&'0'&\N__32472\&'0';
    buf_data_iac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(13);
    buf_data_vac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(9);
    buf_data_iac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(5);
    buf_data_vac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ <= '0'&\N__41843\&\N__39401\&\N__32900\&\N__36080\&\N__41369\&\N__36392\&\N__35921\&\N__39863\&\N__39272\&\N__40994\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ <= '0'&\N__33863\&\N__33977\&\N__34091\&\N__34193\&\N__33182\&\N__33275\&\N__33389\&\N__33500\&\N__33611\&\N__33713\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ <= '0'&'0'&\N__21405\&'0'&'0'&'0'&\N__20040\&'0'&'0'&'0'&\N__20841\&'0'&'0'&'0'&\N__23142\&'0';
    buf_data_iac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(13);
    buf_data_vac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(9);
    buf_data_iac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(5);
    buf_data_vac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ <= '0'&\N__41874\&\N__39432\&\N__32934\&\N__36105\&\N__41394\&\N__36426\&\N__35955\&\N__39891\&\N__39300\&\N__41022\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ <= '0'&\N__33897\&\N__34008\&\N__34116\&\N__34224\&\N__33210\&\N__33312\&\N__33423\&\N__33534\&\N__33642\&\N__33744\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ <= '0'&'0'&\N__22857\&'0'&'0'&'0'&\N__23268\&'0'&'0'&'0'&\N__24300\&'0'&'0'&'0'&\N__23169\&'0';
    buf_data_iac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(13);
    buf_data_vac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(9);
    buf_data_iac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(5);
    buf_data_vac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ <= '0'&\N__41856\&\N__39414\&\N__32916\&\N__36087\&\N__41376\&\N__36408\&\N__35937\&\N__39873\&\N__39282\&\N__41004\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ <= '0'&\N__33879\&\N__33990\&\N__34098\&\N__34206\&\N__33192\&\N__33294\&\N__33405\&\N__33516\&\N__33624\&\N__33726\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ <= '0'&'0'&\N__24759\&'0'&'0'&'0'&\N__24528\&'0'&'0'&'0'&\N__39143\&'0'&'0'&'0'&\N__25782\&'0';
    buf_data_iac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(13);
    buf_data_vac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(9);
    buf_data_iac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(5);
    buf_data_vac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ <= '0'&\N__41868\&\N__39426\&\N__32928\&\N__36099\&\N__41388\&\N__36420\&\N__35949\&\N__39885\&\N__39294\&\N__41016\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ <= '0'&\N__33891\&\N__34002\&\N__34110\&\N__34218\&\N__33204\&\N__33306\&\N__33417\&\N__33528\&\N__33636\&\N__33738\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ <= '0'&'0'&\N__36315\&'0'&'0'&'0'&\N__32184\&'0'&'0'&'0'&\N__27237\&'0'&'0'&'0'&\N__27273\&'0';

    \pll_main.zim_pll_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => OPEN,
            REFERENCECLK => \N__19413\,
            RESETB => \N__58773\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => \clk_16MHz\,
            DYNAMICDELAY => \pll_main.zim_pll_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \clk_32MHz\,
            SCLK => \GNDG0\
        );

    \iac_raw_buf_vac_raw_buf_merged2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56042\,
            RE => \N__58486\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            WE => \N__28614\
        );

    \iac_raw_buf_vac_raw_buf_merged7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56102\,
            RE => \N__58776\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            WE => \N__28626\
        );

    \iac_raw_buf_vac_raw_buf_merged1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55962\,
            RE => \N__58762\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            WE => \N__28631\
        );

    \iac_raw_buf_vac_raw_buf_merged6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56100\,
            RE => \N__58775\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            WE => \N__28621\
        );

    \iac_raw_buf_vac_raw_buf_merged0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55948\,
            RE => \N__58763\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            WE => \N__28632\
        );

    \iac_raw_buf_vac_raw_buf_merged5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56097\,
            RE => \N__58766\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            WE => \N__28610\
        );

    \iac_raw_buf_vac_raw_buf_merged9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55997\,
            RE => \N__58758\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            WE => \N__28571\
        );

    \iac_raw_buf_vac_raw_buf_merged4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56090\,
            RE => \N__58764\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            WE => \N__28575\
        );

    \iac_raw_buf_vac_raw_buf_merged8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55972\,
            RE => \N__58774\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            WE => \N__28602\
        );

    \iac_raw_buf_vac_raw_buf_merged10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55984\,
            RE => \N__58720\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            WE => \N__28627\
        );

    \iac_raw_buf_vac_raw_buf_merged3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56071\,
            RE => \N__58728\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            WE => \N__28603\
        );

    \iac_raw_buf_vac_raw_buf_merged11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__56012\,
            RE => \N__58719\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            WE => \N__28622\
        );

    \ipInertedIOPad_VAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59914\,
            DIN => \N__59913\,
            DOUT => \N__59912\,
            PACKAGEPIN => \VAC_DRDY_wire\
        );

    \ipInertedIOPad_VAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59914\,
            PADOUT => \N__59913\,
            PADIN => \N__59912\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59905\,
            DIN => \N__59904\,
            DOUT => \N__59903\,
            PACKAGEPIN => \IAC_FLT1_wire\
        );

    \ipInertedIOPad_IAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59905\,
            PADOUT => \N__59904\,
            PADIN => \N__59903\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26502\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59896\,
            DIN => \N__59895\,
            DOUT => \N__59894\,
            PACKAGEPIN => \DDS_SCK_wire\
        );

    \ipInertedIOPad_DDS_SCK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59896\,
            PADOUT => \N__59895\,
            PADIN => \N__59894\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39036\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_166_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59887\,
            DIN => \N__59886\,
            DOUT => \N__59885\,
            PACKAGEPIN => \ICE_IOR_166_wire\
        );

    \ipInertedIOPad_ICE_IOR_166_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59887\,
            PADOUT => \N__59886\,
            PADIN => \N__59885\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_119_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59878\,
            DIN => \N__59877\,
            DOUT => \N__59876\,
            PACKAGEPIN => \ICE_IOR_119_wire\
        );

    \ipInertedIOPad_ICE_IOR_119_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59878\,
            PADOUT => \N__59877\,
            PADIN => \N__59876\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59869\,
            DIN => \N__59868\,
            DOUT => \N__59867\,
            PACKAGEPIN => \DDS_MOSI_wire\
        );

    \ipInertedIOPad_DDS_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59869\,
            PADOUT => \N__59868\,
            PADIN => \N__59867\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__38985\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59860\,
            DIN => \N__59859\,
            DOUT => \N__59858\,
            PACKAGEPIN => \VAC_MISO_wire\
        );

    \ipInertedIOPad_VAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59860\,
            PADOUT => \N__59859\,
            PADIN => \N__59858\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59851\,
            DIN => \N__59850\,
            DOUT => \N__59849\,
            PACKAGEPIN => \DDS_MOSI1_wire\
        );

    \ipInertedIOPad_DDS_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59851\,
            PADOUT => \N__59850\,
            PADIN => \N__59849\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__22773\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_146_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59842\,
            DIN => \N__59841\,
            DOUT => \N__59840\,
            PACKAGEPIN => \ICE_IOR_146_wire\
        );

    \ipInertedIOPad_ICE_IOR_146_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59842\,
            PADOUT => \N__59841\,
            PADIN => \N__59840\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59833\,
            DIN => \N__59832\,
            DOUT => \N__59831\,
            PACKAGEPIN => \VDC_CLK_wire\
        );

    \ipInertedIOPad_VDC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59833\,
            PADOUT => \N__59832\,
            PADIN => \N__59831\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__42435\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_222_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59824\,
            DIN => \N__59823\,
            DOUT => \N__59822\,
            PACKAGEPIN => \ICE_IOT_222_wire\
        );

    \ipInertedIOPad_ICE_IOT_222_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59824\,
            PADOUT => \N__59823\,
            PADIN => \N__59822\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59815\,
            DIN => \N__59814\,
            DOUT => \N__59813\,
            PACKAGEPIN => \IAC_CS_wire\
        );

    \ipInertedIOPad_IAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59815\,
            PADOUT => \N__59814\,
            PADIN => \N__59813\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21879\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_18B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59806\,
            DIN => \N__59805\,
            DOUT => \N__59804\,
            PACKAGEPIN => \ICE_IOL_18B_wire\
        );

    \ipInertedIOPad_ICE_IOL_18B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59806\,
            PADOUT => \N__59805\,
            PADIN => \N__59804\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59797\,
            DIN => \N__59796\,
            DOUT => \N__59795\,
            PACKAGEPIN => \ICE_IOL_13A_wire\
        );

    \ipInertedIOPad_ICE_IOL_13A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59797\,
            PADOUT => \N__59796\,
            PADIN => \N__59795\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_81_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59788\,
            DIN => \N__59787\,
            DOUT => \N__59786\,
            PACKAGEPIN => \ICE_IOB_81_wire\
        );

    \ipInertedIOPad_ICE_IOB_81_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59788\,
            PADOUT => \N__59787\,
            PADIN => \N__59786\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59779\,
            DIN => \N__59778\,
            DOUT => \N__59777\,
            PACKAGEPIN => \VAC_OSR1_wire\
        );

    \ipInertedIOPad_VAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59779\,
            PADOUT => \N__59778\,
            PADIN => \N__59777\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27390\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59770\,
            DIN => \N__59769\,
            DOUT => \N__59768\,
            PACKAGEPIN => \IAC_MOSI_wire\
        );

    \ipInertedIOPad_IAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59770\,
            PADOUT => \N__59769\,
            PADIN => \N__59768\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59761\,
            DIN => \N__59760\,
            DOUT => \N__59759\,
            PACKAGEPIN => \DDS_CS1_wire\
        );

    \ipInertedIOPad_DDS_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59761\,
            PADOUT => \N__59760\,
            PADIN => \N__59759\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21858\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59752\,
            DIN => \N__59751\,
            DOUT => \N__59750\,
            PACKAGEPIN => \ICE_IOL_4B_wire\
        );

    \ipInertedIOPad_ICE_IOL_4B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59752\,
            PADOUT => \N__59751\,
            PADIN => \N__59750\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_94_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59743\,
            DIN => \N__59742\,
            DOUT => \N__59741\,
            PACKAGEPIN => \ICE_IOB_94_wire\
        );

    \ipInertedIOPad_ICE_IOB_94_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59743\,
            PADOUT => \N__59742\,
            PADIN => \N__59741\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59734\,
            DIN => \N__59733\,
            DOUT => \N__59732\,
            PACKAGEPIN => \VAC_CS_wire\
        );

    \ipInertedIOPad_VAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59734\,
            PADOUT => \N__59733\,
            PADIN => \N__59732\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21660\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59725\,
            DIN => \N__59724\,
            DOUT => \N__59723\,
            PACKAGEPIN => \VAC_CLK_wire\
        );

    \ipInertedIOPad_VAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59725\,
            PADOUT => \N__59724\,
            PADIN => \N__59723\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31121\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_CE0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59716\,
            DIN => \N__59715\,
            DOUT => \N__59714\,
            PACKAGEPIN => \ICE_SPI_CE0_wire\
        );

    \ipInertedIOPad_ICE_SPI_CE0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59716\,
            PADOUT => \N__59715\,
            PADIN => \N__59714\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_CE0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_167_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59707\,
            DIN => \N__59706\,
            DOUT => \N__59705\,
            PACKAGEPIN => \ICE_IOR_167_wire\
        );

    \ipInertedIOPad_ICE_IOR_167_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59707\,
            PADOUT => \N__59706\,
            PADIN => \N__59705\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_118_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59698\,
            DIN => \N__59697\,
            DOUT => \N__59696\,
            PACKAGEPIN => \ICE_IOR_118_wire\
        );

    \ipInertedIOPad_ICE_IOR_118_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59698\,
            PADOUT => \N__59697\,
            PADIN => \N__59696\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDO_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59689\,
            DIN => \N__59688\,
            DOUT => \N__59687\,
            PACKAGEPIN => \RTD_SDO_wire\
        );

    \ipInertedIOPad_RTD_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59689\,
            PADOUT => \N__59688\,
            PADIN => \N__59687\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59680\,
            DIN => \N__59679\,
            DOUT => \N__59678\,
            PACKAGEPIN => \IAC_OSR0_wire\
        );

    \ipInertedIOPad_IAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59680\,
            PADOUT => \N__59679\,
            PADIN => \N__59678\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__39474\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59671\,
            DIN => \N__59670\,
            DOUT => \N__59669\,
            PACKAGEPIN => \VDC_SCLK_wire\
        );

    \ipInertedIOPad_VDC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59671\,
            PADOUT => \N__59670\,
            PADIN => \N__59669\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__42462\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59662\,
            DIN => \N__59661\,
            DOUT => \N__59660\,
            PACKAGEPIN => \VAC_FLT1_wire\
        );

    \ipInertedIOPad_VAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59662\,
            PADOUT => \N__59661\,
            PADIN => \N__59660\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29007\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MOSI_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59653\,
            DIN => \N__59652\,
            DOUT => \N__59651\,
            PACKAGEPIN => \ICE_SPI_MOSI_wire\
        );

    \ipInertedIOPad_ICE_SPI_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59653\,
            PADOUT => \N__59652\,
            PADIN => \N__59651\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_MOSI\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_165_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59644\,
            DIN => \N__59643\,
            DOUT => \N__59642\,
            PACKAGEPIN => \ICE_IOR_165_wire\
        );

    \ipInertedIOPad_ICE_IOR_165_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59644\,
            PADOUT => \N__59643\,
            PADIN => \N__59642\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_147_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59635\,
            DIN => \N__59634\,
            DOUT => \N__59633\,
            PACKAGEPIN => \ICE_IOR_147_wire\
        );

    \ipInertedIOPad_ICE_IOR_147_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59635\,
            PADOUT => \N__59634\,
            PADIN => \N__59633\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_14A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59626\,
            DIN => \N__59625\,
            DOUT => \N__59624\,
            PACKAGEPIN => \ICE_IOL_14A_wire\
        );

    \ipInertedIOPad_ICE_IOL_14A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59626\,
            PADOUT => \N__59625\,
            PADIN => \N__59624\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59617\,
            DIN => \N__59616\,
            DOUT => \N__59615\,
            PACKAGEPIN => \ICE_IOL_13B_wire\
        );

    \ipInertedIOPad_ICE_IOL_13B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59617\,
            PADOUT => \N__59616\,
            PADIN => \N__59615\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_91_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59608\,
            DIN => \N__59607\,
            DOUT => \N__59606\,
            PACKAGEPIN => \ICE_IOB_91_wire\
        );

    \ipInertedIOPad_ICE_IOB_91_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59608\,
            PADOUT => \N__59607\,
            PADIN => \N__59606\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59599\,
            DIN => \N__59598\,
            DOUT => \N__59597\,
            PACKAGEPIN => \ICE_GPMO_0_wire\
        );

    \ipInertedIOPad_ICE_GPMO_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59599\,
            PADOUT => \N__59598\,
            PADIN => \N__59597\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_RNG_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59590\,
            DIN => \N__59589\,
            DOUT => \N__59588\,
            PACKAGEPIN => \DDS_RNG_0_wire\
        );

    \ipInertedIOPad_DDS_RNG_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59590\,
            PADOUT => \N__59589\,
            PADIN => \N__59588\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__42957\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_RNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59581\,
            DIN => \N__59580\,
            DOUT => \N__59579\,
            PACKAGEPIN => \VDC_RNG0_wire\
        );

    \ipInertedIOPad_VDC_RNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59581\,
            PADOUT => \N__59580\,
            PADIN => \N__59579\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__41517\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_SCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59572\,
            DIN => \N__59571\,
            DOUT => \N__59570\,
            PACKAGEPIN => \ICE_SPI_SCLK_wire\
        );

    \ipInertedIOPad_ICE_SPI_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59572\,
            PADOUT => \N__59571\,
            PADIN => \N__59570\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_SCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_152_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59563\,
            DIN => \N__59562\,
            DOUT => \N__59561\,
            PACKAGEPIN => \ICE_IOR_152_wire\
        );

    \ipInertedIOPad_ICE_IOR_152_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59563\,
            PADOUT => \N__59562\,
            PADIN => \N__59561\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59554\,
            DIN => \N__59553\,
            DOUT => \N__59552\,
            PACKAGEPIN => \ICE_IOL_12A_wire\
        );

    \ipInertedIOPad_ICE_IOL_12A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59554\,
            PADOUT => \N__59553\,
            PADIN => \N__59552\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_DRDY_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59545\,
            DIN => \N__59544\,
            DOUT => \N__59543\,
            PACKAGEPIN => \RTD_DRDY_wire\
        );

    \ipInertedIOPad_RTD_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59545\,
            PADOUT => \N__59544\,
            PADIN => \N__59543\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59536\,
            DIN => \N__59535\,
            DOUT => \N__59534\,
            PACKAGEPIN => \ICE_SPI_MISO_wire\
        );

    \ipInertedIOPad_ICE_SPI_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59536\,
            PADOUT => \N__59535\,
            PADIN => \N__59534\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44283\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_177_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59527\,
            DIN => \N__59526\,
            DOUT => \N__59525\,
            PACKAGEPIN => \ICE_IOT_177_wire\
        );

    \ipInertedIOPad_ICE_IOT_177_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59527\,
            PADOUT => \N__59526\,
            PADIN => \N__59525\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_141_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59518\,
            DIN => \N__59517\,
            DOUT => \N__59516\,
            PACKAGEPIN => \ICE_IOR_141_wire\
        );

    \ipInertedIOPad_ICE_IOR_141_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59518\,
            PADOUT => \N__59517\,
            PADIN => \N__59516\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_80_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59509\,
            DIN => \N__59508\,
            DOUT => \N__59507\,
            PACKAGEPIN => \ICE_IOB_80_wire\
        );

    \ipInertedIOPad_ICE_IOB_80_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59509\,
            PADOUT => \N__59508\,
            PADIN => \N__59507\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_102_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59500\,
            DIN => \N__59499\,
            DOUT => \N__59498\,
            PACKAGEPIN => \ICE_IOB_102_wire\
        );

    \ipInertedIOPad_ICE_IOB_102_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59500\,
            PADOUT => \N__59499\,
            PADIN => \N__59498\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59491\,
            DIN => \N__59490\,
            DOUT => \N__59489\,
            PACKAGEPIN => \ICE_GPMO_2_wire\
        );

    \ipInertedIOPad_ICE_GPMO_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59491\,
            PADOUT => \N__59490\,
            PADIN => \N__59489\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMI_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59482\,
            DIN => \N__59481\,
            DOUT => \N__59480\,
            PACKAGEPIN => \ICE_GPMI_0_wire\
        );

    \ipInertedIOPad_ICE_GPMI_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59482\,
            PADOUT => \N__59481\,
            PADIN => \N__59480\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__56118\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59473\,
            DIN => \N__59472\,
            DOUT => \N__59471\,
            PACKAGEPIN => \IAC_MISO_wire\
        );

    \ipInertedIOPad_IAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59473\,
            PADOUT => \N__59472\,
            PADIN => \N__59471\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59464\,
            DIN => \N__59463\,
            DOUT => \N__59462\,
            PACKAGEPIN => \VAC_OSR0_wire\
        );

    \ipInertedIOPad_VAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59464\,
            PADOUT => \N__59463\,
            PADIN => \N__59462\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32106\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59455\,
            DIN => \N__59454\,
            DOUT => \N__59453\,
            PACKAGEPIN => \VAC_MOSI_wire\
        );

    \ipInertedIOPad_VAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59455\,
            PADOUT => \N__59454\,
            PADIN => \N__59453\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TEST_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59446\,
            DIN => \N__59445\,
            DOUT => \N__59444\,
            PACKAGEPIN => \TEST_LED_wire\
        );

    \ipInertedIOPad_TEST_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59446\,
            PADOUT => \N__59445\,
            PADIN => \N__59444\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__34677\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_148_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59437\,
            DIN => \N__59436\,
            DOUT => \N__59435\,
            PACKAGEPIN => \ICE_IOR_148_wire\
        );

    \ipInertedIOPad_ICE_IOR_148_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59437\,
            PADOUT => \N__59436\,
            PADIN => \N__59435\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_STAT_COMM_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59428\,
            DIN => \N__59427\,
            DOUT => \N__59426\,
            PACKAGEPIN => \STAT_COMM_wire\
        );

    \ipInertedIOPad_STAT_COMM_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59428\,
            PADOUT => \N__59427\,
            PADIN => \N__59426\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19398\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SYSCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59419\,
            DIN => \N__59418\,
            DOUT => \N__59417\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ipInertedIOPad_ICE_SYSCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59419\,
            PADOUT => \N__59418\,
            PADIN => \N__59417\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SYSCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_161_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59410\,
            DIN => \N__59409\,
            DOUT => \N__59408\,
            PACKAGEPIN => \ICE_IOR_161_wire\
        );

    \ipInertedIOPad_ICE_IOR_161_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59410\,
            PADOUT => \N__59409\,
            PADIN => \N__59408\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_95_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59401\,
            DIN => \N__59400\,
            DOUT => \N__59399\,
            PACKAGEPIN => \ICE_IOB_95_wire\
        );

    \ipInertedIOPad_ICE_IOB_95_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59401\,
            PADOUT => \N__59400\,
            PADIN => \N__59399\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_82_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59392\,
            DIN => \N__59391\,
            DOUT => \N__59390\,
            PACKAGEPIN => \ICE_IOB_82_wire\
        );

    \ipInertedIOPad_ICE_IOB_82_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59392\,
            PADOUT => \N__59391\,
            PADIN => \N__59390\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_104_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59383\,
            DIN => \N__59382\,
            DOUT => \N__59381\,
            PACKAGEPIN => \ICE_IOB_104_wire\
        );

    \ipInertedIOPad_ICE_IOB_104_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59383\,
            PADOUT => \N__59382\,
            PADIN => \N__59381\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59374\,
            DIN => \N__59373\,
            DOUT => \N__59372\,
            PACKAGEPIN => \IAC_CLK_wire\
        );

    \ipInertedIOPad_IAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59374\,
            PADOUT => \N__59373\,
            PADIN => \N__59372\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__31125\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59365\,
            DIN => \N__59364\,
            DOUT => \N__59363\,
            PACKAGEPIN => \DDS_CS_wire\
        );

    \ipInertedIOPad_DDS_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59365\,
            PADOUT => \N__59364\,
            PADIN => \N__59363\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__41949\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59356\,
            DIN => \N__59355\,
            DOUT => \N__59354\,
            PACKAGEPIN => \SELIRNG0_wire\
        );

    \ipInertedIOPad_SELIRNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59356\,
            PADOUT => \N__59355\,
            PADIN => \N__59354\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__45738\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59347\,
            DIN => \N__59346\,
            DOUT => \N__59345\,
            PACKAGEPIN => \RTD_SDI_wire\
        );

    \ipInertedIOPad_RTD_SDI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59347\,
            PADOUT => \N__59346\,
            PADIN => \N__59345\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19560\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_221_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59338\,
            DIN => \N__59337\,
            DOUT => \N__59336\,
            PACKAGEPIN => \ICE_IOT_221_wire\
        );

    \ipInertedIOPad_ICE_IOT_221_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59338\,
            PADOUT => \N__59337\,
            PADIN => \N__59336\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_197_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59329\,
            DIN => \N__59328\,
            DOUT => \N__59327\,
            PACKAGEPIN => \ICE_IOT_197_wire\
        );

    \ipInertedIOPad_ICE_IOT_197_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59329\,
            PADOUT => \N__59328\,
            PADIN => \N__59327\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59320\,
            DIN => \N__59319\,
            DOUT => \N__59318\,
            PACKAGEPIN => \DDS_MCLK_wire\
        );

    \ipInertedIOPad_DDS_MCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59320\,
            PADOUT => \N__59319\,
            PADIN => \N__59318\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__50691\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59311\,
            DIN => \N__59310\,
            DOUT => \N__59309\,
            PACKAGEPIN => \RTD_SCLK_wire\
        );

    \ipInertedIOPad_RTD_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59311\,
            PADOUT => \N__59310\,
            PADIN => \N__59309\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19539\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59302\,
            DIN => \N__59301\,
            DOUT => \N__59300\,
            PACKAGEPIN => \RTD_CS_wire\
        );

    \ipInertedIOPad_RTD_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59302\,
            PADOUT => \N__59301\,
            PADIN => \N__59300\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20322\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_137_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59293\,
            DIN => \N__59292\,
            DOUT => \N__59291\,
            PACKAGEPIN => \ICE_IOR_137_wire\
        );

    \ipInertedIOPad_ICE_IOR_137_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59293\,
            PADOUT => \N__59292\,
            PADIN => \N__59291\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59284\,
            DIN => \N__59283\,
            DOUT => \N__59282\,
            PACKAGEPIN => \IAC_OSR1_wire\
        );

    \ipInertedIOPad_IAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59284\,
            PADOUT => \N__59283\,
            PADIN => \N__59282\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26100\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59275\,
            DIN => \N__59274\,
            DOUT => \N__59273\,
            PACKAGEPIN => \VAC_FLT0_wire\
        );

    \ipInertedIOPad_VAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59275\,
            PADOUT => \N__59274\,
            PADIN => \N__59273\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30822\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_144_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59266\,
            DIN => \N__59265\,
            DOUT => \N__59264\,
            PACKAGEPIN => \ICE_IOR_144_wire\
        );

    \ipInertedIOPad_ICE_IOR_144_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59266\,
            PADOUT => \N__59265\,
            PADIN => \N__59264\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_128_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59257\,
            DIN => \N__59256\,
            DOUT => \N__59255\,
            PACKAGEPIN => \ICE_IOR_128_wire\
        );

    \ipInertedIOPad_ICE_IOR_128_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59257\,
            PADOUT => \N__59256\,
            PADIN => \N__59255\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59248\,
            DIN => \N__59247\,
            DOUT => \N__59246\,
            PACKAGEPIN => \ICE_GPMO_1_wire\
        );

    \ipInertedIOPad_ICE_GPMO_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59248\,
            PADOUT => \N__59247\,
            PADIN => \N__59246\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59239\,
            DIN => \N__59238\,
            DOUT => \N__59237\,
            PACKAGEPIN => \IAC_SCLK_wire\
        );

    \ipInertedIOPad_IAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59239\,
            PADOUT => \N__59238\,
            PADIN => \N__59237\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24786\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_EIS_SYNCCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59230\,
            DIN => \N__59229\,
            DOUT => \N__59228\,
            PACKAGEPIN => \EIS_SYNCCLK_wire\
        );

    \ipInertedIOPad_EIS_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59230\,
            PADOUT => \N__59229\,
            PADIN => \N__59228\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \EIS_SYNCCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_139_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59221\,
            DIN => \N__59220\,
            DOUT => \N__59219\,
            PACKAGEPIN => \ICE_IOR_139_wire\
        );

    \ipInertedIOPad_ICE_IOR_139_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59221\,
            PADOUT => \N__59220\,
            PADIN => \N__59219\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59212\,
            DIN => \N__59211\,
            DOUT => \N__59210\,
            PACKAGEPIN => \ICE_IOL_4A_wire\
        );

    \ipInertedIOPad_ICE_IOL_4A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59212\,
            PADOUT => \N__59211\,
            PADIN => \N__59210\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59203\,
            DIN => \N__59202\,
            DOUT => \N__59201\,
            PACKAGEPIN => \VAC_SCLK_wire\
        );

    \ipInertedIOPad_VAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59203\,
            PADOUT => \N__59202\,
            PADIN => \N__59201\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21468\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_THERMOSTAT_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59194\,
            DIN => \N__59193\,
            DOUT => \N__59192\,
            PACKAGEPIN => \THERMOSTAT_wire\
        );

    \ipInertedIOPad_THERMOSTAT_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59194\,
            PADOUT => \N__59193\,
            PADIN => \N__59192\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \THERMOSTAT\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_164_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59185\,
            DIN => \N__59184\,
            DOUT => \N__59183\,
            PACKAGEPIN => \ICE_IOR_164_wire\
        );

    \ipInertedIOPad_ICE_IOR_164_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59185\,
            PADOUT => \N__59184\,
            PADIN => \N__59183\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_103_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59176\,
            DIN => \N__59175\,
            DOUT => \N__59174\,
            PACKAGEPIN => \ICE_IOB_103_wire\
        );

    \ipInertedIOPad_ICE_IOB_103_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59176\,
            PADOUT => \N__59175\,
            PADIN => \N__59174\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AMPV_POW_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59167\,
            DIN => \N__59166\,
            DOUT => \N__59165\,
            PACKAGEPIN => \AMPV_POW_wire\
        );

    \ipInertedIOPad_AMPV_POW_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59167\,
            PADOUT => \N__59166\,
            PADIN => \N__59165\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36015\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SDO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59158\,
            DIN => \N__59157\,
            DOUT => \N__59156\,
            PACKAGEPIN => \VDC_SDO_wire\
        );

    \ipInertedIOPad_VDC_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59158\,
            PADOUT => \N__59157\,
            PADIN => \N__59156\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VDC_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_174_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59149\,
            DIN => \N__59148\,
            DOUT => \N__59147\,
            PACKAGEPIN => \ICE_IOT_174_wire\
        );

    \ipInertedIOPad_ICE_IOT_174_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59149\,
            PADOUT => \N__59148\,
            PADIN => \N__59147\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_140_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59140\,
            DIN => \N__59139\,
            DOUT => \N__59138\,
            PACKAGEPIN => \ICE_IOR_140_wire\
        );

    \ipInertedIOPad_ICE_IOR_140_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59140\,
            PADOUT => \N__59139\,
            PADIN => \N__59138\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_96_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59131\,
            DIN => \N__59130\,
            DOUT => \N__59129\,
            PACKAGEPIN => \ICE_IOB_96_wire\
        );

    \ipInertedIOPad_ICE_IOB_96_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59131\,
            PADOUT => \N__59130\,
            PADIN => \N__59129\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CONT_SD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59122\,
            DIN => \N__59121\,
            DOUT => \N__59120\,
            PACKAGEPIN => \CONT_SD_wire\
        );

    \ipInertedIOPad_CONT_SD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59122\,
            PADOUT => \N__59121\,
            PADIN => \N__59120\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44775\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AC_ADC_SYNC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59113\,
            DIN => \N__59112\,
            DOUT => \N__59111\,
            PACKAGEPIN => \AC_ADC_SYNC_wire\
        );

    \ipInertedIOPad_AC_ADC_SYNC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59113\,
            PADOUT => \N__59112\,
            PADIN => \N__59111\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21903\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59104\,
            DIN => \N__59103\,
            DOUT => \N__59102\,
            PACKAGEPIN => \SELIRNG1_wire\
        );

    \ipInertedIOPad_SELIRNG1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59104\,
            PADOUT => \N__59103\,
            PADIN => \N__59102\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36225\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59095\,
            DIN => \N__59094\,
            DOUT => \N__59093\,
            PACKAGEPIN => \ICE_IOL_12B_wire\
        );

    \ipInertedIOPad_ICE_IOL_12B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59095\,
            PADOUT => \N__59094\,
            PADIN => \N__59093\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_160_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59086\,
            DIN => \N__59085\,
            DOUT => \N__59084\,
            PACKAGEPIN => \ICE_IOR_160_wire\
        );

    \ipInertedIOPad_ICE_IOR_160_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59086\,
            PADOUT => \N__59085\,
            PADIN => \N__59084\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_136_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59077\,
            DIN => \N__59076\,
            DOUT => \N__59075\,
            PACKAGEPIN => \ICE_IOR_136_wire\
        );

    \ipInertedIOPad_ICE_IOR_136_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59077\,
            PADOUT => \N__59076\,
            PADIN => \N__59075\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59068\,
            DIN => \N__59067\,
            DOUT => \N__59066\,
            PACKAGEPIN => \DDS_MCLK1_wire\
        );

    \ipInertedIOPad_DDS_MCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59068\,
            PADOUT => \N__59067\,
            PADIN => \N__59066\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23751\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_198_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59059\,
            DIN => \N__59058\,
            DOUT => \N__59057\,
            PACKAGEPIN => \ICE_IOT_198_wire\
        );

    \ipInertedIOPad_ICE_IOT_198_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59059\,
            PADOUT => \N__59058\,
            PADIN => \N__59057\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_173_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59050\,
            DIN => \N__59049\,
            DOUT => \N__59048\,
            PACKAGEPIN => \ICE_IOT_173_wire\
        );

    \ipInertedIOPad_ICE_IOT_173_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59050\,
            PADOUT => \N__59049\,
            PADIN => \N__59048\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59041\,
            DIN => \N__59040\,
            DOUT => \N__59039\,
            PACKAGEPIN => \IAC_DRDY_wire\
        );

    \ipInertedIOPad_IAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59041\,
            PADOUT => \N__59040\,
            PADIN => \N__59039\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_178_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59032\,
            DIN => \N__59031\,
            DOUT => \N__59030\,
            PACKAGEPIN => \ICE_IOT_178_wire\
        );

    \ipInertedIOPad_ICE_IOT_178_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59032\,
            PADOUT => \N__59031\,
            PADIN => \N__59030\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_138_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59023\,
            DIN => \N__59022\,
            DOUT => \N__59021\,
            PACKAGEPIN => \ICE_IOR_138_wire\
        );

    \ipInertedIOPad_ICE_IOR_138_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59023\,
            PADOUT => \N__59022\,
            PADIN => \N__59021\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_120_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__59014\,
            DIN => \N__59013\,
            DOUT => \N__59012\,
            PACKAGEPIN => \ICE_IOR_120_wire\
        );

    \ipInertedIOPad_ICE_IOR_120_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59014\,
            PADOUT => \N__59013\,
            PADIN => \N__59012\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__59005\,
            DIN => \N__59004\,
            DOUT => \N__59003\,
            PACKAGEPIN => \IAC_FLT0_wire\
        );

    \ipInertedIOPad_IAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__59005\,
            PADOUT => \N__59004\,
            PADIN => \N__59003\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30546\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58996\,
            DIN => \N__58995\,
            DOUT => \N__58994\,
            PACKAGEPIN => \DDS_SCK1_wire\
        );

    \ipInertedIOPad_DDS_SCK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58996\,
            PADOUT => \N__58995\,
            PADIN => \N__58994\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27189\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__14786\ : SRMux
    port map (
            O => \N__58977\,
            I => \N__58974\
        );

    \I__14785\ : LocalMux
    port map (
            O => \N__58974\,
            I => \N__58969\
        );

    \I__14784\ : SRMux
    port map (
            O => \N__58973\,
            I => \N__58965\
        );

    \I__14783\ : SRMux
    port map (
            O => \N__58972\,
            I => \N__58962\
        );

    \I__14782\ : Span4Mux_h
    port map (
            O => \N__58969\,
            I => \N__58959\
        );

    \I__14781\ : SRMux
    port map (
            O => \N__58968\,
            I => \N__58956\
        );

    \I__14780\ : LocalMux
    port map (
            O => \N__58965\,
            I => \N__58953\
        );

    \I__14779\ : LocalMux
    port map (
            O => \N__58962\,
            I => \N__58950\
        );

    \I__14778\ : Span4Mux_h
    port map (
            O => \N__58959\,
            I => \N__58945\
        );

    \I__14777\ : LocalMux
    port map (
            O => \N__58956\,
            I => \N__58945\
        );

    \I__14776\ : Span4Mux_h
    port map (
            O => \N__58953\,
            I => \N__58942\
        );

    \I__14775\ : Span4Mux_v
    port map (
            O => \N__58950\,
            I => \N__58939\
        );

    \I__14774\ : Span4Mux_v
    port map (
            O => \N__58945\,
            I => \N__58934\
        );

    \I__14773\ : Span4Mux_h
    port map (
            O => \N__58942\,
            I => \N__58934\
        );

    \I__14772\ : Span4Mux_h
    port map (
            O => \N__58939\,
            I => \N__58931\
        );

    \I__14771\ : Odrv4
    port map (
            O => \N__58934\,
            I => \ADC_VDC.genclk.n14894\
        );

    \I__14770\ : Odrv4
    port map (
            O => \N__58931\,
            I => \ADC_VDC.genclk.n14894\
        );

    \I__14769\ : SRMux
    port map (
            O => \N__58926\,
            I => \N__58923\
        );

    \I__14768\ : LocalMux
    port map (
            O => \N__58923\,
            I => \N__58920\
        );

    \I__14767\ : Span4Mux_v
    port map (
            O => \N__58920\,
            I => \N__58917\
        );

    \I__14766\ : Odrv4
    port map (
            O => \N__58917\,
            I => \comm_spi.data_tx_7__N_835\
        );

    \I__14765\ : InMux
    port map (
            O => \N__58914\,
            I => \N__58911\
        );

    \I__14764\ : LocalMux
    port map (
            O => \N__58911\,
            I => \N__58907\
        );

    \I__14763\ : InMux
    port map (
            O => \N__58910\,
            I => \N__58904\
        );

    \I__14762\ : Span4Mux_v
    port map (
            O => \N__58907\,
            I => \N__58899\
        );

    \I__14761\ : LocalMux
    port map (
            O => \N__58904\,
            I => \N__58899\
        );

    \I__14760\ : Odrv4
    port map (
            O => \N__58899\,
            I => \comm_spi.n14827\
        );

    \I__14759\ : InMux
    port map (
            O => \N__58896\,
            I => \N__58893\
        );

    \I__14758\ : LocalMux
    port map (
            O => \N__58893\,
            I => \N__58888\
        );

    \I__14757\ : InMux
    port map (
            O => \N__58892\,
            I => \N__58885\
        );

    \I__14756\ : InMux
    port map (
            O => \N__58891\,
            I => \N__58882\
        );

    \I__14755\ : Odrv4
    port map (
            O => \N__58888\,
            I => \comm_spi.n23110\
        );

    \I__14754\ : LocalMux
    port map (
            O => \N__58885\,
            I => \comm_spi.n23110\
        );

    \I__14753\ : LocalMux
    port map (
            O => \N__58882\,
            I => \comm_spi.n23110\
        );

    \I__14752\ : InMux
    port map (
            O => \N__58875\,
            I => \N__58871\
        );

    \I__14751\ : InMux
    port map (
            O => \N__58874\,
            I => \N__58868\
        );

    \I__14750\ : LocalMux
    port map (
            O => \N__58871\,
            I => \N__58863\
        );

    \I__14749\ : LocalMux
    port map (
            O => \N__58868\,
            I => \N__58863\
        );

    \I__14748\ : Odrv12
    port map (
            O => \N__58863\,
            I => \comm_spi.n14801\
        );

    \I__14747\ : InMux
    port map (
            O => \N__58860\,
            I => \N__58857\
        );

    \I__14746\ : LocalMux
    port map (
            O => \N__58857\,
            I => \N__58853\
        );

    \I__14745\ : InMux
    port map (
            O => \N__58856\,
            I => \N__58850\
        );

    \I__14744\ : Span4Mux_v
    port map (
            O => \N__58853\,
            I => \N__58847\
        );

    \I__14743\ : LocalMux
    port map (
            O => \N__58850\,
            I => \N__58844\
        );

    \I__14742\ : Odrv4
    port map (
            O => \N__58847\,
            I => \comm_spi.n14826\
        );

    \I__14741\ : Odrv12
    port map (
            O => \N__58844\,
            I => \comm_spi.n14826\
        );

    \I__14740\ : SRMux
    port map (
            O => \N__58839\,
            I => \N__58836\
        );

    \I__14739\ : LocalMux
    port map (
            O => \N__58836\,
            I => \N__58833\
        );

    \I__14738\ : Odrv4
    port map (
            O => \N__58833\,
            I => \comm_spi.data_tx_7__N_812\
        );

    \I__14737\ : SRMux
    port map (
            O => \N__58830\,
            I => \N__58827\
        );

    \I__14736\ : LocalMux
    port map (
            O => \N__58827\,
            I => \N__58824\
        );

    \I__14735\ : Span4Mux_v
    port map (
            O => \N__58824\,
            I => \N__58821\
        );

    \I__14734\ : Odrv4
    port map (
            O => \N__58821\,
            I => \comm_spi.data_tx_7__N_832\
        );

    \I__14733\ : InMux
    port map (
            O => \N__58818\,
            I => \N__58809\
        );

    \I__14732\ : InMux
    port map (
            O => \N__58817\,
            I => \N__58809\
        );

    \I__14731\ : InMux
    port map (
            O => \N__58816\,
            I => \N__58809\
        );

    \I__14730\ : LocalMux
    port map (
            O => \N__58809\,
            I => \N__58806\
        );

    \I__14729\ : Span4Mux_v
    port map (
            O => \N__58806\,
            I => \N__58803\
        );

    \I__14728\ : Odrv4
    port map (
            O => \N__58803\,
            I => comm_tx_buf_1
        );

    \I__14727\ : InMux
    port map (
            O => \N__58800\,
            I => \N__58797\
        );

    \I__14726\ : LocalMux
    port map (
            O => \N__58797\,
            I => \N__58793\
        );

    \I__14725\ : InMux
    port map (
            O => \N__58796\,
            I => \N__58790\
        );

    \I__14724\ : Span4Mux_v
    port map (
            O => \N__58793\,
            I => \N__58784\
        );

    \I__14723\ : LocalMux
    port map (
            O => \N__58790\,
            I => \N__58784\
        );

    \I__14722\ : InMux
    port map (
            O => \N__58789\,
            I => \N__58781\
        );

    \I__14721\ : Odrv4
    port map (
            O => \N__58784\,
            I => \comm_spi.n23107\
        );

    \I__14720\ : LocalMux
    port map (
            O => \N__58781\,
            I => \comm_spi.n23107\
        );

    \I__14719\ : SRMux
    port map (
            O => \N__58776\,
            I => \N__58770\
        );

    \I__14718\ : SRMux
    port map (
            O => \N__58775\,
            I => \N__58767\
        );

    \I__14717\ : SRMux
    port map (
            O => \N__58774\,
            I => \N__58759\
        );

    \I__14716\ : IoInMux
    port map (
            O => \N__58773\,
            I => \N__58755\
        );

    \I__14715\ : LocalMux
    port map (
            O => \N__58770\,
            I => \N__58738\
        );

    \I__14714\ : LocalMux
    port map (
            O => \N__58767\,
            I => \N__58738\
        );

    \I__14713\ : SRMux
    port map (
            O => \N__58766\,
            I => \N__58735\
        );

    \I__14712\ : InMux
    port map (
            O => \N__58765\,
            I => \N__58732\
        );

    \I__14711\ : SRMux
    port map (
            O => \N__58764\,
            I => \N__58729\
        );

    \I__14710\ : SRMux
    port map (
            O => \N__58763\,
            I => \N__58725\
        );

    \I__14709\ : SRMux
    port map (
            O => \N__58762\,
            I => \N__58722\
        );

    \I__14708\ : LocalMux
    port map (
            O => \N__58759\,
            I => \N__58712\
        );

    \I__14707\ : SRMux
    port map (
            O => \N__58758\,
            I => \N__58709\
        );

    \I__14706\ : LocalMux
    port map (
            O => \N__58755\,
            I => \N__58699\
        );

    \I__14705\ : CascadeMux
    port map (
            O => \N__58754\,
            I => \N__58696\
        );

    \I__14704\ : CascadeMux
    port map (
            O => \N__58753\,
            I => \N__58692\
        );

    \I__14703\ : CascadeMux
    port map (
            O => \N__58752\,
            I => \N__58688\
        );

    \I__14702\ : CascadeMux
    port map (
            O => \N__58751\,
            I => \N__58684\
        );

    \I__14701\ : CascadeMux
    port map (
            O => \N__58750\,
            I => \N__58680\
        );

    \I__14700\ : CascadeMux
    port map (
            O => \N__58749\,
            I => \N__58676\
        );

    \I__14699\ : CascadeMux
    port map (
            O => \N__58748\,
            I => \N__58672\
        );

    \I__14698\ : CascadeMux
    port map (
            O => \N__58747\,
            I => \N__58668\
        );

    \I__14697\ : CascadeMux
    port map (
            O => \N__58746\,
            I => \N__58665\
        );

    \I__14696\ : CascadeMux
    port map (
            O => \N__58745\,
            I => \N__58661\
        );

    \I__14695\ : CascadeMux
    port map (
            O => \N__58744\,
            I => \N__58657\
        );

    \I__14694\ : CascadeMux
    port map (
            O => \N__58743\,
            I => \N__58653\
        );

    \I__14693\ : Span4Mux_v
    port map (
            O => \N__58738\,
            I => \N__58644\
        );

    \I__14692\ : LocalMux
    port map (
            O => \N__58735\,
            I => \N__58644\
        );

    \I__14691\ : LocalMux
    port map (
            O => \N__58732\,
            I => \N__58644\
        );

    \I__14690\ : LocalMux
    port map (
            O => \N__58729\,
            I => \N__58644\
        );

    \I__14689\ : SRMux
    port map (
            O => \N__58728\,
            I => \N__58641\
        );

    \I__14688\ : LocalMux
    port map (
            O => \N__58725\,
            I => \N__58636\
        );

    \I__14687\ : LocalMux
    port map (
            O => \N__58722\,
            I => \N__58636\
        );

    \I__14686\ : InMux
    port map (
            O => \N__58721\,
            I => \N__58633\
        );

    \I__14685\ : SRMux
    port map (
            O => \N__58720\,
            I => \N__58630\
        );

    \I__14684\ : SRMux
    port map (
            O => \N__58719\,
            I => \N__58627\
        );

    \I__14683\ : CascadeMux
    port map (
            O => \N__58718\,
            I => \N__58623\
        );

    \I__14682\ : CascadeMux
    port map (
            O => \N__58717\,
            I => \N__58619\
        );

    \I__14681\ : CascadeMux
    port map (
            O => \N__58716\,
            I => \N__58615\
        );

    \I__14680\ : CascadeMux
    port map (
            O => \N__58715\,
            I => \N__58611\
        );

    \I__14679\ : Span4Mux_v
    port map (
            O => \N__58712\,
            I => \N__58608\
        );

    \I__14678\ : LocalMux
    port map (
            O => \N__58709\,
            I => \N__58605\
        );

    \I__14677\ : InMux
    port map (
            O => \N__58708\,
            I => \N__58598\
        );

    \I__14676\ : InMux
    port map (
            O => \N__58707\,
            I => \N__58598\
        );

    \I__14675\ : InMux
    port map (
            O => \N__58706\,
            I => \N__58598\
        );

    \I__14674\ : InMux
    port map (
            O => \N__58705\,
            I => \N__58589\
        );

    \I__14673\ : InMux
    port map (
            O => \N__58704\,
            I => \N__58589\
        );

    \I__14672\ : InMux
    port map (
            O => \N__58703\,
            I => \N__58589\
        );

    \I__14671\ : InMux
    port map (
            O => \N__58702\,
            I => \N__58589\
        );

    \I__14670\ : Span4Mux_s2_v
    port map (
            O => \N__58699\,
            I => \N__58586\
        );

    \I__14669\ : InMux
    port map (
            O => \N__58696\,
            I => \N__58571\
        );

    \I__14668\ : InMux
    port map (
            O => \N__58695\,
            I => \N__58571\
        );

    \I__14667\ : InMux
    port map (
            O => \N__58692\,
            I => \N__58571\
        );

    \I__14666\ : InMux
    port map (
            O => \N__58691\,
            I => \N__58571\
        );

    \I__14665\ : InMux
    port map (
            O => \N__58688\,
            I => \N__58571\
        );

    \I__14664\ : InMux
    port map (
            O => \N__58687\,
            I => \N__58571\
        );

    \I__14663\ : InMux
    port map (
            O => \N__58684\,
            I => \N__58571\
        );

    \I__14662\ : InMux
    port map (
            O => \N__58683\,
            I => \N__58554\
        );

    \I__14661\ : InMux
    port map (
            O => \N__58680\,
            I => \N__58554\
        );

    \I__14660\ : InMux
    port map (
            O => \N__58679\,
            I => \N__58554\
        );

    \I__14659\ : InMux
    port map (
            O => \N__58676\,
            I => \N__58554\
        );

    \I__14658\ : InMux
    port map (
            O => \N__58675\,
            I => \N__58554\
        );

    \I__14657\ : InMux
    port map (
            O => \N__58672\,
            I => \N__58554\
        );

    \I__14656\ : InMux
    port map (
            O => \N__58671\,
            I => \N__58554\
        );

    \I__14655\ : InMux
    port map (
            O => \N__58668\,
            I => \N__58554\
        );

    \I__14654\ : InMux
    port map (
            O => \N__58665\,
            I => \N__58539\
        );

    \I__14653\ : InMux
    port map (
            O => \N__58664\,
            I => \N__58539\
        );

    \I__14652\ : InMux
    port map (
            O => \N__58661\,
            I => \N__58539\
        );

    \I__14651\ : InMux
    port map (
            O => \N__58660\,
            I => \N__58539\
        );

    \I__14650\ : InMux
    port map (
            O => \N__58657\,
            I => \N__58539\
        );

    \I__14649\ : InMux
    port map (
            O => \N__58656\,
            I => \N__58539\
        );

    \I__14648\ : InMux
    port map (
            O => \N__58653\,
            I => \N__58539\
        );

    \I__14647\ : Span4Mux_v
    port map (
            O => \N__58644\,
            I => \N__58534\
        );

    \I__14646\ : LocalMux
    port map (
            O => \N__58641\,
            I => \N__58534\
        );

    \I__14645\ : Span4Mux_v
    port map (
            O => \N__58636\,
            I => \N__58525\
        );

    \I__14644\ : LocalMux
    port map (
            O => \N__58633\,
            I => \N__58525\
        );

    \I__14643\ : LocalMux
    port map (
            O => \N__58630\,
            I => \N__58525\
        );

    \I__14642\ : LocalMux
    port map (
            O => \N__58627\,
            I => \N__58525\
        );

    \I__14641\ : InMux
    port map (
            O => \N__58626\,
            I => \N__58508\
        );

    \I__14640\ : InMux
    port map (
            O => \N__58623\,
            I => \N__58508\
        );

    \I__14639\ : InMux
    port map (
            O => \N__58622\,
            I => \N__58508\
        );

    \I__14638\ : InMux
    port map (
            O => \N__58619\,
            I => \N__58508\
        );

    \I__14637\ : InMux
    port map (
            O => \N__58618\,
            I => \N__58508\
        );

    \I__14636\ : InMux
    port map (
            O => \N__58615\,
            I => \N__58508\
        );

    \I__14635\ : InMux
    port map (
            O => \N__58614\,
            I => \N__58508\
        );

    \I__14634\ : InMux
    port map (
            O => \N__58611\,
            I => \N__58508\
        );

    \I__14633\ : Span4Mux_v
    port map (
            O => \N__58608\,
            I => \N__58503\
        );

    \I__14632\ : Span4Mux_h
    port map (
            O => \N__58605\,
            I => \N__58503\
        );

    \I__14631\ : LocalMux
    port map (
            O => \N__58598\,
            I => \N__58498\
        );

    \I__14630\ : LocalMux
    port map (
            O => \N__58589\,
            I => \N__58498\
        );

    \I__14629\ : Sp12to4
    port map (
            O => \N__58586\,
            I => \N__58495\
        );

    \I__14628\ : LocalMux
    port map (
            O => \N__58571\,
            I => \N__58490\
        );

    \I__14627\ : LocalMux
    port map (
            O => \N__58554\,
            I => \N__58490\
        );

    \I__14626\ : LocalMux
    port map (
            O => \N__58539\,
            I => \N__58487\
        );

    \I__14625\ : Span4Mux_v
    port map (
            O => \N__58534\,
            I => \N__58481\
        );

    \I__14624\ : Span4Mux_v
    port map (
            O => \N__58525\,
            I => \N__58481\
        );

    \I__14623\ : LocalMux
    port map (
            O => \N__58508\,
            I => \N__58478\
        );

    \I__14622\ : Span4Mux_h
    port map (
            O => \N__58503\,
            I => \N__58475\
        );

    \I__14621\ : Span4Mux_v
    port map (
            O => \N__58498\,
            I => \N__58472\
        );

    \I__14620\ : Span12Mux_h
    port map (
            O => \N__58495\,
            I => \N__58469\
        );

    \I__14619\ : Span4Mux_v
    port map (
            O => \N__58490\,
            I => \N__58466\
        );

    \I__14618\ : Span4Mux_v
    port map (
            O => \N__58487\,
            I => \N__58463\
        );

    \I__14617\ : SRMux
    port map (
            O => \N__58486\,
            I => \N__58460\
        );

    \I__14616\ : Span4Mux_h
    port map (
            O => \N__58481\,
            I => \N__58455\
        );

    \I__14615\ : Span4Mux_h
    port map (
            O => \N__58478\,
            I => \N__58455\
        );

    \I__14614\ : Span4Mux_h
    port map (
            O => \N__58475\,
            I => \N__58450\
        );

    \I__14613\ : Span4Mux_v
    port map (
            O => \N__58472\,
            I => \N__58450\
        );

    \I__14612\ : Span12Mux_v
    port map (
            O => \N__58469\,
            I => \N__58441\
        );

    \I__14611\ : Sp12to4
    port map (
            O => \N__58466\,
            I => \N__58441\
        );

    \I__14610\ : Sp12to4
    port map (
            O => \N__58463\,
            I => \N__58441\
        );

    \I__14609\ : LocalMux
    port map (
            O => \N__58460\,
            I => \N__58441\
        );

    \I__14608\ : Span4Mux_h
    port map (
            O => \N__58455\,
            I => \N__58438\
        );

    \I__14607\ : Odrv4
    port map (
            O => \N__58450\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14606\ : Odrv12
    port map (
            O => \N__58441\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14605\ : Odrv4
    port map (
            O => \N__58438\,
            I => \CONSTANT_ONE_NET\
        );

    \I__14604\ : InMux
    port map (
            O => \N__58431\,
            I => \N__58427\
        );

    \I__14603\ : InMux
    port map (
            O => \N__58430\,
            I => \N__58424\
        );

    \I__14602\ : LocalMux
    port map (
            O => \N__58427\,
            I => \N__58421\
        );

    \I__14601\ : LocalMux
    port map (
            O => \N__58424\,
            I => \N__58418\
        );

    \I__14600\ : Odrv4
    port map (
            O => \N__58421\,
            I => \comm_spi.n14800\
        );

    \I__14599\ : Odrv4
    port map (
            O => \N__58418\,
            I => \comm_spi.n14800\
        );

    \I__14598\ : ClkMux
    port map (
            O => \N__58413\,
            I => \N__58409\
        );

    \I__14597\ : ClkMux
    port map (
            O => \N__58412\,
            I => \N__58403\
        );

    \I__14596\ : LocalMux
    port map (
            O => \N__58409\,
            I => \N__58396\
        );

    \I__14595\ : ClkMux
    port map (
            O => \N__58408\,
            I => \N__58393\
        );

    \I__14594\ : ClkMux
    port map (
            O => \N__58407\,
            I => \N__58388\
        );

    \I__14593\ : ClkMux
    port map (
            O => \N__58406\,
            I => \N__58385\
        );

    \I__14592\ : LocalMux
    port map (
            O => \N__58403\,
            I => \N__58381\
        );

    \I__14591\ : ClkMux
    port map (
            O => \N__58402\,
            I => \N__58378\
        );

    \I__14590\ : ClkMux
    port map (
            O => \N__58401\,
            I => \N__58375\
        );

    \I__14589\ : ClkMux
    port map (
            O => \N__58400\,
            I => \N__58372\
        );

    \I__14588\ : ClkMux
    port map (
            O => \N__58399\,
            I => \N__58368\
        );

    \I__14587\ : Span4Mux_v
    port map (
            O => \N__58396\,
            I => \N__58362\
        );

    \I__14586\ : LocalMux
    port map (
            O => \N__58393\,
            I => \N__58362\
        );

    \I__14585\ : ClkMux
    port map (
            O => \N__58392\,
            I => \N__58359\
        );

    \I__14584\ : ClkMux
    port map (
            O => \N__58391\,
            I => \N__58353\
        );

    \I__14583\ : LocalMux
    port map (
            O => \N__58388\,
            I => \N__58347\
        );

    \I__14582\ : LocalMux
    port map (
            O => \N__58385\,
            I => \N__58347\
        );

    \I__14581\ : ClkMux
    port map (
            O => \N__58384\,
            I => \N__58344\
        );

    \I__14580\ : Span4Mux_v
    port map (
            O => \N__58381\,
            I => \N__58341\
        );

    \I__14579\ : LocalMux
    port map (
            O => \N__58378\,
            I => \N__58338\
        );

    \I__14578\ : LocalMux
    port map (
            O => \N__58375\,
            I => \N__58332\
        );

    \I__14577\ : LocalMux
    port map (
            O => \N__58372\,
            I => \N__58332\
        );

    \I__14576\ : ClkMux
    port map (
            O => \N__58371\,
            I => \N__58329\
        );

    \I__14575\ : LocalMux
    port map (
            O => \N__58368\,
            I => \N__58325\
        );

    \I__14574\ : ClkMux
    port map (
            O => \N__58367\,
            I => \N__58322\
        );

    \I__14573\ : Span4Mux_v
    port map (
            O => \N__58362\,
            I => \N__58317\
        );

    \I__14572\ : LocalMux
    port map (
            O => \N__58359\,
            I => \N__58317\
        );

    \I__14571\ : ClkMux
    port map (
            O => \N__58358\,
            I => \N__58314\
        );

    \I__14570\ : ClkMux
    port map (
            O => \N__58357\,
            I => \N__58311\
        );

    \I__14569\ : ClkMux
    port map (
            O => \N__58356\,
            I => \N__58308\
        );

    \I__14568\ : LocalMux
    port map (
            O => \N__58353\,
            I => \N__58304\
        );

    \I__14567\ : ClkMux
    port map (
            O => \N__58352\,
            I => \N__58301\
        );

    \I__14566\ : Span4Mux_v
    port map (
            O => \N__58347\,
            I => \N__58298\
        );

    \I__14565\ : LocalMux
    port map (
            O => \N__58344\,
            I => \N__58295\
        );

    \I__14564\ : Span4Mux_h
    port map (
            O => \N__58341\,
            I => \N__58290\
        );

    \I__14563\ : Span4Mux_h
    port map (
            O => \N__58338\,
            I => \N__58290\
        );

    \I__14562\ : ClkMux
    port map (
            O => \N__58337\,
            I => \N__58287\
        );

    \I__14561\ : Span4Mux_v
    port map (
            O => \N__58332\,
            I => \N__58284\
        );

    \I__14560\ : LocalMux
    port map (
            O => \N__58329\,
            I => \N__58281\
        );

    \I__14559\ : ClkMux
    port map (
            O => \N__58328\,
            I => \N__58278\
        );

    \I__14558\ : Span4Mux_h
    port map (
            O => \N__58325\,
            I => \N__58273\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__58322\,
            I => \N__58273\
        );

    \I__14556\ : Span4Mux_h
    port map (
            O => \N__58317\,
            I => \N__58270\
        );

    \I__14555\ : LocalMux
    port map (
            O => \N__58314\,
            I => \N__58267\
        );

    \I__14554\ : LocalMux
    port map (
            O => \N__58311\,
            I => \N__58264\
        );

    \I__14553\ : LocalMux
    port map (
            O => \N__58308\,
            I => \N__58261\
        );

    \I__14552\ : ClkMux
    port map (
            O => \N__58307\,
            I => \N__58258\
        );

    \I__14551\ : Span4Mux_v
    port map (
            O => \N__58304\,
            I => \N__58252\
        );

    \I__14550\ : LocalMux
    port map (
            O => \N__58301\,
            I => \N__58252\
        );

    \I__14549\ : Span4Mux_h
    port map (
            O => \N__58298\,
            I => \N__58243\
        );

    \I__14548\ : Span4Mux_h
    port map (
            O => \N__58295\,
            I => \N__58243\
        );

    \I__14547\ : Span4Mux_v
    port map (
            O => \N__58290\,
            I => \N__58243\
        );

    \I__14546\ : LocalMux
    port map (
            O => \N__58287\,
            I => \N__58243\
        );

    \I__14545\ : Span4Mux_h
    port map (
            O => \N__58284\,
            I => \N__58236\
        );

    \I__14544\ : Span4Mux_h
    port map (
            O => \N__58281\,
            I => \N__58236\
        );

    \I__14543\ : LocalMux
    port map (
            O => \N__58278\,
            I => \N__58236\
        );

    \I__14542\ : Span4Mux_h
    port map (
            O => \N__58273\,
            I => \N__58231\
        );

    \I__14541\ : Span4Mux_v
    port map (
            O => \N__58270\,
            I => \N__58231\
        );

    \I__14540\ : Span4Mux_h
    port map (
            O => \N__58267\,
            I => \N__58222\
        );

    \I__14539\ : Span4Mux_v
    port map (
            O => \N__58264\,
            I => \N__58222\
        );

    \I__14538\ : Span4Mux_v
    port map (
            O => \N__58261\,
            I => \N__58222\
        );

    \I__14537\ : LocalMux
    port map (
            O => \N__58258\,
            I => \N__58222\
        );

    \I__14536\ : ClkMux
    port map (
            O => \N__58257\,
            I => \N__58219\
        );

    \I__14535\ : Span4Mux_v
    port map (
            O => \N__58252\,
            I => \N__58216\
        );

    \I__14534\ : Span4Mux_v
    port map (
            O => \N__58243\,
            I => \N__58211\
        );

    \I__14533\ : Span4Mux_h
    port map (
            O => \N__58236\,
            I => \N__58211\
        );

    \I__14532\ : Span4Mux_v
    port map (
            O => \N__58231\,
            I => \N__58206\
        );

    \I__14531\ : Span4Mux_h
    port map (
            O => \N__58222\,
            I => \N__58206\
        );

    \I__14530\ : LocalMux
    port map (
            O => \N__58219\,
            I => \N__58203\
        );

    \I__14529\ : Odrv4
    port map (
            O => \N__58216\,
            I => \comm_spi.iclk\
        );

    \I__14528\ : Odrv4
    port map (
            O => \N__58211\,
            I => \comm_spi.iclk\
        );

    \I__14527\ : Odrv4
    port map (
            O => \N__58206\,
            I => \comm_spi.iclk\
        );

    \I__14526\ : Odrv12
    port map (
            O => \N__58203\,
            I => \comm_spi.iclk\
        );

    \I__14525\ : InMux
    port map (
            O => \N__58194\,
            I => \N__58187\
        );

    \I__14524\ : InMux
    port map (
            O => \N__58193\,
            I => \N__58187\
        );

    \I__14523\ : InMux
    port map (
            O => \N__58192\,
            I => \N__58184\
        );

    \I__14522\ : LocalMux
    port map (
            O => \N__58187\,
            I => \N__58181\
        );

    \I__14521\ : LocalMux
    port map (
            O => \N__58184\,
            I => \N__58178\
        );

    \I__14520\ : Span4Mux_v
    port map (
            O => \N__58181\,
            I => \N__58173\
        );

    \I__14519\ : Span4Mux_v
    port map (
            O => \N__58178\,
            I => \N__58173\
        );

    \I__14518\ : Sp12to4
    port map (
            O => \N__58173\,
            I => \N__58170\
        );

    \I__14517\ : Odrv12
    port map (
            O => \N__58170\,
            I => comm_tx_buf_0
        );

    \I__14516\ : CascadeMux
    port map (
            O => \N__58167\,
            I => \N__58153\
        );

    \I__14515\ : CascadeMux
    port map (
            O => \N__58166\,
            I => \N__58150\
        );

    \I__14514\ : SRMux
    port map (
            O => \N__58165\,
            I => \N__58146\
        );

    \I__14513\ : InMux
    port map (
            O => \N__58164\,
            I => \N__58140\
        );

    \I__14512\ : InMux
    port map (
            O => \N__58163\,
            I => \N__58140\
        );

    \I__14511\ : CascadeMux
    port map (
            O => \N__58162\,
            I => \N__58136\
        );

    \I__14510\ : CascadeMux
    port map (
            O => \N__58161\,
            I => \N__58133\
        );

    \I__14509\ : CascadeMux
    port map (
            O => \N__58160\,
            I => \N__58128\
        );

    \I__14508\ : InMux
    port map (
            O => \N__58159\,
            I => \N__58123\
        );

    \I__14507\ : InMux
    port map (
            O => \N__58158\,
            I => \N__58117\
        );

    \I__14506\ : InMux
    port map (
            O => \N__58157\,
            I => \N__58114\
        );

    \I__14505\ : CascadeMux
    port map (
            O => \N__58156\,
            I => \N__58110\
        );

    \I__14504\ : InMux
    port map (
            O => \N__58153\,
            I => \N__58101\
        );

    \I__14503\ : InMux
    port map (
            O => \N__58150\,
            I => \N__58101\
        );

    \I__14502\ : InMux
    port map (
            O => \N__58149\,
            I => \N__58101\
        );

    \I__14501\ : LocalMux
    port map (
            O => \N__58146\,
            I => \N__58098\
        );

    \I__14500\ : SRMux
    port map (
            O => \N__58145\,
            I => \N__58095\
        );

    \I__14499\ : LocalMux
    port map (
            O => \N__58140\,
            I => \N__58092\
        );

    \I__14498\ : InMux
    port map (
            O => \N__58139\,
            I => \N__58081\
        );

    \I__14497\ : InMux
    port map (
            O => \N__58136\,
            I => \N__58081\
        );

    \I__14496\ : InMux
    port map (
            O => \N__58133\,
            I => \N__58081\
        );

    \I__14495\ : InMux
    port map (
            O => \N__58132\,
            I => \N__58081\
        );

    \I__14494\ : InMux
    port map (
            O => \N__58131\,
            I => \N__58081\
        );

    \I__14493\ : InMux
    port map (
            O => \N__58128\,
            I => \N__58074\
        );

    \I__14492\ : InMux
    port map (
            O => \N__58127\,
            I => \N__58074\
        );

    \I__14491\ : InMux
    port map (
            O => \N__58126\,
            I => \N__58074\
        );

    \I__14490\ : LocalMux
    port map (
            O => \N__58123\,
            I => \N__58071\
        );

    \I__14489\ : SRMux
    port map (
            O => \N__58122\,
            I => \N__58068\
        );

    \I__14488\ : InMux
    port map (
            O => \N__58121\,
            I => \N__58060\
        );

    \I__14487\ : InMux
    port map (
            O => \N__58120\,
            I => \N__58060\
        );

    \I__14486\ : LocalMux
    port map (
            O => \N__58117\,
            I => \N__58055\
        );

    \I__14485\ : LocalMux
    port map (
            O => \N__58114\,
            I => \N__58048\
        );

    \I__14484\ : InMux
    port map (
            O => \N__58113\,
            I => \N__58045\
        );

    \I__14483\ : InMux
    port map (
            O => \N__58110\,
            I => \N__58038\
        );

    \I__14482\ : InMux
    port map (
            O => \N__58109\,
            I => \N__58038\
        );

    \I__14481\ : InMux
    port map (
            O => \N__58108\,
            I => \N__58038\
        );

    \I__14480\ : LocalMux
    port map (
            O => \N__58101\,
            I => \N__58035\
        );

    \I__14479\ : Span4Mux_v
    port map (
            O => \N__58098\,
            I => \N__58030\
        );

    \I__14478\ : LocalMux
    port map (
            O => \N__58095\,
            I => \N__58030\
        );

    \I__14477\ : Span4Mux_h
    port map (
            O => \N__58092\,
            I => \N__58023\
        );

    \I__14476\ : LocalMux
    port map (
            O => \N__58081\,
            I => \N__58023\
        );

    \I__14475\ : LocalMux
    port map (
            O => \N__58074\,
            I => \N__58023\
        );

    \I__14474\ : Span4Mux_v
    port map (
            O => \N__58071\,
            I => \N__58018\
        );

    \I__14473\ : LocalMux
    port map (
            O => \N__58068\,
            I => \N__58018\
        );

    \I__14472\ : InMux
    port map (
            O => \N__58067\,
            I => \N__58013\
        );

    \I__14471\ : InMux
    port map (
            O => \N__58066\,
            I => \N__58013\
        );

    \I__14470\ : InMux
    port map (
            O => \N__58065\,
            I => \N__58010\
        );

    \I__14469\ : LocalMux
    port map (
            O => \N__58060\,
            I => \N__58007\
        );

    \I__14468\ : InMux
    port map (
            O => \N__58059\,
            I => \N__58002\
        );

    \I__14467\ : InMux
    port map (
            O => \N__58058\,
            I => \N__58002\
        );

    \I__14466\ : Span4Mux_v
    port map (
            O => \N__58055\,
            I => \N__57999\
        );

    \I__14465\ : InMux
    port map (
            O => \N__58054\,
            I => \N__57994\
        );

    \I__14464\ : InMux
    port map (
            O => \N__58053\,
            I => \N__57994\
        );

    \I__14463\ : InMux
    port map (
            O => \N__58052\,
            I => \N__57989\
        );

    \I__14462\ : InMux
    port map (
            O => \N__58051\,
            I => \N__57989\
        );

    \I__14461\ : Span4Mux_h
    port map (
            O => \N__58048\,
            I => \N__57982\
        );

    \I__14460\ : LocalMux
    port map (
            O => \N__58045\,
            I => \N__57982\
        );

    \I__14459\ : LocalMux
    port map (
            O => \N__58038\,
            I => \N__57979\
        );

    \I__14458\ : Span4Mux_v
    port map (
            O => \N__58035\,
            I => \N__57976\
        );

    \I__14457\ : Span4Mux_h
    port map (
            O => \N__58030\,
            I => \N__57973\
        );

    \I__14456\ : Span4Mux_v
    port map (
            O => \N__58023\,
            I => \N__57970\
        );

    \I__14455\ : Span4Mux_v
    port map (
            O => \N__58018\,
            I => \N__57967\
        );

    \I__14454\ : LocalMux
    port map (
            O => \N__58013\,
            I => \N__57960\
        );

    \I__14453\ : LocalMux
    port map (
            O => \N__58010\,
            I => \N__57960\
        );

    \I__14452\ : Span12Mux_s10_v
    port map (
            O => \N__58007\,
            I => \N__57960\
        );

    \I__14451\ : LocalMux
    port map (
            O => \N__58002\,
            I => \N__57957\
        );

    \I__14450\ : Sp12to4
    port map (
            O => \N__57999\,
            I => \N__57950\
        );

    \I__14449\ : LocalMux
    port map (
            O => \N__57994\,
            I => \N__57950\
        );

    \I__14448\ : LocalMux
    port map (
            O => \N__57989\,
            I => \N__57950\
        );

    \I__14447\ : InMux
    port map (
            O => \N__57988\,
            I => \N__57945\
        );

    \I__14446\ : InMux
    port map (
            O => \N__57987\,
            I => \N__57945\
        );

    \I__14445\ : Span4Mux_h
    port map (
            O => \N__57982\,
            I => \N__57940\
        );

    \I__14444\ : Span4Mux_v
    port map (
            O => \N__57979\,
            I => \N__57940\
        );

    \I__14443\ : Span4Mux_h
    port map (
            O => \N__57976\,
            I => \N__57935\
        );

    \I__14442\ : Span4Mux_v
    port map (
            O => \N__57973\,
            I => \N__57935\
        );

    \I__14441\ : Span4Mux_v
    port map (
            O => \N__57970\,
            I => \N__57932\
        );

    \I__14440\ : Span4Mux_v
    port map (
            O => \N__57967\,
            I => \N__57929\
        );

    \I__14439\ : Span12Mux_v
    port map (
            O => \N__57960\,
            I => \N__57926\
        );

    \I__14438\ : Span12Mux_h
    port map (
            O => \N__57957\,
            I => \N__57919\
        );

    \I__14437\ : Span12Mux_s11_h
    port map (
            O => \N__57950\,
            I => \N__57919\
        );

    \I__14436\ : LocalMux
    port map (
            O => \N__57945\,
            I => \N__57919\
        );

    \I__14435\ : Span4Mux_v
    port map (
            O => \N__57940\,
            I => \N__57916\
        );

    \I__14434\ : Odrv4
    port map (
            O => \N__57935\,
            I => comm_clear
        );

    \I__14433\ : Odrv4
    port map (
            O => \N__57932\,
            I => comm_clear
        );

    \I__14432\ : Odrv4
    port map (
            O => \N__57929\,
            I => comm_clear
        );

    \I__14431\ : Odrv12
    port map (
            O => \N__57926\,
            I => comm_clear
        );

    \I__14430\ : Odrv12
    port map (
            O => \N__57919\,
            I => comm_clear
        );

    \I__14429\ : Odrv4
    port map (
            O => \N__57916\,
            I => comm_clear
        );

    \I__14428\ : SRMux
    port map (
            O => \N__57903\,
            I => \N__57900\
        );

    \I__14427\ : LocalMux
    port map (
            O => \N__57900\,
            I => \comm_spi.data_tx_7__N_813\
        );

    \I__14426\ : InMux
    port map (
            O => \N__57897\,
            I => \N__57893\
        );

    \I__14425\ : InMux
    port map (
            O => \N__57896\,
            I => \N__57890\
        );

    \I__14424\ : LocalMux
    port map (
            O => \N__57893\,
            I => \N__57887\
        );

    \I__14423\ : LocalMux
    port map (
            O => \N__57890\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__14422\ : Odrv4
    port map (
            O => \N__57887\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__14421\ : InMux
    port map (
            O => \N__57882\,
            I => \bfn_22_8_0_\
        );

    \I__14420\ : CascadeMux
    port map (
            O => \N__57879\,
            I => \N__57875\
        );

    \I__14419\ : InMux
    port map (
            O => \N__57878\,
            I => \N__57872\
        );

    \I__14418\ : InMux
    port map (
            O => \N__57875\,
            I => \N__57869\
        );

    \I__14417\ : LocalMux
    port map (
            O => \N__57872\,
            I => \N__57866\
        );

    \I__14416\ : LocalMux
    port map (
            O => \N__57869\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__14415\ : Odrv4
    port map (
            O => \N__57866\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__14414\ : InMux
    port map (
            O => \N__57861\,
            I => \ADC_VDC.genclk.n19911\
        );

    \I__14413\ : InMux
    port map (
            O => \N__57858\,
            I => \N__57855\
        );

    \I__14412\ : LocalMux
    port map (
            O => \N__57855\,
            I => \N__57851\
        );

    \I__14411\ : InMux
    port map (
            O => \N__57854\,
            I => \N__57848\
        );

    \I__14410\ : Span4Mux_h
    port map (
            O => \N__57851\,
            I => \N__57845\
        );

    \I__14409\ : LocalMux
    port map (
            O => \N__57848\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__14408\ : Odrv4
    port map (
            O => \N__57845\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__14407\ : InMux
    port map (
            O => \N__57840\,
            I => \ADC_VDC.genclk.n19912\
        );

    \I__14406\ : CascadeMux
    port map (
            O => \N__57837\,
            I => \N__57833\
        );

    \I__14405\ : InMux
    port map (
            O => \N__57836\,
            I => \N__57830\
        );

    \I__14404\ : InMux
    port map (
            O => \N__57833\,
            I => \N__57827\
        );

    \I__14403\ : LocalMux
    port map (
            O => \N__57830\,
            I => \N__57824\
        );

    \I__14402\ : LocalMux
    port map (
            O => \N__57827\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__14401\ : Odrv4
    port map (
            O => \N__57824\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__14400\ : InMux
    port map (
            O => \N__57819\,
            I => \ADC_VDC.genclk.n19913\
        );

    \I__14399\ : InMux
    port map (
            O => \N__57816\,
            I => \N__57813\
        );

    \I__14398\ : LocalMux
    port map (
            O => \N__57813\,
            I => \N__57809\
        );

    \I__14397\ : InMux
    port map (
            O => \N__57812\,
            I => \N__57806\
        );

    \I__14396\ : Span4Mux_h
    port map (
            O => \N__57809\,
            I => \N__57803\
        );

    \I__14395\ : LocalMux
    port map (
            O => \N__57806\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__14394\ : Odrv4
    port map (
            O => \N__57803\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__14393\ : InMux
    port map (
            O => \N__57798\,
            I => \ADC_VDC.genclk.n19914\
        );

    \I__14392\ : CascadeMux
    port map (
            O => \N__57795\,
            I => \N__57791\
        );

    \I__14391\ : InMux
    port map (
            O => \N__57794\,
            I => \N__57788\
        );

    \I__14390\ : InMux
    port map (
            O => \N__57791\,
            I => \N__57785\
        );

    \I__14389\ : LocalMux
    port map (
            O => \N__57788\,
            I => \N__57782\
        );

    \I__14388\ : LocalMux
    port map (
            O => \N__57785\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__14387\ : Odrv4
    port map (
            O => \N__57782\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__14386\ : InMux
    port map (
            O => \N__57777\,
            I => \ADC_VDC.genclk.n19915\
        );

    \I__14385\ : InMux
    port map (
            O => \N__57774\,
            I => \N__57770\
        );

    \I__14384\ : InMux
    port map (
            O => \N__57773\,
            I => \N__57767\
        );

    \I__14383\ : LocalMux
    port map (
            O => \N__57770\,
            I => \N__57764\
        );

    \I__14382\ : LocalMux
    port map (
            O => \N__57767\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__14381\ : Odrv4
    port map (
            O => \N__57764\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__14380\ : InMux
    port map (
            O => \N__57759\,
            I => \ADC_VDC.genclk.n19916\
        );

    \I__14379\ : InMux
    port map (
            O => \N__57756\,
            I => \ADC_VDC.genclk.n19917\
        );

    \I__14378\ : CascadeMux
    port map (
            O => \N__57753\,
            I => \N__57750\
        );

    \I__14377\ : InMux
    port map (
            O => \N__57750\,
            I => \N__57746\
        );

    \I__14376\ : InMux
    port map (
            O => \N__57749\,
            I => \N__57743\
        );

    \I__14375\ : LocalMux
    port map (
            O => \N__57746\,
            I => \N__57740\
        );

    \I__14374\ : LocalMux
    port map (
            O => \N__57743\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__14373\ : Odrv4
    port map (
            O => \N__57740\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__14372\ : CEMux
    port map (
            O => \N__57735\,
            I => \N__57731\
        );

    \I__14371\ : CEMux
    port map (
            O => \N__57734\,
            I => \N__57728\
        );

    \I__14370\ : LocalMux
    port map (
            O => \N__57731\,
            I => \N__57725\
        );

    \I__14369\ : LocalMux
    port map (
            O => \N__57728\,
            I => \N__57722\
        );

    \I__14368\ : Span4Mux_h
    port map (
            O => \N__57725\,
            I => \N__57719\
        );

    \I__14367\ : Odrv4
    port map (
            O => \N__57722\,
            I => \ADC_VDC.genclk.div_state_1__N_1432\
        );

    \I__14366\ : Odrv4
    port map (
            O => \N__57719\,
            I => \ADC_VDC.genclk.div_state_1__N_1432\
        );

    \I__14365\ : InMux
    port map (
            O => \N__57714\,
            I => \N__57710\
        );

    \I__14364\ : InMux
    port map (
            O => \N__57713\,
            I => \N__57707\
        );

    \I__14363\ : LocalMux
    port map (
            O => \N__57710\,
            I => \N__57704\
        );

    \I__14362\ : LocalMux
    port map (
            O => \N__57707\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__14361\ : Odrv4
    port map (
            O => \N__57704\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__14360\ : InMux
    port map (
            O => \N__57699\,
            I => \bfn_22_7_0_\
        );

    \I__14359\ : InMux
    port map (
            O => \N__57696\,
            I => \N__57692\
        );

    \I__14358\ : InMux
    port map (
            O => \N__57695\,
            I => \N__57689\
        );

    \I__14357\ : LocalMux
    port map (
            O => \N__57692\,
            I => \N__57686\
        );

    \I__14356\ : LocalMux
    port map (
            O => \N__57689\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__14355\ : Odrv4
    port map (
            O => \N__57686\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__14354\ : InMux
    port map (
            O => \N__57681\,
            I => \ADC_VDC.genclk.n19903\
        );

    \I__14353\ : CascadeMux
    port map (
            O => \N__57678\,
            I => \N__57674\
        );

    \I__14352\ : InMux
    port map (
            O => \N__57677\,
            I => \N__57671\
        );

    \I__14351\ : InMux
    port map (
            O => \N__57674\,
            I => \N__57668\
        );

    \I__14350\ : LocalMux
    port map (
            O => \N__57671\,
            I => \N__57665\
        );

    \I__14349\ : LocalMux
    port map (
            O => \N__57668\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__14348\ : Odrv4
    port map (
            O => \N__57665\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__14347\ : InMux
    port map (
            O => \N__57660\,
            I => \ADC_VDC.genclk.n19904\
        );

    \I__14346\ : InMux
    port map (
            O => \N__57657\,
            I => \N__57654\
        );

    \I__14345\ : LocalMux
    port map (
            O => \N__57654\,
            I => \N__57650\
        );

    \I__14344\ : InMux
    port map (
            O => \N__57653\,
            I => \N__57647\
        );

    \I__14343\ : Span4Mux_h
    port map (
            O => \N__57650\,
            I => \N__57644\
        );

    \I__14342\ : LocalMux
    port map (
            O => \N__57647\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__14341\ : Odrv4
    port map (
            O => \N__57644\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__14340\ : InMux
    port map (
            O => \N__57639\,
            I => \ADC_VDC.genclk.n19905\
        );

    \I__14339\ : CascadeMux
    port map (
            O => \N__57636\,
            I => \N__57632\
        );

    \I__14338\ : CascadeMux
    port map (
            O => \N__57635\,
            I => \N__57629\
        );

    \I__14337\ : InMux
    port map (
            O => \N__57632\,
            I => \N__57626\
        );

    \I__14336\ : InMux
    port map (
            O => \N__57629\,
            I => \N__57623\
        );

    \I__14335\ : LocalMux
    port map (
            O => \N__57626\,
            I => \N__57620\
        );

    \I__14334\ : LocalMux
    port map (
            O => \N__57623\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__14333\ : Odrv4
    port map (
            O => \N__57620\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__14332\ : InMux
    port map (
            O => \N__57615\,
            I => \ADC_VDC.genclk.n19906\
        );

    \I__14331\ : CascadeMux
    port map (
            O => \N__57612\,
            I => \N__57609\
        );

    \I__14330\ : InMux
    port map (
            O => \N__57609\,
            I => \N__57606\
        );

    \I__14329\ : LocalMux
    port map (
            O => \N__57606\,
            I => \N__57602\
        );

    \I__14328\ : InMux
    port map (
            O => \N__57605\,
            I => \N__57599\
        );

    \I__14327\ : Span4Mux_v
    port map (
            O => \N__57602\,
            I => \N__57596\
        );

    \I__14326\ : LocalMux
    port map (
            O => \N__57599\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__14325\ : Odrv4
    port map (
            O => \N__57596\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__14324\ : InMux
    port map (
            O => \N__57591\,
            I => \ADC_VDC.genclk.n19907\
        );

    \I__14323\ : CascadeMux
    port map (
            O => \N__57588\,
            I => \N__57584\
        );

    \I__14322\ : InMux
    port map (
            O => \N__57587\,
            I => \N__57581\
        );

    \I__14321\ : InMux
    port map (
            O => \N__57584\,
            I => \N__57578\
        );

    \I__14320\ : LocalMux
    port map (
            O => \N__57581\,
            I => \N__57575\
        );

    \I__14319\ : LocalMux
    port map (
            O => \N__57578\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__14318\ : Odrv4
    port map (
            O => \N__57575\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__14317\ : InMux
    port map (
            O => \N__57570\,
            I => \ADC_VDC.genclk.n19908\
        );

    \I__14316\ : CascadeMux
    port map (
            O => \N__57567\,
            I => \N__57564\
        );

    \I__14315\ : InMux
    port map (
            O => \N__57564\,
            I => \N__57560\
        );

    \I__14314\ : InMux
    port map (
            O => \N__57563\,
            I => \N__57557\
        );

    \I__14313\ : LocalMux
    port map (
            O => \N__57560\,
            I => \N__57554\
        );

    \I__14312\ : LocalMux
    port map (
            O => \N__57557\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__14311\ : Odrv4
    port map (
            O => \N__57554\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__14310\ : InMux
    port map (
            O => \N__57549\,
            I => \ADC_VDC.genclk.n19909\
        );

    \I__14309\ : SRMux
    port map (
            O => \N__57546\,
            I => \N__57543\
        );

    \I__14308\ : LocalMux
    port map (
            O => \N__57543\,
            I => \N__57540\
        );

    \I__14307\ : Odrv12
    port map (
            O => \N__57540\,
            I => \comm_spi.data_tx_7__N_829\
        );

    \I__14306\ : InMux
    port map (
            O => \N__57537\,
            I => \N__57532\
        );

    \I__14305\ : InMux
    port map (
            O => \N__57536\,
            I => \N__57529\
        );

    \I__14304\ : InMux
    port map (
            O => \N__57535\,
            I => \N__57526\
        );

    \I__14303\ : LocalMux
    port map (
            O => \N__57532\,
            I => \comm_spi.n23098\
        );

    \I__14302\ : LocalMux
    port map (
            O => \N__57529\,
            I => \comm_spi.n23098\
        );

    \I__14301\ : LocalMux
    port map (
            O => \N__57526\,
            I => \comm_spi.n23098\
        );

    \I__14300\ : InMux
    port map (
            O => \N__57519\,
            I => \N__57516\
        );

    \I__14299\ : LocalMux
    port map (
            O => \N__57516\,
            I => \N__57512\
        );

    \I__14298\ : InMux
    port map (
            O => \N__57515\,
            I => \N__57509\
        );

    \I__14297\ : Span4Mux_v
    port map (
            O => \N__57512\,
            I => \N__57506\
        );

    \I__14296\ : LocalMux
    port map (
            O => \N__57509\,
            I => \N__57503\
        );

    \I__14295\ : Span4Mux_h
    port map (
            O => \N__57506\,
            I => \N__57500\
        );

    \I__14294\ : Span4Mux_v
    port map (
            O => \N__57503\,
            I => \N__57497\
        );

    \I__14293\ : Odrv4
    port map (
            O => \N__57500\,
            I => \comm_spi.n14838\
        );

    \I__14292\ : Odrv4
    port map (
            O => \N__57497\,
            I => \comm_spi.n14838\
        );

    \I__14291\ : InMux
    port map (
            O => \N__57492\,
            I => \N__57488\
        );

    \I__14290\ : InMux
    port map (
            O => \N__57491\,
            I => \N__57485\
        );

    \I__14289\ : LocalMux
    port map (
            O => \N__57488\,
            I => \N__57482\
        );

    \I__14288\ : LocalMux
    port map (
            O => \N__57485\,
            I => \N__57479\
        );

    \I__14287\ : Odrv4
    port map (
            O => \N__57482\,
            I => \comm_spi.n14839\
        );

    \I__14286\ : Odrv12
    port map (
            O => \N__57479\,
            I => \comm_spi.n14839\
        );

    \I__14285\ : InMux
    port map (
            O => \N__57474\,
            I => \N__57471\
        );

    \I__14284\ : LocalMux
    port map (
            O => \N__57471\,
            I => \N__57467\
        );

    \I__14283\ : InMux
    port map (
            O => \N__57470\,
            I => \N__57464\
        );

    \I__14282\ : Span4Mux_v
    port map (
            O => \N__57467\,
            I => \N__57459\
        );

    \I__14281\ : LocalMux
    port map (
            O => \N__57464\,
            I => \N__57459\
        );

    \I__14280\ : Span4Mux_h
    port map (
            O => \N__57459\,
            I => \N__57456\
        );

    \I__14279\ : Span4Mux_h
    port map (
            O => \N__57456\,
            I => \N__57453\
        );

    \I__14278\ : Odrv4
    port map (
            O => \N__57453\,
            I => \comm_spi.n14843\
        );

    \I__14277\ : SRMux
    port map (
            O => \N__57450\,
            I => \N__57447\
        );

    \I__14276\ : LocalMux
    port map (
            O => \N__57447\,
            I => \N__57444\
        );

    \I__14275\ : Odrv4
    port map (
            O => \N__57444\,
            I => \comm_spi.data_tx_7__N_820\
        );

    \I__14274\ : InMux
    port map (
            O => \N__57441\,
            I => \N__57438\
        );

    \I__14273\ : LocalMux
    port map (
            O => \N__57438\,
            I => \N__57434\
        );

    \I__14272\ : InMux
    port map (
            O => \N__57437\,
            I => \N__57431\
        );

    \I__14271\ : Sp12to4
    port map (
            O => \N__57434\,
            I => \N__57425\
        );

    \I__14270\ : LocalMux
    port map (
            O => \N__57431\,
            I => \N__57425\
        );

    \I__14269\ : InMux
    port map (
            O => \N__57430\,
            I => \N__57422\
        );

    \I__14268\ : Odrv12
    port map (
            O => \N__57425\,
            I => \comm_spi.n23104\
        );

    \I__14267\ : LocalMux
    port map (
            O => \N__57422\,
            I => \comm_spi.n23104\
        );

    \I__14266\ : InMux
    port map (
            O => \N__57417\,
            I => \N__57414\
        );

    \I__14265\ : LocalMux
    port map (
            O => \N__57414\,
            I => \N__57410\
        );

    \I__14264\ : InMux
    port map (
            O => \N__57413\,
            I => \N__57407\
        );

    \I__14263\ : Sp12to4
    port map (
            O => \N__57410\,
            I => \N__57402\
        );

    \I__14262\ : LocalMux
    port map (
            O => \N__57407\,
            I => \N__57402\
        );

    \I__14261\ : Odrv12
    port map (
            O => \N__57402\,
            I => \comm_spi.n14830\
        );

    \I__14260\ : InMux
    port map (
            O => \N__57399\,
            I => \N__57396\
        );

    \I__14259\ : LocalMux
    port map (
            O => \N__57396\,
            I => \N__57392\
        );

    \I__14258\ : InMux
    port map (
            O => \N__57395\,
            I => \N__57389\
        );

    \I__14257\ : Span4Mux_v
    port map (
            O => \N__57392\,
            I => \N__57386\
        );

    \I__14256\ : LocalMux
    port map (
            O => \N__57389\,
            I => \N__57383\
        );

    \I__14255\ : Odrv4
    port map (
            O => \N__57386\,
            I => \comm_spi.n14831\
        );

    \I__14254\ : Odrv4
    port map (
            O => \N__57383\,
            I => \comm_spi.n14831\
        );

    \I__14253\ : InMux
    port map (
            O => \N__57378\,
            I => \N__57375\
        );

    \I__14252\ : LocalMux
    port map (
            O => \N__57375\,
            I => \N__57372\
        );

    \I__14251\ : Span4Mux_h
    port map (
            O => \N__57372\,
            I => \N__57368\
        );

    \I__14250\ : InMux
    port map (
            O => \N__57371\,
            I => \N__57365\
        );

    \I__14249\ : Span4Mux_v
    port map (
            O => \N__57368\,
            I => \N__57362\
        );

    \I__14248\ : LocalMux
    port map (
            O => \N__57365\,
            I => \N__57359\
        );

    \I__14247\ : Odrv4
    port map (
            O => \N__57362\,
            I => \comm_spi.n14835\
        );

    \I__14246\ : Odrv12
    port map (
            O => \N__57359\,
            I => \comm_spi.n14835\
        );

    \I__14245\ : SRMux
    port map (
            O => \N__57354\,
            I => \N__57351\
        );

    \I__14244\ : LocalMux
    port map (
            O => \N__57351\,
            I => \N__57348\
        );

    \I__14243\ : Span4Mux_h
    port map (
            O => \N__57348\,
            I => \N__57345\
        );

    \I__14242\ : Odrv4
    port map (
            O => \N__57345\,
            I => \comm_spi.data_tx_7__N_826\
        );

    \I__14241\ : InMux
    port map (
            O => \N__57342\,
            I => \N__57339\
        );

    \I__14240\ : LocalMux
    port map (
            O => \N__57339\,
            I => buf_data_iac_13
        );

    \I__14239\ : InMux
    port map (
            O => \N__57336\,
            I => \N__57333\
        );

    \I__14238\ : LocalMux
    port map (
            O => \N__57333\,
            I => \N__57330\
        );

    \I__14237\ : Span12Mux_h
    port map (
            O => \N__57330\,
            I => \N__57327\
        );

    \I__14236\ : Odrv12
    port map (
            O => \N__57327\,
            I => n21456
        );

    \I__14235\ : InMux
    port map (
            O => \N__57324\,
            I => \N__57321\
        );

    \I__14234\ : LocalMux
    port map (
            O => \N__57321\,
            I => buf_data_iac_12
        );

    \I__14233\ : InMux
    port map (
            O => \N__57318\,
            I => \N__57315\
        );

    \I__14232\ : LocalMux
    port map (
            O => \N__57315\,
            I => \N__57312\
        );

    \I__14231\ : Span4Mux_h
    port map (
            O => \N__57312\,
            I => \N__57309\
        );

    \I__14230\ : Span4Mux_h
    port map (
            O => \N__57309\,
            I => \N__57306\
        );

    \I__14229\ : Span4Mux_h
    port map (
            O => \N__57306\,
            I => \N__57303\
        );

    \I__14228\ : Odrv4
    port map (
            O => \N__57303\,
            I => n21447
        );

    \I__14227\ : InMux
    port map (
            O => \N__57300\,
            I => \N__57297\
        );

    \I__14226\ : LocalMux
    port map (
            O => \N__57297\,
            I => \N__57294\
        );

    \I__14225\ : Odrv4
    port map (
            O => \N__57294\,
            I => buf_data_iac_9
        );

    \I__14224\ : InMux
    port map (
            O => \N__57291\,
            I => \N__57288\
        );

    \I__14223\ : LocalMux
    port map (
            O => \N__57288\,
            I => \N__57285\
        );

    \I__14222\ : Span4Mux_h
    port map (
            O => \N__57285\,
            I => \N__57282\
        );

    \I__14221\ : Odrv4
    port map (
            O => \N__57282\,
            I => n21512
        );

    \I__14220\ : InMux
    port map (
            O => \N__57279\,
            I => \N__57276\
        );

    \I__14219\ : LocalMux
    port map (
            O => \N__57276\,
            I => buf_data_iac_11
        );

    \I__14218\ : CascadeMux
    port map (
            O => \N__57273\,
            I => \N__57254\
        );

    \I__14217\ : InMux
    port map (
            O => \N__57272\,
            I => \N__57246\
        );

    \I__14216\ : InMux
    port map (
            O => \N__57271\,
            I => \N__57243\
        );

    \I__14215\ : InMux
    port map (
            O => \N__57270\,
            I => \N__57240\
        );

    \I__14214\ : InMux
    port map (
            O => \N__57269\,
            I => \N__57233\
        );

    \I__14213\ : InMux
    port map (
            O => \N__57268\,
            I => \N__57233\
        );

    \I__14212\ : InMux
    port map (
            O => \N__57267\,
            I => \N__57230\
        );

    \I__14211\ : InMux
    port map (
            O => \N__57266\,
            I => \N__57227\
        );

    \I__14210\ : InMux
    port map (
            O => \N__57265\,
            I => \N__57224\
        );

    \I__14209\ : InMux
    port map (
            O => \N__57264\,
            I => \N__57221\
        );

    \I__14208\ : InMux
    port map (
            O => \N__57263\,
            I => \N__57218\
        );

    \I__14207\ : CascadeMux
    port map (
            O => \N__57262\,
            I => \N__57214\
        );

    \I__14206\ : CascadeMux
    port map (
            O => \N__57261\,
            I => \N__57199\
        );

    \I__14205\ : InMux
    port map (
            O => \N__57260\,
            I => \N__57191\
        );

    \I__14204\ : CascadeMux
    port map (
            O => \N__57259\,
            I => \N__57188\
        );

    \I__14203\ : CascadeMux
    port map (
            O => \N__57258\,
            I => \N__57181\
        );

    \I__14202\ : InMux
    port map (
            O => \N__57257\,
            I => \N__57170\
        );

    \I__14201\ : InMux
    port map (
            O => \N__57254\,
            I => \N__57170\
        );

    \I__14200\ : InMux
    port map (
            O => \N__57253\,
            I => \N__57170\
        );

    \I__14199\ : InMux
    port map (
            O => \N__57252\,
            I => \N__57170\
        );

    \I__14198\ : InMux
    port map (
            O => \N__57251\,
            I => \N__57167\
        );

    \I__14197\ : InMux
    port map (
            O => \N__57250\,
            I => \N__57164\
        );

    \I__14196\ : CascadeMux
    port map (
            O => \N__57249\,
            I => \N__57159\
        );

    \I__14195\ : LocalMux
    port map (
            O => \N__57246\,
            I => \N__57152\
        );

    \I__14194\ : LocalMux
    port map (
            O => \N__57243\,
            I => \N__57152\
        );

    \I__14193\ : LocalMux
    port map (
            O => \N__57240\,
            I => \N__57152\
        );

    \I__14192\ : InMux
    port map (
            O => \N__57239\,
            I => \N__57143\
        );

    \I__14191\ : InMux
    port map (
            O => \N__57238\,
            I => \N__57140\
        );

    \I__14190\ : LocalMux
    port map (
            O => \N__57233\,
            I => \N__57137\
        );

    \I__14189\ : LocalMux
    port map (
            O => \N__57230\,
            I => \N__57122\
        );

    \I__14188\ : LocalMux
    port map (
            O => \N__57227\,
            I => \N__57122\
        );

    \I__14187\ : LocalMux
    port map (
            O => \N__57224\,
            I => \N__57115\
        );

    \I__14186\ : LocalMux
    port map (
            O => \N__57221\,
            I => \N__57115\
        );

    \I__14185\ : LocalMux
    port map (
            O => \N__57218\,
            I => \N__57115\
        );

    \I__14184\ : CascadeMux
    port map (
            O => \N__57217\,
            I => \N__57106\
        );

    \I__14183\ : InMux
    port map (
            O => \N__57214\,
            I => \N__57102\
        );

    \I__14182\ : InMux
    port map (
            O => \N__57213\,
            I => \N__57094\
        );

    \I__14181\ : InMux
    port map (
            O => \N__57212\,
            I => \N__57088\
        );

    \I__14180\ : InMux
    port map (
            O => \N__57211\,
            I => \N__57083\
        );

    \I__14179\ : InMux
    port map (
            O => \N__57210\,
            I => \N__57083\
        );

    \I__14178\ : CascadeMux
    port map (
            O => \N__57209\,
            I => \N__57080\
        );

    \I__14177\ : InMux
    port map (
            O => \N__57208\,
            I => \N__57077\
        );

    \I__14176\ : InMux
    port map (
            O => \N__57207\,
            I => \N__57072\
        );

    \I__14175\ : InMux
    port map (
            O => \N__57206\,
            I => \N__57072\
        );

    \I__14174\ : InMux
    port map (
            O => \N__57205\,
            I => \N__57067\
        );

    \I__14173\ : InMux
    port map (
            O => \N__57204\,
            I => \N__57067\
        );

    \I__14172\ : InMux
    port map (
            O => \N__57203\,
            I => \N__57062\
        );

    \I__14171\ : InMux
    port map (
            O => \N__57202\,
            I => \N__57062\
        );

    \I__14170\ : InMux
    port map (
            O => \N__57199\,
            I => \N__57059\
        );

    \I__14169\ : InMux
    port map (
            O => \N__57198\,
            I => \N__57052\
        );

    \I__14168\ : InMux
    port map (
            O => \N__57197\,
            I => \N__57052\
        );

    \I__14167\ : InMux
    port map (
            O => \N__57196\,
            I => \N__57052\
        );

    \I__14166\ : InMux
    port map (
            O => \N__57195\,
            I => \N__57049\
        );

    \I__14165\ : InMux
    port map (
            O => \N__57194\,
            I => \N__57046\
        );

    \I__14164\ : LocalMux
    port map (
            O => \N__57191\,
            I => \N__57043\
        );

    \I__14163\ : InMux
    port map (
            O => \N__57188\,
            I => \N__57038\
        );

    \I__14162\ : InMux
    port map (
            O => \N__57187\,
            I => \N__57038\
        );

    \I__14161\ : InMux
    port map (
            O => \N__57186\,
            I => \N__57035\
        );

    \I__14160\ : InMux
    port map (
            O => \N__57185\,
            I => \N__57032\
        );

    \I__14159\ : InMux
    port map (
            O => \N__57184\,
            I => \N__57029\
        );

    \I__14158\ : InMux
    port map (
            O => \N__57181\,
            I => \N__57018\
        );

    \I__14157\ : InMux
    port map (
            O => \N__57180\,
            I => \N__57018\
        );

    \I__14156\ : InMux
    port map (
            O => \N__57179\,
            I => \N__57015\
        );

    \I__14155\ : LocalMux
    port map (
            O => \N__57170\,
            I => \N__57012\
        );

    \I__14154\ : LocalMux
    port map (
            O => \N__57167\,
            I => \N__57007\
        );

    \I__14153\ : LocalMux
    port map (
            O => \N__57164\,
            I => \N__57007\
        );

    \I__14152\ : InMux
    port map (
            O => \N__57163\,
            I => \N__57004\
        );

    \I__14151\ : InMux
    port map (
            O => \N__57162\,
            I => \N__56999\
        );

    \I__14150\ : InMux
    port map (
            O => \N__57159\,
            I => \N__56999\
        );

    \I__14149\ : Span4Mux_v
    port map (
            O => \N__57152\,
            I => \N__56996\
        );

    \I__14148\ : InMux
    port map (
            O => \N__57151\,
            I => \N__56993\
        );

    \I__14147\ : InMux
    port map (
            O => \N__57150\,
            I => \N__56986\
        );

    \I__14146\ : InMux
    port map (
            O => \N__57149\,
            I => \N__56986\
        );

    \I__14145\ : InMux
    port map (
            O => \N__57148\,
            I => \N__56986\
        );

    \I__14144\ : InMux
    port map (
            O => \N__57147\,
            I => \N__56983\
        );

    \I__14143\ : InMux
    port map (
            O => \N__57146\,
            I => \N__56980\
        );

    \I__14142\ : LocalMux
    port map (
            O => \N__57143\,
            I => \N__56975\
        );

    \I__14141\ : LocalMux
    port map (
            O => \N__57140\,
            I => \N__56975\
        );

    \I__14140\ : Span4Mux_h
    port map (
            O => \N__57137\,
            I => \N__56972\
        );

    \I__14139\ : InMux
    port map (
            O => \N__57136\,
            I => \N__56961\
        );

    \I__14138\ : InMux
    port map (
            O => \N__57135\,
            I => \N__56961\
        );

    \I__14137\ : InMux
    port map (
            O => \N__57134\,
            I => \N__56961\
        );

    \I__14136\ : InMux
    port map (
            O => \N__57133\,
            I => \N__56961\
        );

    \I__14135\ : InMux
    port map (
            O => \N__57132\,
            I => \N__56961\
        );

    \I__14134\ : InMux
    port map (
            O => \N__57131\,
            I => \N__56954\
        );

    \I__14133\ : InMux
    port map (
            O => \N__57130\,
            I => \N__56949\
        );

    \I__14132\ : InMux
    port map (
            O => \N__57129\,
            I => \N__56949\
        );

    \I__14131\ : InMux
    port map (
            O => \N__57128\,
            I => \N__56946\
        );

    \I__14130\ : InMux
    port map (
            O => \N__57127\,
            I => \N__56943\
        );

    \I__14129\ : Span4Mux_v
    port map (
            O => \N__57122\,
            I => \N__56938\
        );

    \I__14128\ : Span4Mux_v
    port map (
            O => \N__57115\,
            I => \N__56938\
        );

    \I__14127\ : InMux
    port map (
            O => \N__57114\,
            I => \N__56934\
        );

    \I__14126\ : InMux
    port map (
            O => \N__57113\,
            I => \N__56931\
        );

    \I__14125\ : InMux
    port map (
            O => \N__57112\,
            I => \N__56928\
        );

    \I__14124\ : InMux
    port map (
            O => \N__57111\,
            I => \N__56925\
        );

    \I__14123\ : InMux
    port map (
            O => \N__57110\,
            I => \N__56918\
        );

    \I__14122\ : InMux
    port map (
            O => \N__57109\,
            I => \N__56918\
        );

    \I__14121\ : InMux
    port map (
            O => \N__57106\,
            I => \N__56918\
        );

    \I__14120\ : InMux
    port map (
            O => \N__57105\,
            I => \N__56915\
        );

    \I__14119\ : LocalMux
    port map (
            O => \N__57102\,
            I => \N__56910\
        );

    \I__14118\ : InMux
    port map (
            O => \N__57101\,
            I => \N__56901\
        );

    \I__14117\ : InMux
    port map (
            O => \N__57100\,
            I => \N__56901\
        );

    \I__14116\ : InMux
    port map (
            O => \N__57099\,
            I => \N__56901\
        );

    \I__14115\ : InMux
    port map (
            O => \N__57098\,
            I => \N__56901\
        );

    \I__14114\ : InMux
    port map (
            O => \N__57097\,
            I => \N__56895\
        );

    \I__14113\ : LocalMux
    port map (
            O => \N__57094\,
            I => \N__56892\
        );

    \I__14112\ : InMux
    port map (
            O => \N__57093\,
            I => \N__56889\
        );

    \I__14111\ : InMux
    port map (
            O => \N__57092\,
            I => \N__56884\
        );

    \I__14110\ : InMux
    port map (
            O => \N__57091\,
            I => \N__56884\
        );

    \I__14109\ : LocalMux
    port map (
            O => \N__57088\,
            I => \N__56881\
        );

    \I__14108\ : LocalMux
    port map (
            O => \N__57083\,
            I => \N__56878\
        );

    \I__14107\ : InMux
    port map (
            O => \N__57080\,
            I => \N__56875\
        );

    \I__14106\ : LocalMux
    port map (
            O => \N__57077\,
            I => \N__56870\
        );

    \I__14105\ : LocalMux
    port map (
            O => \N__57072\,
            I => \N__56856\
        );

    \I__14104\ : LocalMux
    port map (
            O => \N__57067\,
            I => \N__56856\
        );

    \I__14103\ : LocalMux
    port map (
            O => \N__57062\,
            I => \N__56856\
        );

    \I__14102\ : LocalMux
    port map (
            O => \N__57059\,
            I => \N__56856\
        );

    \I__14101\ : LocalMux
    port map (
            O => \N__57052\,
            I => \N__56853\
        );

    \I__14100\ : LocalMux
    port map (
            O => \N__57049\,
            I => \N__56848\
        );

    \I__14099\ : LocalMux
    port map (
            O => \N__57046\,
            I => \N__56848\
        );

    \I__14098\ : Span4Mux_h
    port map (
            O => \N__57043\,
            I => \N__56843\
        );

    \I__14097\ : LocalMux
    port map (
            O => \N__57038\,
            I => \N__56843\
        );

    \I__14096\ : LocalMux
    port map (
            O => \N__57035\,
            I => \N__56836\
        );

    \I__14095\ : LocalMux
    port map (
            O => \N__57032\,
            I => \N__56836\
        );

    \I__14094\ : LocalMux
    port map (
            O => \N__57029\,
            I => \N__56836\
        );

    \I__14093\ : InMux
    port map (
            O => \N__57028\,
            I => \N__56827\
        );

    \I__14092\ : InMux
    port map (
            O => \N__57027\,
            I => \N__56827\
        );

    \I__14091\ : InMux
    port map (
            O => \N__57026\,
            I => \N__56827\
        );

    \I__14090\ : InMux
    port map (
            O => \N__57025\,
            I => \N__56827\
        );

    \I__14089\ : InMux
    port map (
            O => \N__57024\,
            I => \N__56822\
        );

    \I__14088\ : InMux
    port map (
            O => \N__57023\,
            I => \N__56822\
        );

    \I__14087\ : LocalMux
    port map (
            O => \N__57018\,
            I => \N__56807\
        );

    \I__14086\ : LocalMux
    port map (
            O => \N__57015\,
            I => \N__56807\
        );

    \I__14085\ : Span4Mux_v
    port map (
            O => \N__57012\,
            I => \N__56807\
        );

    \I__14084\ : Span4Mux_v
    port map (
            O => \N__57007\,
            I => \N__56807\
        );

    \I__14083\ : LocalMux
    port map (
            O => \N__57004\,
            I => \N__56807\
        );

    \I__14082\ : LocalMux
    port map (
            O => \N__56999\,
            I => \N__56807\
        );

    \I__14081\ : Span4Mux_v
    port map (
            O => \N__56996\,
            I => \N__56807\
        );

    \I__14080\ : LocalMux
    port map (
            O => \N__56993\,
            I => \N__56802\
        );

    \I__14079\ : LocalMux
    port map (
            O => \N__56986\,
            I => \N__56802\
        );

    \I__14078\ : LocalMux
    port map (
            O => \N__56983\,
            I => \N__56791\
        );

    \I__14077\ : LocalMux
    port map (
            O => \N__56980\,
            I => \N__56791\
        );

    \I__14076\ : Span4Mux_v
    port map (
            O => \N__56975\,
            I => \N__56791\
        );

    \I__14075\ : Span4Mux_h
    port map (
            O => \N__56972\,
            I => \N__56791\
        );

    \I__14074\ : LocalMux
    port map (
            O => \N__56961\,
            I => \N__56791\
        );

    \I__14073\ : CascadeMux
    port map (
            O => \N__56960\,
            I => \N__56788\
        );

    \I__14072\ : CascadeMux
    port map (
            O => \N__56959\,
            I => \N__56784\
        );

    \I__14071\ : InMux
    port map (
            O => \N__56958\,
            I => \N__56778\
        );

    \I__14070\ : InMux
    port map (
            O => \N__56957\,
            I => \N__56778\
        );

    \I__14069\ : LocalMux
    port map (
            O => \N__56954\,
            I => \N__56767\
        );

    \I__14068\ : LocalMux
    port map (
            O => \N__56949\,
            I => \N__56767\
        );

    \I__14067\ : LocalMux
    port map (
            O => \N__56946\,
            I => \N__56767\
        );

    \I__14066\ : LocalMux
    port map (
            O => \N__56943\,
            I => \N__56767\
        );

    \I__14065\ : Sp12to4
    port map (
            O => \N__56938\,
            I => \N__56767\
        );

    \I__14064\ : InMux
    port map (
            O => \N__56937\,
            I => \N__56764\
        );

    \I__14063\ : LocalMux
    port map (
            O => \N__56934\,
            I => \N__56753\
        );

    \I__14062\ : LocalMux
    port map (
            O => \N__56931\,
            I => \N__56753\
        );

    \I__14061\ : LocalMux
    port map (
            O => \N__56928\,
            I => \N__56753\
        );

    \I__14060\ : LocalMux
    port map (
            O => \N__56925\,
            I => \N__56753\
        );

    \I__14059\ : LocalMux
    port map (
            O => \N__56918\,
            I => \N__56753\
        );

    \I__14058\ : LocalMux
    port map (
            O => \N__56915\,
            I => \N__56748\
        );

    \I__14057\ : InMux
    port map (
            O => \N__56914\,
            I => \N__56743\
        );

    \I__14056\ : InMux
    port map (
            O => \N__56913\,
            I => \N__56743\
        );

    \I__14055\ : Span4Mux_v
    port map (
            O => \N__56910\,
            I => \N__56738\
        );

    \I__14054\ : LocalMux
    port map (
            O => \N__56901\,
            I => \N__56738\
        );

    \I__14053\ : InMux
    port map (
            O => \N__56900\,
            I => \N__56731\
        );

    \I__14052\ : InMux
    port map (
            O => \N__56899\,
            I => \N__56731\
        );

    \I__14051\ : InMux
    port map (
            O => \N__56898\,
            I => \N__56731\
        );

    \I__14050\ : LocalMux
    port map (
            O => \N__56895\,
            I => \N__56728\
        );

    \I__14049\ : Span4Mux_v
    port map (
            O => \N__56892\,
            I => \N__56723\
        );

    \I__14048\ : LocalMux
    port map (
            O => \N__56889\,
            I => \N__56723\
        );

    \I__14047\ : LocalMux
    port map (
            O => \N__56884\,
            I => \N__56720\
        );

    \I__14046\ : Span4Mux_v
    port map (
            O => \N__56881\,
            I => \N__56713\
        );

    \I__14045\ : Span4Mux_h
    port map (
            O => \N__56878\,
            I => \N__56713\
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__56875\,
            I => \N__56713\
        );

    \I__14043\ : InMux
    port map (
            O => \N__56874\,
            I => \N__56710\
        );

    \I__14042\ : InMux
    port map (
            O => \N__56873\,
            I => \N__56707\
        );

    \I__14041\ : Span4Mux_v
    port map (
            O => \N__56870\,
            I => \N__56704\
        );

    \I__14040\ : InMux
    port map (
            O => \N__56869\,
            I => \N__56697\
        );

    \I__14039\ : InMux
    port map (
            O => \N__56868\,
            I => \N__56697\
        );

    \I__14038\ : InMux
    port map (
            O => \N__56867\,
            I => \N__56697\
        );

    \I__14037\ : InMux
    port map (
            O => \N__56866\,
            I => \N__56692\
        );

    \I__14036\ : InMux
    port map (
            O => \N__56865\,
            I => \N__56692\
        );

    \I__14035\ : Span4Mux_v
    port map (
            O => \N__56856\,
            I => \N__56687\
        );

    \I__14034\ : Span4Mux_v
    port map (
            O => \N__56853\,
            I => \N__56687\
        );

    \I__14033\ : Span4Mux_h
    port map (
            O => \N__56848\,
            I => \N__56680\
        );

    \I__14032\ : Span4Mux_h
    port map (
            O => \N__56843\,
            I => \N__56680\
        );

    \I__14031\ : Span4Mux_h
    port map (
            O => \N__56836\,
            I => \N__56680\
        );

    \I__14030\ : LocalMux
    port map (
            O => \N__56827\,
            I => \N__56669\
        );

    \I__14029\ : LocalMux
    port map (
            O => \N__56822\,
            I => \N__56669\
        );

    \I__14028\ : Span4Mux_h
    port map (
            O => \N__56807\,
            I => \N__56669\
        );

    \I__14027\ : Span4Mux_h
    port map (
            O => \N__56802\,
            I => \N__56669\
        );

    \I__14026\ : Span4Mux_v
    port map (
            O => \N__56791\,
            I => \N__56669\
        );

    \I__14025\ : InMux
    port map (
            O => \N__56788\,
            I => \N__56660\
        );

    \I__14024\ : InMux
    port map (
            O => \N__56787\,
            I => \N__56660\
        );

    \I__14023\ : InMux
    port map (
            O => \N__56784\,
            I => \N__56660\
        );

    \I__14022\ : InMux
    port map (
            O => \N__56783\,
            I => \N__56660\
        );

    \I__14021\ : LocalMux
    port map (
            O => \N__56778\,
            I => \N__56655\
        );

    \I__14020\ : Span12Mux_h
    port map (
            O => \N__56767\,
            I => \N__56655\
        );

    \I__14019\ : LocalMux
    port map (
            O => \N__56764\,
            I => \N__56650\
        );

    \I__14018\ : Span12Mux_v
    port map (
            O => \N__56753\,
            I => \N__56650\
        );

    \I__14017\ : InMux
    port map (
            O => \N__56752\,
            I => \N__56645\
        );

    \I__14016\ : InMux
    port map (
            O => \N__56751\,
            I => \N__56645\
        );

    \I__14015\ : Span4Mux_v
    port map (
            O => \N__56748\,
            I => \N__56628\
        );

    \I__14014\ : LocalMux
    port map (
            O => \N__56743\,
            I => \N__56628\
        );

    \I__14013\ : Span4Mux_h
    port map (
            O => \N__56738\,
            I => \N__56628\
        );

    \I__14012\ : LocalMux
    port map (
            O => \N__56731\,
            I => \N__56628\
        );

    \I__14011\ : Span4Mux_v
    port map (
            O => \N__56728\,
            I => \N__56628\
        );

    \I__14010\ : Span4Mux_h
    port map (
            O => \N__56723\,
            I => \N__56628\
        );

    \I__14009\ : Span4Mux_h
    port map (
            O => \N__56720\,
            I => \N__56628\
        );

    \I__14008\ : Span4Mux_h
    port map (
            O => \N__56713\,
            I => \N__56628\
        );

    \I__14007\ : LocalMux
    port map (
            O => \N__56710\,
            I => comm_cmd_0
        );

    \I__14006\ : LocalMux
    port map (
            O => \N__56707\,
            I => comm_cmd_0
        );

    \I__14005\ : Odrv4
    port map (
            O => \N__56704\,
            I => comm_cmd_0
        );

    \I__14004\ : LocalMux
    port map (
            O => \N__56697\,
            I => comm_cmd_0
        );

    \I__14003\ : LocalMux
    port map (
            O => \N__56692\,
            I => comm_cmd_0
        );

    \I__14002\ : Odrv4
    port map (
            O => \N__56687\,
            I => comm_cmd_0
        );

    \I__14001\ : Odrv4
    port map (
            O => \N__56680\,
            I => comm_cmd_0
        );

    \I__14000\ : Odrv4
    port map (
            O => \N__56669\,
            I => comm_cmd_0
        );

    \I__13999\ : LocalMux
    port map (
            O => \N__56660\,
            I => comm_cmd_0
        );

    \I__13998\ : Odrv12
    port map (
            O => \N__56655\,
            I => comm_cmd_0
        );

    \I__13997\ : Odrv12
    port map (
            O => \N__56650\,
            I => comm_cmd_0
        );

    \I__13996\ : LocalMux
    port map (
            O => \N__56645\,
            I => comm_cmd_0
        );

    \I__13995\ : Odrv4
    port map (
            O => \N__56628\,
            I => comm_cmd_0
        );

    \I__13994\ : InMux
    port map (
            O => \N__56601\,
            I => \N__56598\
        );

    \I__13993\ : LocalMux
    port map (
            O => \N__56598\,
            I => \N__56595\
        );

    \I__13992\ : Span4Mux_v
    port map (
            O => \N__56595\,
            I => \N__56592\
        );

    \I__13991\ : Span4Mux_h
    port map (
            O => \N__56592\,
            I => \N__56589\
        );

    \I__13990\ : Odrv4
    port map (
            O => \N__56589\,
            I => n21434
        );

    \I__13989\ : InMux
    port map (
            O => \N__56586\,
            I => \N__56583\
        );

    \I__13988\ : LocalMux
    port map (
            O => \N__56583\,
            I => \N__56579\
        );

    \I__13987\ : InMux
    port map (
            O => \N__56582\,
            I => \N__56575\
        );

    \I__13986\ : Span12Mux_s11_v
    port map (
            O => \N__56579\,
            I => \N__56568\
        );

    \I__13985\ : InMux
    port map (
            O => \N__56578\,
            I => \N__56565\
        );

    \I__13984\ : LocalMux
    port map (
            O => \N__56575\,
            I => \N__56562\
        );

    \I__13983\ : InMux
    port map (
            O => \N__56574\,
            I => \N__56557\
        );

    \I__13982\ : InMux
    port map (
            O => \N__56573\,
            I => \N__56557\
        );

    \I__13981\ : InMux
    port map (
            O => \N__56572\,
            I => \N__56552\
        );

    \I__13980\ : InMux
    port map (
            O => \N__56571\,
            I => \N__56552\
        );

    \I__13979\ : Odrv12
    port map (
            O => \N__56568\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__13978\ : LocalMux
    port map (
            O => \N__56565\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__13977\ : Odrv4
    port map (
            O => \N__56562\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__13976\ : LocalMux
    port map (
            O => \N__56557\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__13975\ : LocalMux
    port map (
            O => \N__56552\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__13974\ : CascadeMux
    port map (
            O => \N__56541\,
            I => \N__56538\
        );

    \I__13973\ : InMux
    port map (
            O => \N__56538\,
            I => \N__56534\
        );

    \I__13972\ : InMux
    port map (
            O => \N__56537\,
            I => \N__56531\
        );

    \I__13971\ : LocalMux
    port map (
            O => \N__56534\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__13970\ : LocalMux
    port map (
            O => \N__56531\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__13969\ : InMux
    port map (
            O => \N__56526\,
            I => \N__56523\
        );

    \I__13968\ : LocalMux
    port map (
            O => \N__56523\,
            I => \N__56520\
        );

    \I__13967\ : Odrv4
    port map (
            O => \N__56520\,
            I => \ADC_VDC.genclk.n28\
        );

    \I__13966\ : InMux
    port map (
            O => \N__56517\,
            I => \N__56514\
        );

    \I__13965\ : LocalMux
    port map (
            O => \N__56514\,
            I => \ADC_VDC.genclk.n26_adj_1448\
        );

    \I__13964\ : InMux
    port map (
            O => \N__56511\,
            I => \N__56508\
        );

    \I__13963\ : LocalMux
    port map (
            O => \N__56508\,
            I => \N__56505\
        );

    \I__13962\ : Span4Mux_v
    port map (
            O => \N__56505\,
            I => \N__56500\
        );

    \I__13961\ : InMux
    port map (
            O => \N__56504\,
            I => \N__56497\
        );

    \I__13960\ : InMux
    port map (
            O => \N__56503\,
            I => \N__56494\
        );

    \I__13959\ : Odrv4
    port map (
            O => \N__56500\,
            I => \comm_spi.n23101\
        );

    \I__13958\ : LocalMux
    port map (
            O => \N__56497\,
            I => \comm_spi.n23101\
        );

    \I__13957\ : LocalMux
    port map (
            O => \N__56494\,
            I => \comm_spi.n23101\
        );

    \I__13956\ : InMux
    port map (
            O => \N__56487\,
            I => \N__56483\
        );

    \I__13955\ : InMux
    port map (
            O => \N__56486\,
            I => \N__56480\
        );

    \I__13954\ : LocalMux
    port map (
            O => \N__56483\,
            I => \N__56477\
        );

    \I__13953\ : LocalMux
    port map (
            O => \N__56480\,
            I => \N__56474\
        );

    \I__13952\ : Span4Mux_h
    port map (
            O => \N__56477\,
            I => \N__56469\
        );

    \I__13951\ : Span4Mux_v
    port map (
            O => \N__56474\,
            I => \N__56469\
        );

    \I__13950\ : Odrv4
    port map (
            O => \N__56469\,
            I => \comm_spi.n14834\
        );

    \I__13949\ : SRMux
    port map (
            O => \N__56466\,
            I => \N__56463\
        );

    \I__13948\ : LocalMux
    port map (
            O => \N__56463\,
            I => \N__56460\
        );

    \I__13947\ : Odrv12
    port map (
            O => \N__56460\,
            I => \comm_spi.data_tx_7__N_823\
        );

    \I__13946\ : SRMux
    port map (
            O => \N__56457\,
            I => \N__56454\
        );

    \I__13945\ : LocalMux
    port map (
            O => \N__56454\,
            I => \N__56451\
        );

    \I__13944\ : Odrv12
    port map (
            O => \N__56451\,
            I => \comm_spi.data_tx_7__N_811\
        );

    \I__13943\ : InMux
    port map (
            O => \N__56448\,
            I => \N__56443\
        );

    \I__13942\ : InMux
    port map (
            O => \N__56447\,
            I => \N__56438\
        );

    \I__13941\ : InMux
    port map (
            O => \N__56446\,
            I => \N__56438\
        );

    \I__13940\ : LocalMux
    port map (
            O => \N__56443\,
            I => \N__56435\
        );

    \I__13939\ : LocalMux
    port map (
            O => \N__56438\,
            I => \N__56432\
        );

    \I__13938\ : Span4Mux_h
    port map (
            O => \N__56435\,
            I => \N__56429\
        );

    \I__13937\ : Span4Mux_h
    port map (
            O => \N__56432\,
            I => \N__56426\
        );

    \I__13936\ : Odrv4
    port map (
            O => \N__56429\,
            I => comm_tx_buf_4
        );

    \I__13935\ : Odrv4
    port map (
            O => \N__56426\,
            I => comm_tx_buf_4
        );

    \I__13934\ : SRMux
    port map (
            O => \N__56421\,
            I => \N__56418\
        );

    \I__13933\ : LocalMux
    port map (
            O => \N__56418\,
            I => \N__56415\
        );

    \I__13932\ : Span4Mux_v
    port map (
            O => \N__56415\,
            I => \N__56412\
        );

    \I__13931\ : Span4Mux_h
    port map (
            O => \N__56412\,
            I => \N__56409\
        );

    \I__13930\ : Span4Mux_h
    port map (
            O => \N__56409\,
            I => \N__56406\
        );

    \I__13929\ : Odrv4
    port map (
            O => \N__56406\,
            I => \comm_spi.data_tx_7__N_809\
        );

    \I__13928\ : InMux
    port map (
            O => \N__56403\,
            I => \N__56394\
        );

    \I__13927\ : InMux
    port map (
            O => \N__56402\,
            I => \N__56394\
        );

    \I__13926\ : InMux
    port map (
            O => \N__56401\,
            I => \N__56394\
        );

    \I__13925\ : LocalMux
    port map (
            O => \N__56394\,
            I => \N__56391\
        );

    \I__13924\ : Span4Mux_v
    port map (
            O => \N__56391\,
            I => \N__56388\
        );

    \I__13923\ : Odrv4
    port map (
            O => \N__56388\,
            I => comm_tx_buf_2
        );

    \I__13922\ : CascadeMux
    port map (
            O => \N__56385\,
            I => \N__56382\
        );

    \I__13921\ : InMux
    port map (
            O => \N__56382\,
            I => \N__56378\
        );

    \I__13920\ : InMux
    port map (
            O => \N__56381\,
            I => \N__56375\
        );

    \I__13919\ : LocalMux
    port map (
            O => \N__56378\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__13918\ : LocalMux
    port map (
            O => \N__56375\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__13917\ : InMux
    port map (
            O => \N__56370\,
            I => \N__56366\
        );

    \I__13916\ : InMux
    port map (
            O => \N__56369\,
            I => \N__56363\
        );

    \I__13915\ : LocalMux
    port map (
            O => \N__56366\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__13914\ : LocalMux
    port map (
            O => \N__56363\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__13913\ : CascadeMux
    port map (
            O => \N__56358\,
            I => \N__56354\
        );

    \I__13912\ : CascadeMux
    port map (
            O => \N__56357\,
            I => \N__56351\
        );

    \I__13911\ : InMux
    port map (
            O => \N__56354\,
            I => \N__56348\
        );

    \I__13910\ : InMux
    port map (
            O => \N__56351\,
            I => \N__56345\
        );

    \I__13909\ : LocalMux
    port map (
            O => \N__56348\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__13908\ : LocalMux
    port map (
            O => \N__56345\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__13907\ : InMux
    port map (
            O => \N__56340\,
            I => \N__56336\
        );

    \I__13906\ : InMux
    port map (
            O => \N__56339\,
            I => \N__56333\
        );

    \I__13905\ : LocalMux
    port map (
            O => \N__56336\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__13904\ : LocalMux
    port map (
            O => \N__56333\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__13903\ : InMux
    port map (
            O => \N__56328\,
            I => \N__56325\
        );

    \I__13902\ : LocalMux
    port map (
            O => \N__56325\,
            I => \ADC_VDC.genclk.n21600\
        );

    \I__13901\ : CascadeMux
    port map (
            O => \N__56322\,
            I => \ADC_VDC.genclk.n27_adj_1449_cascade_\
        );

    \I__13900\ : InMux
    port map (
            O => \N__56319\,
            I => \N__56316\
        );

    \I__13899\ : LocalMux
    port map (
            O => \N__56316\,
            I => \ADC_VDC.genclk.n21597\
        );

    \I__13898\ : InMux
    port map (
            O => \N__56313\,
            I => \N__56310\
        );

    \I__13897\ : LocalMux
    port map (
            O => \N__56310\,
            I => \ADC_VDC.genclk.n21598\
        );

    \I__13896\ : CascadeMux
    port map (
            O => \N__56307\,
            I => \ADC_VDC.genclk.n21597_cascade_\
        );

    \I__13895\ : InMux
    port map (
            O => \N__56304\,
            I => \N__56301\
        );

    \I__13894\ : LocalMux
    port map (
            O => \N__56301\,
            I => \ADC_VDC.genclk.n21603\
        );

    \I__13893\ : CascadeMux
    port map (
            O => \N__56298\,
            I => \N__56294\
        );

    \I__13892\ : InMux
    port map (
            O => \N__56297\,
            I => \N__56291\
        );

    \I__13891\ : InMux
    port map (
            O => \N__56294\,
            I => \N__56288\
        );

    \I__13890\ : LocalMux
    port map (
            O => \N__56291\,
            I => \N__56285\
        );

    \I__13889\ : LocalMux
    port map (
            O => \N__56288\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__13888\ : Odrv4
    port map (
            O => \N__56285\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__13887\ : InMux
    port map (
            O => \N__56280\,
            I => \N__56276\
        );

    \I__13886\ : InMux
    port map (
            O => \N__56279\,
            I => \N__56273\
        );

    \I__13885\ : LocalMux
    port map (
            O => \N__56276\,
            I => \N__56270\
        );

    \I__13884\ : LocalMux
    port map (
            O => \N__56273\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__13883\ : Odrv4
    port map (
            O => \N__56270\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__13882\ : CascadeMux
    port map (
            O => \N__56265\,
            I => \N__56261\
        );

    \I__13881\ : InMux
    port map (
            O => \N__56264\,
            I => \N__56258\
        );

    \I__13880\ : InMux
    port map (
            O => \N__56261\,
            I => \N__56255\
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__56258\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__13878\ : LocalMux
    port map (
            O => \N__56255\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__13877\ : InMux
    port map (
            O => \N__56250\,
            I => \N__56246\
        );

    \I__13876\ : InMux
    port map (
            O => \N__56249\,
            I => \N__56243\
        );

    \I__13875\ : LocalMux
    port map (
            O => \N__56246\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__13874\ : LocalMux
    port map (
            O => \N__56243\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__13873\ : InMux
    port map (
            O => \N__56238\,
            I => \N__56235\
        );

    \I__13872\ : LocalMux
    port map (
            O => \N__56235\,
            I => \ADC_VDC.genclk.n26\
        );

    \I__13871\ : InMux
    port map (
            O => \N__56232\,
            I => \N__56225\
        );

    \I__13870\ : InMux
    port map (
            O => \N__56231\,
            I => \N__56222\
        );

    \I__13869\ : InMux
    port map (
            O => \N__56230\,
            I => \N__56217\
        );

    \I__13868\ : InMux
    port map (
            O => \N__56229\,
            I => \N__56217\
        );

    \I__13867\ : InMux
    port map (
            O => \N__56228\,
            I => \N__56214\
        );

    \I__13866\ : LocalMux
    port map (
            O => \N__56225\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__13865\ : LocalMux
    port map (
            O => \N__56222\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__13864\ : LocalMux
    port map (
            O => \N__56217\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__13863\ : LocalMux
    port map (
            O => \N__56214\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__13862\ : InMux
    port map (
            O => \N__56205\,
            I => \N__56202\
        );

    \I__13861\ : LocalMux
    port map (
            O => \N__56202\,
            I => \ADC_VDC.genclk.n28_adj_1447\
        );

    \I__13860\ : InMux
    port map (
            O => \N__56199\,
            I => \N__56195\
        );

    \I__13859\ : InMux
    port map (
            O => \N__56198\,
            I => \N__56192\
        );

    \I__13858\ : LocalMux
    port map (
            O => \N__56195\,
            I => \N__56187\
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__56192\,
            I => \N__56187\
        );

    \I__13856\ : Odrv4
    port map (
            O => \N__56187\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__13855\ : CascadeMux
    port map (
            O => \N__56184\,
            I => \N__56181\
        );

    \I__13854\ : InMux
    port map (
            O => \N__56181\,
            I => \N__56177\
        );

    \I__13853\ : InMux
    port map (
            O => \N__56180\,
            I => \N__56174\
        );

    \I__13852\ : LocalMux
    port map (
            O => \N__56177\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__13851\ : LocalMux
    port map (
            O => \N__56174\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__13850\ : CascadeMux
    port map (
            O => \N__56169\,
            I => \N__56165\
        );

    \I__13849\ : InMux
    port map (
            O => \N__56168\,
            I => \N__56162\
        );

    \I__13848\ : InMux
    port map (
            O => \N__56165\,
            I => \N__56159\
        );

    \I__13847\ : LocalMux
    port map (
            O => \N__56162\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__13846\ : LocalMux
    port map (
            O => \N__56159\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__13845\ : InMux
    port map (
            O => \N__56154\,
            I => \N__56151\
        );

    \I__13844\ : LocalMux
    port map (
            O => \N__56151\,
            I => \N__56148\
        );

    \I__13843\ : Span4Mux_v
    port map (
            O => \N__56148\,
            I => \N__56144\
        );

    \I__13842\ : InMux
    port map (
            O => \N__56147\,
            I => \N__56141\
        );

    \I__13841\ : Span4Mux_v
    port map (
            O => \N__56144\,
            I => \N__56135\
        );

    \I__13840\ : LocalMux
    port map (
            O => \N__56141\,
            I => \N__56135\
        );

    \I__13839\ : InMux
    port map (
            O => \N__56140\,
            I => \N__56132\
        );

    \I__13838\ : Span4Mux_v
    port map (
            O => \N__56135\,
            I => \N__56129\
        );

    \I__13837\ : LocalMux
    port map (
            O => \N__56132\,
            I => \N__56126\
        );

    \I__13836\ : Sp12to4
    port map (
            O => \N__56129\,
            I => \N__56121\
        );

    \I__13835\ : Span12Mux_v
    port map (
            O => \N__56126\,
            I => \N__56121\
        );

    \I__13834\ : Odrv12
    port map (
            O => \N__56121\,
            I => comm_tx_buf_3
        );

    \I__13833\ : IoInMux
    port map (
            O => \N__56118\,
            I => \N__56115\
        );

    \I__13832\ : LocalMux
    port map (
            O => \N__56115\,
            I => \N__56112\
        );

    \I__13831\ : Span12Mux_s9_h
    port map (
            O => \N__56112\,
            I => \N__56109\
        );

    \I__13830\ : Span12Mux_v
    port map (
            O => \N__56109\,
            I => \N__56106\
        );

    \I__13829\ : Odrv12
    port map (
            O => \N__56106\,
            I => \ICE_GPMI_0\
        );

    \I__13828\ : ClkMux
    port map (
            O => \N__56103\,
            I => \N__55602\
        );

    \I__13827\ : ClkMux
    port map (
            O => \N__56102\,
            I => \N__55602\
        );

    \I__13826\ : ClkMux
    port map (
            O => \N__56101\,
            I => \N__55602\
        );

    \I__13825\ : ClkMux
    port map (
            O => \N__56100\,
            I => \N__55602\
        );

    \I__13824\ : ClkMux
    port map (
            O => \N__56099\,
            I => \N__55602\
        );

    \I__13823\ : ClkMux
    port map (
            O => \N__56098\,
            I => \N__55602\
        );

    \I__13822\ : ClkMux
    port map (
            O => \N__56097\,
            I => \N__55602\
        );

    \I__13821\ : ClkMux
    port map (
            O => \N__56096\,
            I => \N__55602\
        );

    \I__13820\ : ClkMux
    port map (
            O => \N__56095\,
            I => \N__55602\
        );

    \I__13819\ : ClkMux
    port map (
            O => \N__56094\,
            I => \N__55602\
        );

    \I__13818\ : ClkMux
    port map (
            O => \N__56093\,
            I => \N__55602\
        );

    \I__13817\ : ClkMux
    port map (
            O => \N__56092\,
            I => \N__55602\
        );

    \I__13816\ : ClkMux
    port map (
            O => \N__56091\,
            I => \N__55602\
        );

    \I__13815\ : ClkMux
    port map (
            O => \N__56090\,
            I => \N__55602\
        );

    \I__13814\ : ClkMux
    port map (
            O => \N__56089\,
            I => \N__55602\
        );

    \I__13813\ : ClkMux
    port map (
            O => \N__56088\,
            I => \N__55602\
        );

    \I__13812\ : ClkMux
    port map (
            O => \N__56087\,
            I => \N__55602\
        );

    \I__13811\ : ClkMux
    port map (
            O => \N__56086\,
            I => \N__55602\
        );

    \I__13810\ : ClkMux
    port map (
            O => \N__56085\,
            I => \N__55602\
        );

    \I__13809\ : ClkMux
    port map (
            O => \N__56084\,
            I => \N__55602\
        );

    \I__13808\ : ClkMux
    port map (
            O => \N__56083\,
            I => \N__55602\
        );

    \I__13807\ : ClkMux
    port map (
            O => \N__56082\,
            I => \N__55602\
        );

    \I__13806\ : ClkMux
    port map (
            O => \N__56081\,
            I => \N__55602\
        );

    \I__13805\ : ClkMux
    port map (
            O => \N__56080\,
            I => \N__55602\
        );

    \I__13804\ : ClkMux
    port map (
            O => \N__56079\,
            I => \N__55602\
        );

    \I__13803\ : ClkMux
    port map (
            O => \N__56078\,
            I => \N__55602\
        );

    \I__13802\ : ClkMux
    port map (
            O => \N__56077\,
            I => \N__55602\
        );

    \I__13801\ : ClkMux
    port map (
            O => \N__56076\,
            I => \N__55602\
        );

    \I__13800\ : ClkMux
    port map (
            O => \N__56075\,
            I => \N__55602\
        );

    \I__13799\ : ClkMux
    port map (
            O => \N__56074\,
            I => \N__55602\
        );

    \I__13798\ : ClkMux
    port map (
            O => \N__56073\,
            I => \N__55602\
        );

    \I__13797\ : ClkMux
    port map (
            O => \N__56072\,
            I => \N__55602\
        );

    \I__13796\ : ClkMux
    port map (
            O => \N__56071\,
            I => \N__55602\
        );

    \I__13795\ : ClkMux
    port map (
            O => \N__56070\,
            I => \N__55602\
        );

    \I__13794\ : ClkMux
    port map (
            O => \N__56069\,
            I => \N__55602\
        );

    \I__13793\ : ClkMux
    port map (
            O => \N__56068\,
            I => \N__55602\
        );

    \I__13792\ : ClkMux
    port map (
            O => \N__56067\,
            I => \N__55602\
        );

    \I__13791\ : ClkMux
    port map (
            O => \N__56066\,
            I => \N__55602\
        );

    \I__13790\ : ClkMux
    port map (
            O => \N__56065\,
            I => \N__55602\
        );

    \I__13789\ : ClkMux
    port map (
            O => \N__56064\,
            I => \N__55602\
        );

    \I__13788\ : ClkMux
    port map (
            O => \N__56063\,
            I => \N__55602\
        );

    \I__13787\ : ClkMux
    port map (
            O => \N__56062\,
            I => \N__55602\
        );

    \I__13786\ : ClkMux
    port map (
            O => \N__56061\,
            I => \N__55602\
        );

    \I__13785\ : ClkMux
    port map (
            O => \N__56060\,
            I => \N__55602\
        );

    \I__13784\ : ClkMux
    port map (
            O => \N__56059\,
            I => \N__55602\
        );

    \I__13783\ : ClkMux
    port map (
            O => \N__56058\,
            I => \N__55602\
        );

    \I__13782\ : ClkMux
    port map (
            O => \N__56057\,
            I => \N__55602\
        );

    \I__13781\ : ClkMux
    port map (
            O => \N__56056\,
            I => \N__55602\
        );

    \I__13780\ : ClkMux
    port map (
            O => \N__56055\,
            I => \N__55602\
        );

    \I__13779\ : ClkMux
    port map (
            O => \N__56054\,
            I => \N__55602\
        );

    \I__13778\ : ClkMux
    port map (
            O => \N__56053\,
            I => \N__55602\
        );

    \I__13777\ : ClkMux
    port map (
            O => \N__56052\,
            I => \N__55602\
        );

    \I__13776\ : ClkMux
    port map (
            O => \N__56051\,
            I => \N__55602\
        );

    \I__13775\ : ClkMux
    port map (
            O => \N__56050\,
            I => \N__55602\
        );

    \I__13774\ : ClkMux
    port map (
            O => \N__56049\,
            I => \N__55602\
        );

    \I__13773\ : ClkMux
    port map (
            O => \N__56048\,
            I => \N__55602\
        );

    \I__13772\ : ClkMux
    port map (
            O => \N__56047\,
            I => \N__55602\
        );

    \I__13771\ : ClkMux
    port map (
            O => \N__56046\,
            I => \N__55602\
        );

    \I__13770\ : ClkMux
    port map (
            O => \N__56045\,
            I => \N__55602\
        );

    \I__13769\ : ClkMux
    port map (
            O => \N__56044\,
            I => \N__55602\
        );

    \I__13768\ : ClkMux
    port map (
            O => \N__56043\,
            I => \N__55602\
        );

    \I__13767\ : ClkMux
    port map (
            O => \N__56042\,
            I => \N__55602\
        );

    \I__13766\ : ClkMux
    port map (
            O => \N__56041\,
            I => \N__55602\
        );

    \I__13765\ : ClkMux
    port map (
            O => \N__56040\,
            I => \N__55602\
        );

    \I__13764\ : ClkMux
    port map (
            O => \N__56039\,
            I => \N__55602\
        );

    \I__13763\ : ClkMux
    port map (
            O => \N__56038\,
            I => \N__55602\
        );

    \I__13762\ : ClkMux
    port map (
            O => \N__56037\,
            I => \N__55602\
        );

    \I__13761\ : ClkMux
    port map (
            O => \N__56036\,
            I => \N__55602\
        );

    \I__13760\ : ClkMux
    port map (
            O => \N__56035\,
            I => \N__55602\
        );

    \I__13759\ : ClkMux
    port map (
            O => \N__56034\,
            I => \N__55602\
        );

    \I__13758\ : ClkMux
    port map (
            O => \N__56033\,
            I => \N__55602\
        );

    \I__13757\ : ClkMux
    port map (
            O => \N__56032\,
            I => \N__55602\
        );

    \I__13756\ : ClkMux
    port map (
            O => \N__56031\,
            I => \N__55602\
        );

    \I__13755\ : ClkMux
    port map (
            O => \N__56030\,
            I => \N__55602\
        );

    \I__13754\ : ClkMux
    port map (
            O => \N__56029\,
            I => \N__55602\
        );

    \I__13753\ : ClkMux
    port map (
            O => \N__56028\,
            I => \N__55602\
        );

    \I__13752\ : ClkMux
    port map (
            O => \N__56027\,
            I => \N__55602\
        );

    \I__13751\ : ClkMux
    port map (
            O => \N__56026\,
            I => \N__55602\
        );

    \I__13750\ : ClkMux
    port map (
            O => \N__56025\,
            I => \N__55602\
        );

    \I__13749\ : ClkMux
    port map (
            O => \N__56024\,
            I => \N__55602\
        );

    \I__13748\ : ClkMux
    port map (
            O => \N__56023\,
            I => \N__55602\
        );

    \I__13747\ : ClkMux
    port map (
            O => \N__56022\,
            I => \N__55602\
        );

    \I__13746\ : ClkMux
    port map (
            O => \N__56021\,
            I => \N__55602\
        );

    \I__13745\ : ClkMux
    port map (
            O => \N__56020\,
            I => \N__55602\
        );

    \I__13744\ : ClkMux
    port map (
            O => \N__56019\,
            I => \N__55602\
        );

    \I__13743\ : ClkMux
    port map (
            O => \N__56018\,
            I => \N__55602\
        );

    \I__13742\ : ClkMux
    port map (
            O => \N__56017\,
            I => \N__55602\
        );

    \I__13741\ : ClkMux
    port map (
            O => \N__56016\,
            I => \N__55602\
        );

    \I__13740\ : ClkMux
    port map (
            O => \N__56015\,
            I => \N__55602\
        );

    \I__13739\ : ClkMux
    port map (
            O => \N__56014\,
            I => \N__55602\
        );

    \I__13738\ : ClkMux
    port map (
            O => \N__56013\,
            I => \N__55602\
        );

    \I__13737\ : ClkMux
    port map (
            O => \N__56012\,
            I => \N__55602\
        );

    \I__13736\ : ClkMux
    port map (
            O => \N__56011\,
            I => \N__55602\
        );

    \I__13735\ : ClkMux
    port map (
            O => \N__56010\,
            I => \N__55602\
        );

    \I__13734\ : ClkMux
    port map (
            O => \N__56009\,
            I => \N__55602\
        );

    \I__13733\ : ClkMux
    port map (
            O => \N__56008\,
            I => \N__55602\
        );

    \I__13732\ : ClkMux
    port map (
            O => \N__56007\,
            I => \N__55602\
        );

    \I__13731\ : ClkMux
    port map (
            O => \N__56006\,
            I => \N__55602\
        );

    \I__13730\ : ClkMux
    port map (
            O => \N__56005\,
            I => \N__55602\
        );

    \I__13729\ : ClkMux
    port map (
            O => \N__56004\,
            I => \N__55602\
        );

    \I__13728\ : ClkMux
    port map (
            O => \N__56003\,
            I => \N__55602\
        );

    \I__13727\ : ClkMux
    port map (
            O => \N__56002\,
            I => \N__55602\
        );

    \I__13726\ : ClkMux
    port map (
            O => \N__56001\,
            I => \N__55602\
        );

    \I__13725\ : ClkMux
    port map (
            O => \N__56000\,
            I => \N__55602\
        );

    \I__13724\ : ClkMux
    port map (
            O => \N__55999\,
            I => \N__55602\
        );

    \I__13723\ : ClkMux
    port map (
            O => \N__55998\,
            I => \N__55602\
        );

    \I__13722\ : ClkMux
    port map (
            O => \N__55997\,
            I => \N__55602\
        );

    \I__13721\ : ClkMux
    port map (
            O => \N__55996\,
            I => \N__55602\
        );

    \I__13720\ : ClkMux
    port map (
            O => \N__55995\,
            I => \N__55602\
        );

    \I__13719\ : ClkMux
    port map (
            O => \N__55994\,
            I => \N__55602\
        );

    \I__13718\ : ClkMux
    port map (
            O => \N__55993\,
            I => \N__55602\
        );

    \I__13717\ : ClkMux
    port map (
            O => \N__55992\,
            I => \N__55602\
        );

    \I__13716\ : ClkMux
    port map (
            O => \N__55991\,
            I => \N__55602\
        );

    \I__13715\ : ClkMux
    port map (
            O => \N__55990\,
            I => \N__55602\
        );

    \I__13714\ : ClkMux
    port map (
            O => \N__55989\,
            I => \N__55602\
        );

    \I__13713\ : ClkMux
    port map (
            O => \N__55988\,
            I => \N__55602\
        );

    \I__13712\ : ClkMux
    port map (
            O => \N__55987\,
            I => \N__55602\
        );

    \I__13711\ : ClkMux
    port map (
            O => \N__55986\,
            I => \N__55602\
        );

    \I__13710\ : ClkMux
    port map (
            O => \N__55985\,
            I => \N__55602\
        );

    \I__13709\ : ClkMux
    port map (
            O => \N__55984\,
            I => \N__55602\
        );

    \I__13708\ : ClkMux
    port map (
            O => \N__55983\,
            I => \N__55602\
        );

    \I__13707\ : ClkMux
    port map (
            O => \N__55982\,
            I => \N__55602\
        );

    \I__13706\ : ClkMux
    port map (
            O => \N__55981\,
            I => \N__55602\
        );

    \I__13705\ : ClkMux
    port map (
            O => \N__55980\,
            I => \N__55602\
        );

    \I__13704\ : ClkMux
    port map (
            O => \N__55979\,
            I => \N__55602\
        );

    \I__13703\ : ClkMux
    port map (
            O => \N__55978\,
            I => \N__55602\
        );

    \I__13702\ : ClkMux
    port map (
            O => \N__55977\,
            I => \N__55602\
        );

    \I__13701\ : ClkMux
    port map (
            O => \N__55976\,
            I => \N__55602\
        );

    \I__13700\ : ClkMux
    port map (
            O => \N__55975\,
            I => \N__55602\
        );

    \I__13699\ : ClkMux
    port map (
            O => \N__55974\,
            I => \N__55602\
        );

    \I__13698\ : ClkMux
    port map (
            O => \N__55973\,
            I => \N__55602\
        );

    \I__13697\ : ClkMux
    port map (
            O => \N__55972\,
            I => \N__55602\
        );

    \I__13696\ : ClkMux
    port map (
            O => \N__55971\,
            I => \N__55602\
        );

    \I__13695\ : ClkMux
    port map (
            O => \N__55970\,
            I => \N__55602\
        );

    \I__13694\ : ClkMux
    port map (
            O => \N__55969\,
            I => \N__55602\
        );

    \I__13693\ : ClkMux
    port map (
            O => \N__55968\,
            I => \N__55602\
        );

    \I__13692\ : ClkMux
    port map (
            O => \N__55967\,
            I => \N__55602\
        );

    \I__13691\ : ClkMux
    port map (
            O => \N__55966\,
            I => \N__55602\
        );

    \I__13690\ : ClkMux
    port map (
            O => \N__55965\,
            I => \N__55602\
        );

    \I__13689\ : ClkMux
    port map (
            O => \N__55964\,
            I => \N__55602\
        );

    \I__13688\ : ClkMux
    port map (
            O => \N__55963\,
            I => \N__55602\
        );

    \I__13687\ : ClkMux
    port map (
            O => \N__55962\,
            I => \N__55602\
        );

    \I__13686\ : ClkMux
    port map (
            O => \N__55961\,
            I => \N__55602\
        );

    \I__13685\ : ClkMux
    port map (
            O => \N__55960\,
            I => \N__55602\
        );

    \I__13684\ : ClkMux
    port map (
            O => \N__55959\,
            I => \N__55602\
        );

    \I__13683\ : ClkMux
    port map (
            O => \N__55958\,
            I => \N__55602\
        );

    \I__13682\ : ClkMux
    port map (
            O => \N__55957\,
            I => \N__55602\
        );

    \I__13681\ : ClkMux
    port map (
            O => \N__55956\,
            I => \N__55602\
        );

    \I__13680\ : ClkMux
    port map (
            O => \N__55955\,
            I => \N__55602\
        );

    \I__13679\ : ClkMux
    port map (
            O => \N__55954\,
            I => \N__55602\
        );

    \I__13678\ : ClkMux
    port map (
            O => \N__55953\,
            I => \N__55602\
        );

    \I__13677\ : ClkMux
    port map (
            O => \N__55952\,
            I => \N__55602\
        );

    \I__13676\ : ClkMux
    port map (
            O => \N__55951\,
            I => \N__55602\
        );

    \I__13675\ : ClkMux
    port map (
            O => \N__55950\,
            I => \N__55602\
        );

    \I__13674\ : ClkMux
    port map (
            O => \N__55949\,
            I => \N__55602\
        );

    \I__13673\ : ClkMux
    port map (
            O => \N__55948\,
            I => \N__55602\
        );

    \I__13672\ : ClkMux
    port map (
            O => \N__55947\,
            I => \N__55602\
        );

    \I__13671\ : ClkMux
    port map (
            O => \N__55946\,
            I => \N__55602\
        );

    \I__13670\ : ClkMux
    port map (
            O => \N__55945\,
            I => \N__55602\
        );

    \I__13669\ : ClkMux
    port map (
            O => \N__55944\,
            I => \N__55602\
        );

    \I__13668\ : ClkMux
    port map (
            O => \N__55943\,
            I => \N__55602\
        );

    \I__13667\ : ClkMux
    port map (
            O => \N__55942\,
            I => \N__55602\
        );

    \I__13666\ : ClkMux
    port map (
            O => \N__55941\,
            I => \N__55602\
        );

    \I__13665\ : ClkMux
    port map (
            O => \N__55940\,
            I => \N__55602\
        );

    \I__13664\ : ClkMux
    port map (
            O => \N__55939\,
            I => \N__55602\
        );

    \I__13663\ : ClkMux
    port map (
            O => \N__55938\,
            I => \N__55602\
        );

    \I__13662\ : ClkMux
    port map (
            O => \N__55937\,
            I => \N__55602\
        );

    \I__13661\ : GlobalMux
    port map (
            O => \N__55602\,
            I => \clk_32MHz\
        );

    \I__13660\ : CEMux
    port map (
            O => \N__55599\,
            I => \N__55596\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__55596\,
            I => \N__55593\
        );

    \I__13658\ : Span4Mux_v
    port map (
            O => \N__55593\,
            I => \N__55590\
        );

    \I__13657\ : Span4Mux_h
    port map (
            O => \N__55590\,
            I => \N__55587\
        );

    \I__13656\ : Sp12to4
    port map (
            O => \N__55587\,
            I => \N__55584\
        );

    \I__13655\ : Span12Mux_s10_h
    port map (
            O => \N__55584\,
            I => \N__55581\
        );

    \I__13654\ : Odrv12
    port map (
            O => \N__55581\,
            I => n11600
        );

    \I__13653\ : InMux
    port map (
            O => \N__55578\,
            I => \N__55575\
        );

    \I__13652\ : LocalMux
    port map (
            O => \N__55575\,
            I => \N__55568\
        );

    \I__13651\ : InMux
    port map (
            O => \N__55574\,
            I => \N__55565\
        );

    \I__13650\ : InMux
    port map (
            O => \N__55573\,
            I => \N__55559\
        );

    \I__13649\ : InMux
    port map (
            O => \N__55572\,
            I => \N__55554\
        );

    \I__13648\ : InMux
    port map (
            O => \N__55571\,
            I => \N__55554\
        );

    \I__13647\ : Span4Mux_v
    port map (
            O => \N__55568\,
            I => \N__55548\
        );

    \I__13646\ : LocalMux
    port map (
            O => \N__55565\,
            I => \N__55548\
        );

    \I__13645\ : InMux
    port map (
            O => \N__55564\,
            I => \N__55545\
        );

    \I__13644\ : InMux
    port map (
            O => \N__55563\,
            I => \N__55541\
        );

    \I__13643\ : InMux
    port map (
            O => \N__55562\,
            I => \N__55538\
        );

    \I__13642\ : LocalMux
    port map (
            O => \N__55559\,
            I => \N__55533\
        );

    \I__13641\ : LocalMux
    port map (
            O => \N__55554\,
            I => \N__55530\
        );

    \I__13640\ : InMux
    port map (
            O => \N__55553\,
            I => \N__55527\
        );

    \I__13639\ : Span4Mux_h
    port map (
            O => \N__55548\,
            I => \N__55524\
        );

    \I__13638\ : LocalMux
    port map (
            O => \N__55545\,
            I => \N__55521\
        );

    \I__13637\ : InMux
    port map (
            O => \N__55544\,
            I => \N__55518\
        );

    \I__13636\ : LocalMux
    port map (
            O => \N__55541\,
            I => \N__55513\
        );

    \I__13635\ : LocalMux
    port map (
            O => \N__55538\,
            I => \N__55513\
        );

    \I__13634\ : InMux
    port map (
            O => \N__55537\,
            I => \N__55508\
        );

    \I__13633\ : InMux
    port map (
            O => \N__55536\,
            I => \N__55508\
        );

    \I__13632\ : Span4Mux_h
    port map (
            O => \N__55533\,
            I => \N__55503\
        );

    \I__13631\ : Span4Mux_v
    port map (
            O => \N__55530\,
            I => \N__55503\
        );

    \I__13630\ : LocalMux
    port map (
            O => \N__55527\,
            I => \N__55496\
        );

    \I__13629\ : Span4Mux_v
    port map (
            O => \N__55524\,
            I => \N__55496\
        );

    \I__13628\ : Span4Mux_h
    port map (
            O => \N__55521\,
            I => \N__55496\
        );

    \I__13627\ : LocalMux
    port map (
            O => \N__55518\,
            I => \N__55489\
        );

    \I__13626\ : Span12Mux_v
    port map (
            O => \N__55513\,
            I => \N__55489\
        );

    \I__13625\ : LocalMux
    port map (
            O => \N__55508\,
            I => \N__55489\
        );

    \I__13624\ : Odrv4
    port map (
            O => \N__55503\,
            I => n12433
        );

    \I__13623\ : Odrv4
    port map (
            O => \N__55496\,
            I => n12433
        );

    \I__13622\ : Odrv12
    port map (
            O => \N__55489\,
            I => n12433
        );

    \I__13621\ : CascadeMux
    port map (
            O => \N__55482\,
            I => \n10_adj_1619_cascade_\
        );

    \I__13620\ : CascadeMux
    port map (
            O => \N__55479\,
            I => \N__55475\
        );

    \I__13619\ : SRMux
    port map (
            O => \N__55478\,
            I => \N__55456\
        );

    \I__13618\ : InMux
    port map (
            O => \N__55475\,
            I => \N__55452\
        );

    \I__13617\ : InMux
    port map (
            O => \N__55474\,
            I => \N__55441\
        );

    \I__13616\ : InMux
    port map (
            O => \N__55473\,
            I => \N__55441\
        );

    \I__13615\ : InMux
    port map (
            O => \N__55472\,
            I => \N__55441\
        );

    \I__13614\ : InMux
    port map (
            O => \N__55471\,
            I => \N__55441\
        );

    \I__13613\ : InMux
    port map (
            O => \N__55470\,
            I => \N__55441\
        );

    \I__13612\ : CascadeMux
    port map (
            O => \N__55469\,
            I => \N__55424\
        );

    \I__13611\ : CascadeMux
    port map (
            O => \N__55468\,
            I => \N__55415\
        );

    \I__13610\ : CascadeMux
    port map (
            O => \N__55467\,
            I => \N__55411\
        );

    \I__13609\ : CascadeMux
    port map (
            O => \N__55466\,
            I => \N__55407\
        );

    \I__13608\ : CascadeMux
    port map (
            O => \N__55465\,
            I => \N__55403\
        );

    \I__13607\ : InMux
    port map (
            O => \N__55464\,
            I => \N__55399\
        );

    \I__13606\ : CascadeMux
    port map (
            O => \N__55463\,
            I => \N__55396\
        );

    \I__13605\ : InMux
    port map (
            O => \N__55462\,
            I => \N__55389\
        );

    \I__13604\ : InMux
    port map (
            O => \N__55461\,
            I => \N__55389\
        );

    \I__13603\ : InMux
    port map (
            O => \N__55460\,
            I => \N__55389\
        );

    \I__13602\ : InMux
    port map (
            O => \N__55459\,
            I => \N__55384\
        );

    \I__13601\ : LocalMux
    port map (
            O => \N__55456\,
            I => \N__55381\
        );

    \I__13600\ : InMux
    port map (
            O => \N__55455\,
            I => \N__55378\
        );

    \I__13599\ : LocalMux
    port map (
            O => \N__55452\,
            I => \N__55373\
        );

    \I__13598\ : LocalMux
    port map (
            O => \N__55441\,
            I => \N__55373\
        );

    \I__13597\ : InMux
    port map (
            O => \N__55440\,
            I => \N__55368\
        );

    \I__13596\ : InMux
    port map (
            O => \N__55439\,
            I => \N__55368\
        );

    \I__13595\ : InMux
    port map (
            O => \N__55438\,
            I => \N__55359\
        );

    \I__13594\ : InMux
    port map (
            O => \N__55437\,
            I => \N__55359\
        );

    \I__13593\ : InMux
    port map (
            O => \N__55436\,
            I => \N__55359\
        );

    \I__13592\ : InMux
    port map (
            O => \N__55435\,
            I => \N__55359\
        );

    \I__13591\ : CascadeMux
    port map (
            O => \N__55434\,
            I => \N__55355\
        );

    \I__13590\ : InMux
    port map (
            O => \N__55433\,
            I => \N__55352\
        );

    \I__13589\ : InMux
    port map (
            O => \N__55432\,
            I => \N__55347\
        );

    \I__13588\ : InMux
    port map (
            O => \N__55431\,
            I => \N__55347\
        );

    \I__13587\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55343\
        );

    \I__13586\ : InMux
    port map (
            O => \N__55429\,
            I => \N__55336\
        );

    \I__13585\ : InMux
    port map (
            O => \N__55428\,
            I => \N__55336\
        );

    \I__13584\ : InMux
    port map (
            O => \N__55427\,
            I => \N__55336\
        );

    \I__13583\ : InMux
    port map (
            O => \N__55424\,
            I => \N__55325\
        );

    \I__13582\ : InMux
    port map (
            O => \N__55423\,
            I => \N__55325\
        );

    \I__13581\ : InMux
    port map (
            O => \N__55422\,
            I => \N__55325\
        );

    \I__13580\ : InMux
    port map (
            O => \N__55421\,
            I => \N__55325\
        );

    \I__13579\ : InMux
    port map (
            O => \N__55420\,
            I => \N__55325\
        );

    \I__13578\ : InMux
    port map (
            O => \N__55419\,
            I => \N__55322\
        );

    \I__13577\ : InMux
    port map (
            O => \N__55418\,
            I => \N__55319\
        );

    \I__13576\ : InMux
    port map (
            O => \N__55415\,
            I => \N__55302\
        );

    \I__13575\ : InMux
    port map (
            O => \N__55414\,
            I => \N__55302\
        );

    \I__13574\ : InMux
    port map (
            O => \N__55411\,
            I => \N__55302\
        );

    \I__13573\ : InMux
    port map (
            O => \N__55410\,
            I => \N__55302\
        );

    \I__13572\ : InMux
    port map (
            O => \N__55407\,
            I => \N__55302\
        );

    \I__13571\ : InMux
    port map (
            O => \N__55406\,
            I => \N__55302\
        );

    \I__13570\ : InMux
    port map (
            O => \N__55403\,
            I => \N__55302\
        );

    \I__13569\ : InMux
    port map (
            O => \N__55402\,
            I => \N__55302\
        );

    \I__13568\ : LocalMux
    port map (
            O => \N__55399\,
            I => \N__55299\
        );

    \I__13567\ : InMux
    port map (
            O => \N__55396\,
            I => \N__55289\
        );

    \I__13566\ : LocalMux
    port map (
            O => \N__55389\,
            I => \N__55282\
        );

    \I__13565\ : CascadeMux
    port map (
            O => \N__55388\,
            I => \N__55276\
        );

    \I__13564\ : InMux
    port map (
            O => \N__55387\,
            I => \N__55273\
        );

    \I__13563\ : LocalMux
    port map (
            O => \N__55384\,
            I => \N__55255\
        );

    \I__13562\ : Span4Mux_v
    port map (
            O => \N__55381\,
            I => \N__55255\
        );

    \I__13561\ : LocalMux
    port map (
            O => \N__55378\,
            I => \N__55255\
        );

    \I__13560\ : Span4Mux_v
    port map (
            O => \N__55373\,
            I => \N__55255\
        );

    \I__13559\ : LocalMux
    port map (
            O => \N__55368\,
            I => \N__55255\
        );

    \I__13558\ : LocalMux
    port map (
            O => \N__55359\,
            I => \N__55255\
        );

    \I__13557\ : CascadeMux
    port map (
            O => \N__55358\,
            I => \N__55252\
        );

    \I__13556\ : InMux
    port map (
            O => \N__55355\,
            I => \N__55244\
        );

    \I__13555\ : LocalMux
    port map (
            O => \N__55352\,
            I => \N__55239\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__55347\,
            I => \N__55239\
        );

    \I__13553\ : InMux
    port map (
            O => \N__55346\,
            I => \N__55230\
        );

    \I__13552\ : LocalMux
    port map (
            O => \N__55343\,
            I => \N__55227\
        );

    \I__13551\ : LocalMux
    port map (
            O => \N__55336\,
            I => \N__55216\
        );

    \I__13550\ : LocalMux
    port map (
            O => \N__55325\,
            I => \N__55216\
        );

    \I__13549\ : LocalMux
    port map (
            O => \N__55322\,
            I => \N__55216\
        );

    \I__13548\ : LocalMux
    port map (
            O => \N__55319\,
            I => \N__55216\
        );

    \I__13547\ : LocalMux
    port map (
            O => \N__55302\,
            I => \N__55216\
        );

    \I__13546\ : Span4Mux_v
    port map (
            O => \N__55299\,
            I => \N__55213\
        );

    \I__13545\ : InMux
    port map (
            O => \N__55298\,
            I => \N__55208\
        );

    \I__13544\ : InMux
    port map (
            O => \N__55297\,
            I => \N__55208\
        );

    \I__13543\ : InMux
    port map (
            O => \N__55296\,
            I => \N__55204\
        );

    \I__13542\ : InMux
    port map (
            O => \N__55295\,
            I => \N__55195\
        );

    \I__13541\ : InMux
    port map (
            O => \N__55294\,
            I => \N__55195\
        );

    \I__13540\ : InMux
    port map (
            O => \N__55293\,
            I => \N__55195\
        );

    \I__13539\ : InMux
    port map (
            O => \N__55292\,
            I => \N__55195\
        );

    \I__13538\ : LocalMux
    port map (
            O => \N__55289\,
            I => \N__55192\
        );

    \I__13537\ : InMux
    port map (
            O => \N__55288\,
            I => \N__55187\
        );

    \I__13536\ : InMux
    port map (
            O => \N__55287\,
            I => \N__55187\
        );

    \I__13535\ : InMux
    port map (
            O => \N__55286\,
            I => \N__55184\
        );

    \I__13534\ : CascadeMux
    port map (
            O => \N__55285\,
            I => \N__55177\
        );

    \I__13533\ : Span4Mux_h
    port map (
            O => \N__55282\,
            I => \N__55174\
        );

    \I__13532\ : InMux
    port map (
            O => \N__55281\,
            I => \N__55171\
        );

    \I__13531\ : InMux
    port map (
            O => \N__55280\,
            I => \N__55166\
        );

    \I__13530\ : InMux
    port map (
            O => \N__55279\,
            I => \N__55166\
        );

    \I__13529\ : InMux
    port map (
            O => \N__55276\,
            I => \N__55160\
        );

    \I__13528\ : LocalMux
    port map (
            O => \N__55273\,
            I => \N__55157\
        );

    \I__13527\ : InMux
    port map (
            O => \N__55272\,
            I => \N__55154\
        );

    \I__13526\ : InMux
    port map (
            O => \N__55271\,
            I => \N__55149\
        );

    \I__13525\ : InMux
    port map (
            O => \N__55270\,
            I => \N__55149\
        );

    \I__13524\ : InMux
    port map (
            O => \N__55269\,
            I => \N__55144\
        );

    \I__13523\ : InMux
    port map (
            O => \N__55268\,
            I => \N__55144\
        );

    \I__13522\ : Span4Mux_v
    port map (
            O => \N__55255\,
            I => \N__55141\
        );

    \I__13521\ : InMux
    port map (
            O => \N__55252\,
            I => \N__55136\
        );

    \I__13520\ : InMux
    port map (
            O => \N__55251\,
            I => \N__55136\
        );

    \I__13519\ : InMux
    port map (
            O => \N__55250\,
            I => \N__55131\
        );

    \I__13518\ : InMux
    port map (
            O => \N__55249\,
            I => \N__55131\
        );

    \I__13517\ : InMux
    port map (
            O => \N__55248\,
            I => \N__55126\
        );

    \I__13516\ : InMux
    port map (
            O => \N__55247\,
            I => \N__55126\
        );

    \I__13515\ : LocalMux
    port map (
            O => \N__55244\,
            I => \N__55121\
        );

    \I__13514\ : Span4Mux_v
    port map (
            O => \N__55239\,
            I => \N__55121\
        );

    \I__13513\ : InMux
    port map (
            O => \N__55238\,
            I => \N__55109\
        );

    \I__13512\ : InMux
    port map (
            O => \N__55237\,
            I => \N__55109\
        );

    \I__13511\ : InMux
    port map (
            O => \N__55236\,
            I => \N__55109\
        );

    \I__13510\ : InMux
    port map (
            O => \N__55235\,
            I => \N__55109\
        );

    \I__13509\ : InMux
    port map (
            O => \N__55234\,
            I => \N__55109\
        );

    \I__13508\ : InMux
    port map (
            O => \N__55233\,
            I => \N__55105\
        );

    \I__13507\ : LocalMux
    port map (
            O => \N__55230\,
            I => \N__55101\
        );

    \I__13506\ : Span4Mux_h
    port map (
            O => \N__55227\,
            I => \N__55096\
        );

    \I__13505\ : Span4Mux_v
    port map (
            O => \N__55216\,
            I => \N__55096\
        );

    \I__13504\ : Span4Mux_h
    port map (
            O => \N__55213\,
            I => \N__55091\
        );

    \I__13503\ : LocalMux
    port map (
            O => \N__55208\,
            I => \N__55091\
        );

    \I__13502\ : InMux
    port map (
            O => \N__55207\,
            I => \N__55088\
        );

    \I__13501\ : LocalMux
    port map (
            O => \N__55204\,
            I => \N__55085\
        );

    \I__13500\ : LocalMux
    port map (
            O => \N__55195\,
            I => \N__55076\
        );

    \I__13499\ : Span4Mux_v
    port map (
            O => \N__55192\,
            I => \N__55076\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__55187\,
            I => \N__55076\
        );

    \I__13497\ : LocalMux
    port map (
            O => \N__55184\,
            I => \N__55076\
        );

    \I__13496\ : InMux
    port map (
            O => \N__55183\,
            I => \N__55069\
        );

    \I__13495\ : InMux
    port map (
            O => \N__55182\,
            I => \N__55069\
        );

    \I__13494\ : InMux
    port map (
            O => \N__55181\,
            I => \N__55069\
        );

    \I__13493\ : InMux
    port map (
            O => \N__55180\,
            I => \N__55062\
        );

    \I__13492\ : InMux
    port map (
            O => \N__55177\,
            I => \N__55059\
        );

    \I__13491\ : Span4Mux_h
    port map (
            O => \N__55174\,
            I => \N__55056\
        );

    \I__13490\ : LocalMux
    port map (
            O => \N__55171\,
            I => \N__55051\
        );

    \I__13489\ : LocalMux
    port map (
            O => \N__55166\,
            I => \N__55051\
        );

    \I__13488\ : InMux
    port map (
            O => \N__55165\,
            I => \N__55044\
        );

    \I__13487\ : InMux
    port map (
            O => \N__55164\,
            I => \N__55044\
        );

    \I__13486\ : InMux
    port map (
            O => \N__55163\,
            I => \N__55044\
        );

    \I__13485\ : LocalMux
    port map (
            O => \N__55160\,
            I => \N__55033\
        );

    \I__13484\ : Span4Mux_v
    port map (
            O => \N__55157\,
            I => \N__55033\
        );

    \I__13483\ : LocalMux
    port map (
            O => \N__55154\,
            I => \N__55033\
        );

    \I__13482\ : LocalMux
    port map (
            O => \N__55149\,
            I => \N__55033\
        );

    \I__13481\ : LocalMux
    port map (
            O => \N__55144\,
            I => \N__55033\
        );

    \I__13480\ : Span4Mux_h
    port map (
            O => \N__55141\,
            I => \N__55030\
        );

    \I__13479\ : LocalMux
    port map (
            O => \N__55136\,
            I => \N__55024\
        );

    \I__13478\ : LocalMux
    port map (
            O => \N__55131\,
            I => \N__55017\
        );

    \I__13477\ : LocalMux
    port map (
            O => \N__55126\,
            I => \N__55017\
        );

    \I__13476\ : Span4Mux_h
    port map (
            O => \N__55121\,
            I => \N__55017\
        );

    \I__13475\ : InMux
    port map (
            O => \N__55120\,
            I => \N__55014\
        );

    \I__13474\ : LocalMux
    port map (
            O => \N__55109\,
            I => \N__55011\
        );

    \I__13473\ : InMux
    port map (
            O => \N__55108\,
            I => \N__55008\
        );

    \I__13472\ : LocalMux
    port map (
            O => \N__55105\,
            I => \N__55005\
        );

    \I__13471\ : InMux
    port map (
            O => \N__55104\,
            I => \N__55002\
        );

    \I__13470\ : Span4Mux_v
    port map (
            O => \N__55101\,
            I => \N__54995\
        );

    \I__13469\ : Span4Mux_h
    port map (
            O => \N__55096\,
            I => \N__54995\
        );

    \I__13468\ : Span4Mux_v
    port map (
            O => \N__55091\,
            I => \N__54995\
        );

    \I__13467\ : LocalMux
    port map (
            O => \N__55088\,
            I => \N__54990\
        );

    \I__13466\ : Span4Mux_v
    port map (
            O => \N__55085\,
            I => \N__54990\
        );

    \I__13465\ : Span4Mux_v
    port map (
            O => \N__55076\,
            I => \N__54985\
        );

    \I__13464\ : LocalMux
    port map (
            O => \N__55069\,
            I => \N__54985\
        );

    \I__13463\ : InMux
    port map (
            O => \N__55068\,
            I => \N__54980\
        );

    \I__13462\ : InMux
    port map (
            O => \N__55067\,
            I => \N__54980\
        );

    \I__13461\ : InMux
    port map (
            O => \N__55066\,
            I => \N__54977\
        );

    \I__13460\ : InMux
    port map (
            O => \N__55065\,
            I => \N__54974\
        );

    \I__13459\ : LocalMux
    port map (
            O => \N__55062\,
            I => \N__54965\
        );

    \I__13458\ : LocalMux
    port map (
            O => \N__55059\,
            I => \N__54965\
        );

    \I__13457\ : Span4Mux_h
    port map (
            O => \N__55056\,
            I => \N__54965\
        );

    \I__13456\ : Span4Mux_v
    port map (
            O => \N__55051\,
            I => \N__54965\
        );

    \I__13455\ : LocalMux
    port map (
            O => \N__55044\,
            I => \N__54958\
        );

    \I__13454\ : Span4Mux_v
    port map (
            O => \N__55033\,
            I => \N__54958\
        );

    \I__13453\ : Span4Mux_h
    port map (
            O => \N__55030\,
            I => \N__54958\
        );

    \I__13452\ : InMux
    port map (
            O => \N__55029\,
            I => \N__54951\
        );

    \I__13451\ : InMux
    port map (
            O => \N__55028\,
            I => \N__54951\
        );

    \I__13450\ : InMux
    port map (
            O => \N__55027\,
            I => \N__54951\
        );

    \I__13449\ : Span4Mux_v
    port map (
            O => \N__55024\,
            I => \N__54946\
        );

    \I__13448\ : Span4Mux_v
    port map (
            O => \N__55017\,
            I => \N__54946\
        );

    \I__13447\ : LocalMux
    port map (
            O => \N__55014\,
            I => \N__54941\
        );

    \I__13446\ : Span4Mux_h
    port map (
            O => \N__55011\,
            I => \N__54941\
        );

    \I__13445\ : LocalMux
    port map (
            O => \N__55008\,
            I => \N__54934\
        );

    \I__13444\ : Span12Mux_v
    port map (
            O => \N__55005\,
            I => \N__54934\
        );

    \I__13443\ : LocalMux
    port map (
            O => \N__55002\,
            I => \N__54934\
        );

    \I__13442\ : Span4Mux_h
    port map (
            O => \N__54995\,
            I => \N__54931\
        );

    \I__13441\ : Span4Mux_h
    port map (
            O => \N__54990\,
            I => \N__54924\
        );

    \I__13440\ : Span4Mux_v
    port map (
            O => \N__54985\,
            I => \N__54924\
        );

    \I__13439\ : LocalMux
    port map (
            O => \N__54980\,
            I => \N__54924\
        );

    \I__13438\ : LocalMux
    port map (
            O => \N__54977\,
            I => comm_state_3
        );

    \I__13437\ : LocalMux
    port map (
            O => \N__54974\,
            I => comm_state_3
        );

    \I__13436\ : Odrv4
    port map (
            O => \N__54965\,
            I => comm_state_3
        );

    \I__13435\ : Odrv4
    port map (
            O => \N__54958\,
            I => comm_state_3
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__54951\,
            I => comm_state_3
        );

    \I__13433\ : Odrv4
    port map (
            O => \N__54946\,
            I => comm_state_3
        );

    \I__13432\ : Odrv4
    port map (
            O => \N__54941\,
            I => comm_state_3
        );

    \I__13431\ : Odrv12
    port map (
            O => \N__54934\,
            I => comm_state_3
        );

    \I__13430\ : Odrv4
    port map (
            O => \N__54931\,
            I => comm_state_3
        );

    \I__13429\ : Odrv4
    port map (
            O => \N__54924\,
            I => comm_state_3
        );

    \I__13428\ : CEMux
    port map (
            O => \N__54903\,
            I => \N__54900\
        );

    \I__13427\ : LocalMux
    port map (
            O => \N__54900\,
            I => \N__54897\
        );

    \I__13426\ : Odrv12
    port map (
            O => \N__54897\,
            I => n12079
        );

    \I__13425\ : CascadeMux
    port map (
            O => \N__54894\,
            I => \N__54888\
        );

    \I__13424\ : InMux
    port map (
            O => \N__54893\,
            I => \N__54881\
        );

    \I__13423\ : InMux
    port map (
            O => \N__54892\,
            I => \N__54876\
        );

    \I__13422\ : InMux
    port map (
            O => \N__54891\,
            I => \N__54876\
        );

    \I__13421\ : InMux
    port map (
            O => \N__54888\,
            I => \N__54871\
        );

    \I__13420\ : InMux
    port map (
            O => \N__54887\,
            I => \N__54864\
        );

    \I__13419\ : InMux
    port map (
            O => \N__54886\,
            I => \N__54864\
        );

    \I__13418\ : InMux
    port map (
            O => \N__54885\,
            I => \N__54864\
        );

    \I__13417\ : InMux
    port map (
            O => \N__54884\,
            I => \N__54854\
        );

    \I__13416\ : LocalMux
    port map (
            O => \N__54881\,
            I => \N__54848\
        );

    \I__13415\ : LocalMux
    port map (
            O => \N__54876\,
            I => \N__54844\
        );

    \I__13414\ : InMux
    port map (
            O => \N__54875\,
            I => \N__54836\
        );

    \I__13413\ : InMux
    port map (
            O => \N__54874\,
            I => \N__54833\
        );

    \I__13412\ : LocalMux
    port map (
            O => \N__54871\,
            I => \N__54828\
        );

    \I__13411\ : LocalMux
    port map (
            O => \N__54864\,
            I => \N__54828\
        );

    \I__13410\ : InMux
    port map (
            O => \N__54863\,
            I => \N__54822\
        );

    \I__13409\ : InMux
    port map (
            O => \N__54862\,
            I => \N__54811\
        );

    \I__13408\ : InMux
    port map (
            O => \N__54861\,
            I => \N__54811\
        );

    \I__13407\ : InMux
    port map (
            O => \N__54860\,
            I => \N__54811\
        );

    \I__13406\ : InMux
    port map (
            O => \N__54859\,
            I => \N__54811\
        );

    \I__13405\ : InMux
    port map (
            O => \N__54858\,
            I => \N__54811\
        );

    \I__13404\ : InMux
    port map (
            O => \N__54857\,
            I => \N__54807\
        );

    \I__13403\ : LocalMux
    port map (
            O => \N__54854\,
            I => \N__54804\
        );

    \I__13402\ : CascadeMux
    port map (
            O => \N__54853\,
            I => \N__54800\
        );

    \I__13401\ : CascadeMux
    port map (
            O => \N__54852\,
            I => \N__54797\
        );

    \I__13400\ : InMux
    port map (
            O => \N__54851\,
            I => \N__54792\
        );

    \I__13399\ : Span4Mux_h
    port map (
            O => \N__54848\,
            I => \N__54789\
        );

    \I__13398\ : InMux
    port map (
            O => \N__54847\,
            I => \N__54784\
        );

    \I__13397\ : Span4Mux_h
    port map (
            O => \N__54844\,
            I => \N__54781\
        );

    \I__13396\ : InMux
    port map (
            O => \N__54843\,
            I => \N__54778\
        );

    \I__13395\ : CascadeMux
    port map (
            O => \N__54842\,
            I => \N__54774\
        );

    \I__13394\ : InMux
    port map (
            O => \N__54841\,
            I => \N__54771\
        );

    \I__13393\ : InMux
    port map (
            O => \N__54840\,
            I => \N__54766\
        );

    \I__13392\ : InMux
    port map (
            O => \N__54839\,
            I => \N__54766\
        );

    \I__13391\ : LocalMux
    port map (
            O => \N__54836\,
            I => \N__54761\
        );

    \I__13390\ : LocalMux
    port map (
            O => \N__54833\,
            I => \N__54761\
        );

    \I__13389\ : Span4Mux_v
    port map (
            O => \N__54828\,
            I => \N__54758\
        );

    \I__13388\ : InMux
    port map (
            O => \N__54827\,
            I => \N__54755\
        );

    \I__13387\ : InMux
    port map (
            O => \N__54826\,
            I => \N__54750\
        );

    \I__13386\ : InMux
    port map (
            O => \N__54825\,
            I => \N__54747\
        );

    \I__13385\ : LocalMux
    port map (
            O => \N__54822\,
            I => \N__54744\
        );

    \I__13384\ : LocalMux
    port map (
            O => \N__54811\,
            I => \N__54741\
        );

    \I__13383\ : CascadeMux
    port map (
            O => \N__54810\,
            I => \N__54734\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__54807\,
            I => \N__54731\
        );

    \I__13381\ : Span4Mux_v
    port map (
            O => \N__54804\,
            I => \N__54728\
        );

    \I__13380\ : InMux
    port map (
            O => \N__54803\,
            I => \N__54725\
        );

    \I__13379\ : InMux
    port map (
            O => \N__54800\,
            I => \N__54716\
        );

    \I__13378\ : InMux
    port map (
            O => \N__54797\,
            I => \N__54716\
        );

    \I__13377\ : InMux
    port map (
            O => \N__54796\,
            I => \N__54716\
        );

    \I__13376\ : InMux
    port map (
            O => \N__54795\,
            I => \N__54716\
        );

    \I__13375\ : LocalMux
    port map (
            O => \N__54792\,
            I => \N__54711\
        );

    \I__13374\ : Span4Mux_h
    port map (
            O => \N__54789\,
            I => \N__54711\
        );

    \I__13373\ : CascadeMux
    port map (
            O => \N__54788\,
            I => \N__54707\
        );

    \I__13372\ : InMux
    port map (
            O => \N__54787\,
            I => \N__54703\
        );

    \I__13371\ : LocalMux
    port map (
            O => \N__54784\,
            I => \N__54696\
        );

    \I__13370\ : Span4Mux_v
    port map (
            O => \N__54781\,
            I => \N__54696\
        );

    \I__13369\ : LocalMux
    port map (
            O => \N__54778\,
            I => \N__54696\
        );

    \I__13368\ : InMux
    port map (
            O => \N__54777\,
            I => \N__54691\
        );

    \I__13367\ : InMux
    port map (
            O => \N__54774\,
            I => \N__54691\
        );

    \I__13366\ : LocalMux
    port map (
            O => \N__54771\,
            I => \N__54686\
        );

    \I__13365\ : LocalMux
    port map (
            O => \N__54766\,
            I => \N__54686\
        );

    \I__13364\ : Span4Mux_v
    port map (
            O => \N__54761\,
            I => \N__54680\
        );

    \I__13363\ : Span4Mux_h
    port map (
            O => \N__54758\,
            I => \N__54675\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__54755\,
            I => \N__54675\
        );

    \I__13361\ : InMux
    port map (
            O => \N__54754\,
            I => \N__54670\
        );

    \I__13360\ : InMux
    port map (
            O => \N__54753\,
            I => \N__54670\
        );

    \I__13359\ : LocalMux
    port map (
            O => \N__54750\,
            I => \N__54667\
        );

    \I__13358\ : LocalMux
    port map (
            O => \N__54747\,
            I => \N__54662\
        );

    \I__13357\ : Span4Mux_v
    port map (
            O => \N__54744\,
            I => \N__54662\
        );

    \I__13356\ : Span4Mux_h
    port map (
            O => \N__54741\,
            I => \N__54659\
        );

    \I__13355\ : InMux
    port map (
            O => \N__54740\,
            I => \N__54652\
        );

    \I__13354\ : InMux
    port map (
            O => \N__54739\,
            I => \N__54652\
        );

    \I__13353\ : InMux
    port map (
            O => \N__54738\,
            I => \N__54652\
        );

    \I__13352\ : InMux
    port map (
            O => \N__54737\,
            I => \N__54649\
        );

    \I__13351\ : InMux
    port map (
            O => \N__54734\,
            I => \N__54646\
        );

    \I__13350\ : Span12Mux_h
    port map (
            O => \N__54731\,
            I => \N__54643\
        );

    \I__13349\ : Span4Mux_h
    port map (
            O => \N__54728\,
            I => \N__54640\
        );

    \I__13348\ : LocalMux
    port map (
            O => \N__54725\,
            I => \N__54633\
        );

    \I__13347\ : LocalMux
    port map (
            O => \N__54716\,
            I => \N__54633\
        );

    \I__13346\ : Span4Mux_h
    port map (
            O => \N__54711\,
            I => \N__54633\
        );

    \I__13345\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54626\
        );

    \I__13344\ : InMux
    port map (
            O => \N__54707\,
            I => \N__54626\
        );

    \I__13343\ : InMux
    port map (
            O => \N__54706\,
            I => \N__54626\
        );

    \I__13342\ : LocalMux
    port map (
            O => \N__54703\,
            I => \N__54617\
        );

    \I__13341\ : Span4Mux_v
    port map (
            O => \N__54696\,
            I => \N__54617\
        );

    \I__13340\ : LocalMux
    port map (
            O => \N__54691\,
            I => \N__54617\
        );

    \I__13339\ : Span4Mux_v
    port map (
            O => \N__54686\,
            I => \N__54617\
        );

    \I__13338\ : InMux
    port map (
            O => \N__54685\,
            I => \N__54610\
        );

    \I__13337\ : InMux
    port map (
            O => \N__54684\,
            I => \N__54610\
        );

    \I__13336\ : InMux
    port map (
            O => \N__54683\,
            I => \N__54610\
        );

    \I__13335\ : Span4Mux_h
    port map (
            O => \N__54680\,
            I => \N__54603\
        );

    \I__13334\ : Span4Mux_v
    port map (
            O => \N__54675\,
            I => \N__54603\
        );

    \I__13333\ : LocalMux
    port map (
            O => \N__54670\,
            I => \N__54603\
        );

    \I__13332\ : Span4Mux_v
    port map (
            O => \N__54667\,
            I => \N__54594\
        );

    \I__13331\ : Span4Mux_h
    port map (
            O => \N__54662\,
            I => \N__54594\
        );

    \I__13330\ : Span4Mux_v
    port map (
            O => \N__54659\,
            I => \N__54594\
        );

    \I__13329\ : LocalMux
    port map (
            O => \N__54652\,
            I => \N__54594\
        );

    \I__13328\ : LocalMux
    port map (
            O => \N__54649\,
            I => comm_state_2
        );

    \I__13327\ : LocalMux
    port map (
            O => \N__54646\,
            I => comm_state_2
        );

    \I__13326\ : Odrv12
    port map (
            O => \N__54643\,
            I => comm_state_2
        );

    \I__13325\ : Odrv4
    port map (
            O => \N__54640\,
            I => comm_state_2
        );

    \I__13324\ : Odrv4
    port map (
            O => \N__54633\,
            I => comm_state_2
        );

    \I__13323\ : LocalMux
    port map (
            O => \N__54626\,
            I => comm_state_2
        );

    \I__13322\ : Odrv4
    port map (
            O => \N__54617\,
            I => comm_state_2
        );

    \I__13321\ : LocalMux
    port map (
            O => \N__54610\,
            I => comm_state_2
        );

    \I__13320\ : Odrv4
    port map (
            O => \N__54603\,
            I => comm_state_2
        );

    \I__13319\ : Odrv4
    port map (
            O => \N__54594\,
            I => comm_state_2
        );

    \I__13318\ : InMux
    port map (
            O => \N__54573\,
            I => \N__54568\
        );

    \I__13317\ : InMux
    port map (
            O => \N__54572\,
            I => \N__54563\
        );

    \I__13316\ : InMux
    port map (
            O => \N__54571\,
            I => \N__54560\
        );

    \I__13315\ : LocalMux
    port map (
            O => \N__54568\,
            I => \N__54557\
        );

    \I__13314\ : InMux
    port map (
            O => \N__54567\,
            I => \N__54538\
        );

    \I__13313\ : InMux
    port map (
            O => \N__54566\,
            I => \N__54535\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__54563\,
            I => \N__54531\
        );

    \I__13311\ : LocalMux
    port map (
            O => \N__54560\,
            I => \N__54526\
        );

    \I__13310\ : Span4Mux_v
    port map (
            O => \N__54557\,
            I => \N__54526\
        );

    \I__13309\ : InMux
    port map (
            O => \N__54556\,
            I => \N__54522\
        );

    \I__13308\ : InMux
    port map (
            O => \N__54555\,
            I => \N__54519\
        );

    \I__13307\ : InMux
    port map (
            O => \N__54554\,
            I => \N__54511\
        );

    \I__13306\ : InMux
    port map (
            O => \N__54553\,
            I => \N__54495\
        );

    \I__13305\ : CascadeMux
    port map (
            O => \N__54552\,
            I => \N__54491\
        );

    \I__13304\ : InMux
    port map (
            O => \N__54551\,
            I => \N__54467\
        );

    \I__13303\ : InMux
    port map (
            O => \N__54550\,
            I => \N__54467\
        );

    \I__13302\ : InMux
    port map (
            O => \N__54549\,
            I => \N__54467\
        );

    \I__13301\ : InMux
    port map (
            O => \N__54548\,
            I => \N__54467\
        );

    \I__13300\ : InMux
    port map (
            O => \N__54547\,
            I => \N__54467\
        );

    \I__13299\ : InMux
    port map (
            O => \N__54546\,
            I => \N__54467\
        );

    \I__13298\ : InMux
    port map (
            O => \N__54545\,
            I => \N__54467\
        );

    \I__13297\ : InMux
    port map (
            O => \N__54544\,
            I => \N__54467\
        );

    \I__13296\ : InMux
    port map (
            O => \N__54543\,
            I => \N__54464\
        );

    \I__13295\ : InMux
    port map (
            O => \N__54542\,
            I => \N__54461\
        );

    \I__13294\ : InMux
    port map (
            O => \N__54541\,
            I => \N__54458\
        );

    \I__13293\ : LocalMux
    port map (
            O => \N__54538\,
            I => \N__54455\
        );

    \I__13292\ : LocalMux
    port map (
            O => \N__54535\,
            I => \N__54452\
        );

    \I__13291\ : InMux
    port map (
            O => \N__54534\,
            I => \N__54449\
        );

    \I__13290\ : Span4Mux_h
    port map (
            O => \N__54531\,
            I => \N__54444\
        );

    \I__13289\ : Span4Mux_h
    port map (
            O => \N__54526\,
            I => \N__54444\
        );

    \I__13288\ : InMux
    port map (
            O => \N__54525\,
            I => \N__54441\
        );

    \I__13287\ : LocalMux
    port map (
            O => \N__54522\,
            I => \N__54426\
        );

    \I__13286\ : LocalMux
    port map (
            O => \N__54519\,
            I => \N__54423\
        );

    \I__13285\ : InMux
    port map (
            O => \N__54518\,
            I => \N__54418\
        );

    \I__13284\ : InMux
    port map (
            O => \N__54517\,
            I => \N__54418\
        );

    \I__13283\ : InMux
    port map (
            O => \N__54516\,
            I => \N__54414\
        );

    \I__13282\ : CascadeMux
    port map (
            O => \N__54515\,
            I => \N__54411\
        );

    \I__13281\ : InMux
    port map (
            O => \N__54514\,
            I => \N__54406\
        );

    \I__13280\ : LocalMux
    port map (
            O => \N__54511\,
            I => \N__54403\
        );

    \I__13279\ : InMux
    port map (
            O => \N__54510\,
            I => \N__54397\
        );

    \I__13278\ : InMux
    port map (
            O => \N__54509\,
            I => \N__54390\
        );

    \I__13277\ : InMux
    port map (
            O => \N__54508\,
            I => \N__54390\
        );

    \I__13276\ : InMux
    port map (
            O => \N__54507\,
            I => \N__54390\
        );

    \I__13275\ : InMux
    port map (
            O => \N__54506\,
            I => \N__54381\
        );

    \I__13274\ : InMux
    port map (
            O => \N__54505\,
            I => \N__54381\
        );

    \I__13273\ : InMux
    port map (
            O => \N__54504\,
            I => \N__54381\
        );

    \I__13272\ : InMux
    port map (
            O => \N__54503\,
            I => \N__54381\
        );

    \I__13271\ : CascadeMux
    port map (
            O => \N__54502\,
            I => \N__54376\
        );

    \I__13270\ : InMux
    port map (
            O => \N__54501\,
            I => \N__54371\
        );

    \I__13269\ : InMux
    port map (
            O => \N__54500\,
            I => \N__54368\
        );

    \I__13268\ : InMux
    port map (
            O => \N__54499\,
            I => \N__54363\
        );

    \I__13267\ : InMux
    port map (
            O => \N__54498\,
            I => \N__54360\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__54495\,
            I => \N__54357\
        );

    \I__13265\ : InMux
    port map (
            O => \N__54494\,
            I => \N__54350\
        );

    \I__13264\ : InMux
    port map (
            O => \N__54491\,
            I => \N__54350\
        );

    \I__13263\ : InMux
    port map (
            O => \N__54490\,
            I => \N__54350\
        );

    \I__13262\ : InMux
    port map (
            O => \N__54489\,
            I => \N__54343\
        );

    \I__13261\ : InMux
    port map (
            O => \N__54488\,
            I => \N__54343\
        );

    \I__13260\ : InMux
    port map (
            O => \N__54487\,
            I => \N__54343\
        );

    \I__13259\ : InMux
    port map (
            O => \N__54486\,
            I => \N__54326\
        );

    \I__13258\ : InMux
    port map (
            O => \N__54485\,
            I => \N__54326\
        );

    \I__13257\ : InMux
    port map (
            O => \N__54484\,
            I => \N__54323\
        );

    \I__13256\ : LocalMux
    port map (
            O => \N__54467\,
            I => \N__54308\
        );

    \I__13255\ : LocalMux
    port map (
            O => \N__54464\,
            I => \N__54308\
        );

    \I__13254\ : LocalMux
    port map (
            O => \N__54461\,
            I => \N__54308\
        );

    \I__13253\ : LocalMux
    port map (
            O => \N__54458\,
            I => \N__54308\
        );

    \I__13252\ : Span4Mux_h
    port map (
            O => \N__54455\,
            I => \N__54308\
        );

    \I__13251\ : Span4Mux_v
    port map (
            O => \N__54452\,
            I => \N__54308\
        );

    \I__13250\ : LocalMux
    port map (
            O => \N__54449\,
            I => \N__54308\
        );

    \I__13249\ : Span4Mux_h
    port map (
            O => \N__54444\,
            I => \N__54303\
        );

    \I__13248\ : LocalMux
    port map (
            O => \N__54441\,
            I => \N__54303\
        );

    \I__13247\ : InMux
    port map (
            O => \N__54440\,
            I => \N__54300\
        );

    \I__13246\ : InMux
    port map (
            O => \N__54439\,
            I => \N__54293\
        );

    \I__13245\ : InMux
    port map (
            O => \N__54438\,
            I => \N__54293\
        );

    \I__13244\ : InMux
    port map (
            O => \N__54437\,
            I => \N__54293\
        );

    \I__13243\ : InMux
    port map (
            O => \N__54436\,
            I => \N__54276\
        );

    \I__13242\ : InMux
    port map (
            O => \N__54435\,
            I => \N__54276\
        );

    \I__13241\ : InMux
    port map (
            O => \N__54434\,
            I => \N__54276\
        );

    \I__13240\ : InMux
    port map (
            O => \N__54433\,
            I => \N__54276\
        );

    \I__13239\ : InMux
    port map (
            O => \N__54432\,
            I => \N__54276\
        );

    \I__13238\ : InMux
    port map (
            O => \N__54431\,
            I => \N__54276\
        );

    \I__13237\ : InMux
    port map (
            O => \N__54430\,
            I => \N__54276\
        );

    \I__13236\ : InMux
    port map (
            O => \N__54429\,
            I => \N__54276\
        );

    \I__13235\ : Span4Mux_v
    port map (
            O => \N__54426\,
            I => \N__54269\
        );

    \I__13234\ : Span4Mux_h
    port map (
            O => \N__54423\,
            I => \N__54269\
        );

    \I__13233\ : LocalMux
    port map (
            O => \N__54418\,
            I => \N__54269\
        );

    \I__13232\ : InMux
    port map (
            O => \N__54417\,
            I => \N__54266\
        );

    \I__13231\ : LocalMux
    port map (
            O => \N__54414\,
            I => \N__54263\
        );

    \I__13230\ : InMux
    port map (
            O => \N__54411\,
            I => \N__54256\
        );

    \I__13229\ : InMux
    port map (
            O => \N__54410\,
            I => \N__54256\
        );

    \I__13228\ : InMux
    port map (
            O => \N__54409\,
            I => \N__54256\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__54406\,
            I => \N__54251\
        );

    \I__13226\ : Span4Mux_v
    port map (
            O => \N__54403\,
            I => \N__54251\
        );

    \I__13225\ : InMux
    port map (
            O => \N__54402\,
            I => \N__54248\
        );

    \I__13224\ : InMux
    port map (
            O => \N__54401\,
            I => \N__54245\
        );

    \I__13223\ : InMux
    port map (
            O => \N__54400\,
            I => \N__54242\
        );

    \I__13222\ : LocalMux
    port map (
            O => \N__54397\,
            I => \N__54235\
        );

    \I__13221\ : LocalMux
    port map (
            O => \N__54390\,
            I => \N__54235\
        );

    \I__13220\ : LocalMux
    port map (
            O => \N__54381\,
            I => \N__54235\
        );

    \I__13219\ : InMux
    port map (
            O => \N__54380\,
            I => \N__54232\
        );

    \I__13218\ : InMux
    port map (
            O => \N__54379\,
            I => \N__54225\
        );

    \I__13217\ : InMux
    port map (
            O => \N__54376\,
            I => \N__54225\
        );

    \I__13216\ : InMux
    port map (
            O => \N__54375\,
            I => \N__54225\
        );

    \I__13215\ : InMux
    port map (
            O => \N__54374\,
            I => \N__54222\
        );

    \I__13214\ : LocalMux
    port map (
            O => \N__54371\,
            I => \N__54217\
        );

    \I__13213\ : LocalMux
    port map (
            O => \N__54368\,
            I => \N__54217\
        );

    \I__13212\ : InMux
    port map (
            O => \N__54367\,
            I => \N__54212\
        );

    \I__13211\ : InMux
    port map (
            O => \N__54366\,
            I => \N__54212\
        );

    \I__13210\ : LocalMux
    port map (
            O => \N__54363\,
            I => \N__54201\
        );

    \I__13209\ : LocalMux
    port map (
            O => \N__54360\,
            I => \N__54201\
        );

    \I__13208\ : Span4Mux_v
    port map (
            O => \N__54357\,
            I => \N__54201\
        );

    \I__13207\ : LocalMux
    port map (
            O => \N__54350\,
            I => \N__54201\
        );

    \I__13206\ : LocalMux
    port map (
            O => \N__54343\,
            I => \N__54201\
        );

    \I__13205\ : InMux
    port map (
            O => \N__54342\,
            I => \N__54188\
        );

    \I__13204\ : InMux
    port map (
            O => \N__54341\,
            I => \N__54185\
        );

    \I__13203\ : CascadeMux
    port map (
            O => \N__54340\,
            I => \N__54180\
        );

    \I__13202\ : CascadeMux
    port map (
            O => \N__54339\,
            I => \N__54174\
        );

    \I__13201\ : InMux
    port map (
            O => \N__54338\,
            I => \N__54155\
        );

    \I__13200\ : InMux
    port map (
            O => \N__54337\,
            I => \N__54155\
        );

    \I__13199\ : InMux
    port map (
            O => \N__54336\,
            I => \N__54155\
        );

    \I__13198\ : InMux
    port map (
            O => \N__54335\,
            I => \N__54155\
        );

    \I__13197\ : InMux
    port map (
            O => \N__54334\,
            I => \N__54155\
        );

    \I__13196\ : InMux
    port map (
            O => \N__54333\,
            I => \N__54155\
        );

    \I__13195\ : InMux
    port map (
            O => \N__54332\,
            I => \N__54155\
        );

    \I__13194\ : InMux
    port map (
            O => \N__54331\,
            I => \N__54155\
        );

    \I__13193\ : LocalMux
    port map (
            O => \N__54326\,
            I => \N__54152\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__54323\,
            I => \N__54141\
        );

    \I__13191\ : Span4Mux_v
    port map (
            O => \N__54308\,
            I => \N__54141\
        );

    \I__13190\ : Span4Mux_h
    port map (
            O => \N__54303\,
            I => \N__54141\
        );

    \I__13189\ : LocalMux
    port map (
            O => \N__54300\,
            I => \N__54141\
        );

    \I__13188\ : LocalMux
    port map (
            O => \N__54293\,
            I => \N__54141\
        );

    \I__13187\ : LocalMux
    port map (
            O => \N__54276\,
            I => \N__54136\
        );

    \I__13186\ : Span4Mux_h
    port map (
            O => \N__54269\,
            I => \N__54136\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__54266\,
            I => \N__54129\
        );

    \I__13184\ : Span4Mux_v
    port map (
            O => \N__54263\,
            I => \N__54129\
        );

    \I__13183\ : LocalMux
    port map (
            O => \N__54256\,
            I => \N__54129\
        );

    \I__13182\ : Sp12to4
    port map (
            O => \N__54251\,
            I => \N__54126\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__54248\,
            I => \N__54115\
        );

    \I__13180\ : LocalMux
    port map (
            O => \N__54245\,
            I => \N__54115\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__54242\,
            I => \N__54115\
        );

    \I__13178\ : Sp12to4
    port map (
            O => \N__54235\,
            I => \N__54115\
        );

    \I__13177\ : LocalMux
    port map (
            O => \N__54232\,
            I => \N__54115\
        );

    \I__13176\ : LocalMux
    port map (
            O => \N__54225\,
            I => \N__54112\
        );

    \I__13175\ : LocalMux
    port map (
            O => \N__54222\,
            I => \N__54103\
        );

    \I__13174\ : Span4Mux_h
    port map (
            O => \N__54217\,
            I => \N__54103\
        );

    \I__13173\ : LocalMux
    port map (
            O => \N__54212\,
            I => \N__54103\
        );

    \I__13172\ : Span4Mux_v
    port map (
            O => \N__54201\,
            I => \N__54103\
        );

    \I__13171\ : InMux
    port map (
            O => \N__54200\,
            I => \N__54086\
        );

    \I__13170\ : InMux
    port map (
            O => \N__54199\,
            I => \N__54086\
        );

    \I__13169\ : InMux
    port map (
            O => \N__54198\,
            I => \N__54086\
        );

    \I__13168\ : InMux
    port map (
            O => \N__54197\,
            I => \N__54086\
        );

    \I__13167\ : InMux
    port map (
            O => \N__54196\,
            I => \N__54086\
        );

    \I__13166\ : InMux
    port map (
            O => \N__54195\,
            I => \N__54086\
        );

    \I__13165\ : InMux
    port map (
            O => \N__54194\,
            I => \N__54086\
        );

    \I__13164\ : InMux
    port map (
            O => \N__54193\,
            I => \N__54086\
        );

    \I__13163\ : InMux
    port map (
            O => \N__54192\,
            I => \N__54081\
        );

    \I__13162\ : InMux
    port map (
            O => \N__54191\,
            I => \N__54081\
        );

    \I__13161\ : LocalMux
    port map (
            O => \N__54188\,
            I => \N__54078\
        );

    \I__13160\ : LocalMux
    port map (
            O => \N__54185\,
            I => \N__54075\
        );

    \I__13159\ : InMux
    port map (
            O => \N__54184\,
            I => \N__54068\
        );

    \I__13158\ : InMux
    port map (
            O => \N__54183\,
            I => \N__54068\
        );

    \I__13157\ : InMux
    port map (
            O => \N__54180\,
            I => \N__54068\
        );

    \I__13156\ : InMux
    port map (
            O => \N__54179\,
            I => \N__54063\
        );

    \I__13155\ : InMux
    port map (
            O => \N__54178\,
            I => \N__54063\
        );

    \I__13154\ : InMux
    port map (
            O => \N__54177\,
            I => \N__54054\
        );

    \I__13153\ : InMux
    port map (
            O => \N__54174\,
            I => \N__54054\
        );

    \I__13152\ : InMux
    port map (
            O => \N__54173\,
            I => \N__54054\
        );

    \I__13151\ : InMux
    port map (
            O => \N__54172\,
            I => \N__54054\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__54155\,
            I => \N__54047\
        );

    \I__13149\ : Span4Mux_v
    port map (
            O => \N__54152\,
            I => \N__54047\
        );

    \I__13148\ : Span4Mux_v
    port map (
            O => \N__54141\,
            I => \N__54047\
        );

    \I__13147\ : Span4Mux_h
    port map (
            O => \N__54136\,
            I => \N__54042\
        );

    \I__13146\ : Span4Mux_v
    port map (
            O => \N__54129\,
            I => \N__54042\
        );

    \I__13145\ : Span12Mux_h
    port map (
            O => \N__54126\,
            I => \N__54037\
        );

    \I__13144\ : Span12Mux_v
    port map (
            O => \N__54115\,
            I => \N__54037\
        );

    \I__13143\ : Span4Mux_h
    port map (
            O => \N__54112\,
            I => \N__54032\
        );

    \I__13142\ : Span4Mux_h
    port map (
            O => \N__54103\,
            I => \N__54032\
        );

    \I__13141\ : LocalMux
    port map (
            O => \N__54086\,
            I => comm_state_1
        );

    \I__13140\ : LocalMux
    port map (
            O => \N__54081\,
            I => comm_state_1
        );

    \I__13139\ : Odrv12
    port map (
            O => \N__54078\,
            I => comm_state_1
        );

    \I__13138\ : Odrv12
    port map (
            O => \N__54075\,
            I => comm_state_1
        );

    \I__13137\ : LocalMux
    port map (
            O => \N__54068\,
            I => comm_state_1
        );

    \I__13136\ : LocalMux
    port map (
            O => \N__54063\,
            I => comm_state_1
        );

    \I__13135\ : LocalMux
    port map (
            O => \N__54054\,
            I => comm_state_1
        );

    \I__13134\ : Odrv4
    port map (
            O => \N__54047\,
            I => comm_state_1
        );

    \I__13133\ : Odrv4
    port map (
            O => \N__54042\,
            I => comm_state_1
        );

    \I__13132\ : Odrv12
    port map (
            O => \N__54037\,
            I => comm_state_1
        );

    \I__13131\ : Odrv4
    port map (
            O => \N__54032\,
            I => comm_state_1
        );

    \I__13130\ : InMux
    port map (
            O => \N__54009\,
            I => \N__53998\
        );

    \I__13129\ : InMux
    port map (
            O => \N__54008\,
            I => \N__53994\
        );

    \I__13128\ : InMux
    port map (
            O => \N__54007\,
            I => \N__53989\
        );

    \I__13127\ : InMux
    port map (
            O => \N__54006\,
            I => \N__53989\
        );

    \I__13126\ : CascadeMux
    port map (
            O => \N__54005\,
            I => \N__53983\
        );

    \I__13125\ : InMux
    port map (
            O => \N__54004\,
            I => \N__53970\
        );

    \I__13124\ : InMux
    port map (
            O => \N__54003\,
            I => \N__53970\
        );

    \I__13123\ : InMux
    port map (
            O => \N__54002\,
            I => \N__53970\
        );

    \I__13122\ : InMux
    port map (
            O => \N__54001\,
            I => \N__53966\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__53998\,
            I => \N__53959\
        );

    \I__13120\ : InMux
    port map (
            O => \N__53997\,
            I => \N__53956\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__53994\,
            I => \N__53951\
        );

    \I__13118\ : LocalMux
    port map (
            O => \N__53989\,
            I => \N__53951\
        );

    \I__13117\ : InMux
    port map (
            O => \N__53988\,
            I => \N__53948\
        );

    \I__13116\ : InMux
    port map (
            O => \N__53987\,
            I => \N__53943\
        );

    \I__13115\ : CascadeMux
    port map (
            O => \N__53986\,
            I => \N__53940\
        );

    \I__13114\ : InMux
    port map (
            O => \N__53983\,
            I => \N__53931\
        );

    \I__13113\ : InMux
    port map (
            O => \N__53982\,
            I => \N__53931\
        );

    \I__13112\ : InMux
    port map (
            O => \N__53981\,
            I => \N__53931\
        );

    \I__13111\ : InMux
    port map (
            O => \N__53980\,
            I => \N__53931\
        );

    \I__13110\ : InMux
    port map (
            O => \N__53979\,
            I => \N__53924\
        );

    \I__13109\ : InMux
    port map (
            O => \N__53978\,
            I => \N__53924\
        );

    \I__13108\ : InMux
    port map (
            O => \N__53977\,
            I => \N__53924\
        );

    \I__13107\ : LocalMux
    port map (
            O => \N__53970\,
            I => \N__53916\
        );

    \I__13106\ : InMux
    port map (
            O => \N__53969\,
            I => \N__53913\
        );

    \I__13105\ : LocalMux
    port map (
            O => \N__53966\,
            I => \N__53910\
        );

    \I__13104\ : InMux
    port map (
            O => \N__53965\,
            I => \N__53905\
        );

    \I__13103\ : InMux
    port map (
            O => \N__53964\,
            I => \N__53905\
        );

    \I__13102\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53900\
        );

    \I__13101\ : InMux
    port map (
            O => \N__53962\,
            I => \N__53900\
        );

    \I__13100\ : Span4Mux_v
    port map (
            O => \N__53959\,
            I => \N__53897\
        );

    \I__13099\ : LocalMux
    port map (
            O => \N__53956\,
            I => \N__53894\
        );

    \I__13098\ : Span4Mux_h
    port map (
            O => \N__53951\,
            I => \N__53889\
        );

    \I__13097\ : LocalMux
    port map (
            O => \N__53948\,
            I => \N__53889\
        );

    \I__13096\ : InMux
    port map (
            O => \N__53947\,
            I => \N__53886\
        );

    \I__13095\ : InMux
    port map (
            O => \N__53946\,
            I => \N__53883\
        );

    \I__13094\ : LocalMux
    port map (
            O => \N__53943\,
            I => \N__53880\
        );

    \I__13093\ : InMux
    port map (
            O => \N__53940\,
            I => \N__53877\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__53931\,
            I => \N__53874\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__53924\,
            I => \N__53865\
        );

    \I__13090\ : InMux
    port map (
            O => \N__53923\,
            I => \N__53860\
        );

    \I__13089\ : InMux
    port map (
            O => \N__53922\,
            I => \N__53860\
        );

    \I__13088\ : InMux
    port map (
            O => \N__53921\,
            I => \N__53853\
        );

    \I__13087\ : InMux
    port map (
            O => \N__53920\,
            I => \N__53853\
        );

    \I__13086\ : InMux
    port map (
            O => \N__53919\,
            I => \N__53853\
        );

    \I__13085\ : Span4Mux_v
    port map (
            O => \N__53916\,
            I => \N__53850\
        );

    \I__13084\ : LocalMux
    port map (
            O => \N__53913\,
            I => \N__53845\
        );

    \I__13083\ : Span4Mux_v
    port map (
            O => \N__53910\,
            I => \N__53845\
        );

    \I__13082\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53838\
        );

    \I__13081\ : LocalMux
    port map (
            O => \N__53900\,
            I => \N__53838\
        );

    \I__13080\ : Span4Mux_h
    port map (
            O => \N__53897\,
            I => \N__53838\
        );

    \I__13079\ : Span4Mux_v
    port map (
            O => \N__53894\,
            I => \N__53833\
        );

    \I__13078\ : Span4Mux_v
    port map (
            O => \N__53889\,
            I => \N__53833\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__53886\,
            I => \N__53830\
        );

    \I__13076\ : LocalMux
    port map (
            O => \N__53883\,
            I => \N__53823\
        );

    \I__13075\ : Span4Mux_v
    port map (
            O => \N__53880\,
            I => \N__53823\
        );

    \I__13074\ : LocalMux
    port map (
            O => \N__53877\,
            I => \N__53823\
        );

    \I__13073\ : Span4Mux_v
    port map (
            O => \N__53874\,
            I => \N__53820\
        );

    \I__13072\ : InMux
    port map (
            O => \N__53873\,
            I => \N__53811\
        );

    \I__13071\ : InMux
    port map (
            O => \N__53872\,
            I => \N__53811\
        );

    \I__13070\ : InMux
    port map (
            O => \N__53871\,
            I => \N__53811\
        );

    \I__13069\ : InMux
    port map (
            O => \N__53870\,
            I => \N__53811\
        );

    \I__13068\ : InMux
    port map (
            O => \N__53869\,
            I => \N__53806\
        );

    \I__13067\ : InMux
    port map (
            O => \N__53868\,
            I => \N__53806\
        );

    \I__13066\ : Span4Mux_v
    port map (
            O => \N__53865\,
            I => \N__53793\
        );

    \I__13065\ : LocalMux
    port map (
            O => \N__53860\,
            I => \N__53793\
        );

    \I__13064\ : LocalMux
    port map (
            O => \N__53853\,
            I => \N__53793\
        );

    \I__13063\ : Span4Mux_v
    port map (
            O => \N__53850\,
            I => \N__53793\
        );

    \I__13062\ : Span4Mux_h
    port map (
            O => \N__53845\,
            I => \N__53793\
        );

    \I__13061\ : Span4Mux_v
    port map (
            O => \N__53838\,
            I => \N__53793\
        );

    \I__13060\ : Span4Mux_h
    port map (
            O => \N__53833\,
            I => \N__53790\
        );

    \I__13059\ : Odrv12
    port map (
            O => \N__53830\,
            I => comm_state_0
        );

    \I__13058\ : Odrv4
    port map (
            O => \N__53823\,
            I => comm_state_0
        );

    \I__13057\ : Odrv4
    port map (
            O => \N__53820\,
            I => comm_state_0
        );

    \I__13056\ : LocalMux
    port map (
            O => \N__53811\,
            I => comm_state_0
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__53806\,
            I => comm_state_0
        );

    \I__13054\ : Odrv4
    port map (
            O => \N__53793\,
            I => comm_state_0
        );

    \I__13053\ : Odrv4
    port map (
            O => \N__53790\,
            I => comm_state_0
        );

    \I__13052\ : InMux
    port map (
            O => \N__53775\,
            I => \N__53772\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__53772\,
            I => \N__53769\
        );

    \I__13050\ : Span4Mux_v
    port map (
            O => \N__53769\,
            I => \N__53766\
        );

    \I__13049\ : Span4Mux_h
    port map (
            O => \N__53766\,
            I => \N__53763\
        );

    \I__13048\ : Odrv4
    port map (
            O => \N__53763\,
            I => n10804
        );

    \I__13047\ : InMux
    port map (
            O => \N__53760\,
            I => \N__53757\
        );

    \I__13046\ : LocalMux
    port map (
            O => \N__53757\,
            I => \N__53753\
        );

    \I__13045\ : InMux
    port map (
            O => \N__53756\,
            I => \N__53750\
        );

    \I__13044\ : Span4Mux_h
    port map (
            O => \N__53753\,
            I => \N__53747\
        );

    \I__13043\ : LocalMux
    port map (
            O => \N__53750\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__13042\ : Odrv4
    port map (
            O => \N__53747\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__13041\ : CascadeMux
    port map (
            O => \N__53742\,
            I => \N__53738\
        );

    \I__13040\ : InMux
    port map (
            O => \N__53741\,
            I => \N__53735\
        );

    \I__13039\ : InMux
    port map (
            O => \N__53738\,
            I => \N__53732\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__53735\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__13037\ : LocalMux
    port map (
            O => \N__53732\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__13036\ : CascadeMux
    port map (
            O => \N__53727\,
            I => \N__53723\
        );

    \I__13035\ : InMux
    port map (
            O => \N__53726\,
            I => \N__53720\
        );

    \I__13034\ : InMux
    port map (
            O => \N__53723\,
            I => \N__53717\
        );

    \I__13033\ : LocalMux
    port map (
            O => \N__53720\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__13032\ : LocalMux
    port map (
            O => \N__53717\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__13031\ : InMux
    port map (
            O => \N__53712\,
            I => \N__53708\
        );

    \I__13030\ : InMux
    port map (
            O => \N__53711\,
            I => \N__53705\
        );

    \I__13029\ : LocalMux
    port map (
            O => \N__53708\,
            I => \N__53702\
        );

    \I__13028\ : LocalMux
    port map (
            O => \N__53705\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__13027\ : Odrv4
    port map (
            O => \N__53702\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__13026\ : CascadeMux
    port map (
            O => \N__53697\,
            I => \ADC_VDC.genclk.n27_cascade_\
        );

    \I__13025\ : CascadeMux
    port map (
            O => \N__53694\,
            I => \ADC_VDC.genclk.n21598_cascade_\
        );

    \I__13024\ : CEMux
    port map (
            O => \N__53691\,
            I => \N__53688\
        );

    \I__13023\ : LocalMux
    port map (
            O => \N__53688\,
            I => \ADC_VDC.genclk.n6\
        );

    \I__13022\ : InMux
    port map (
            O => \N__53685\,
            I => \N__53682\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__53682\,
            I => \N__53679\
        );

    \I__13020\ : Span4Mux_h
    port map (
            O => \N__53679\,
            I => \N__53676\
        );

    \I__13019\ : Span4Mux_h
    port map (
            O => \N__53676\,
            I => \N__53671\
        );

    \I__13018\ : InMux
    port map (
            O => \N__53675\,
            I => \N__53666\
        );

    \I__13017\ : InMux
    port map (
            O => \N__53674\,
            I => \N__53666\
        );

    \I__13016\ : Span4Mux_v
    port map (
            O => \N__53671\,
            I => \N__53663\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__53666\,
            I => \N__53660\
        );

    \I__13014\ : Odrv4
    port map (
            O => \N__53663\,
            I => comm_tx_buf_5
        );

    \I__13013\ : Odrv4
    port map (
            O => \N__53660\,
            I => comm_tx_buf_5
        );

    \I__13012\ : SRMux
    port map (
            O => \N__53655\,
            I => \N__53652\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__53652\,
            I => \comm_spi.data_tx_7__N_808\
        );

    \I__13010\ : InMux
    port map (
            O => \N__53649\,
            I => \N__53646\
        );

    \I__13009\ : LocalMux
    port map (
            O => \N__53646\,
            I => \N__53641\
        );

    \I__13008\ : InMux
    port map (
            O => \N__53645\,
            I => \N__53637\
        );

    \I__13007\ : InMux
    port map (
            O => \N__53644\,
            I => \N__53633\
        );

    \I__13006\ : Span4Mux_h
    port map (
            O => \N__53641\,
            I => \N__53630\
        );

    \I__13005\ : InMux
    port map (
            O => \N__53640\,
            I => \N__53627\
        );

    \I__13004\ : LocalMux
    port map (
            O => \N__53637\,
            I => \N__53624\
        );

    \I__13003\ : InMux
    port map (
            O => \N__53636\,
            I => \N__53621\
        );

    \I__13002\ : LocalMux
    port map (
            O => \N__53633\,
            I => \N__53612\
        );

    \I__13001\ : Span4Mux_h
    port map (
            O => \N__53630\,
            I => \N__53612\
        );

    \I__13000\ : LocalMux
    port map (
            O => \N__53627\,
            I => \N__53612\
        );

    \I__12999\ : Span4Mux_v
    port map (
            O => \N__53624\,
            I => \N__53607\
        );

    \I__12998\ : LocalMux
    port map (
            O => \N__53621\,
            I => \N__53607\
        );

    \I__12997\ : InMux
    port map (
            O => \N__53620\,
            I => \N__53604\
        );

    \I__12996\ : InMux
    port map (
            O => \N__53619\,
            I => \N__53601\
        );

    \I__12995\ : Span4Mux_v
    port map (
            O => \N__53612\,
            I => \N__53597\
        );

    \I__12994\ : Span4Mux_v
    port map (
            O => \N__53607\,
            I => \N__53594\
        );

    \I__12993\ : LocalMux
    port map (
            O => \N__53604\,
            I => \N__53591\
        );

    \I__12992\ : LocalMux
    port map (
            O => \N__53601\,
            I => \N__53588\
        );

    \I__12991\ : InMux
    port map (
            O => \N__53600\,
            I => \N__53585\
        );

    \I__12990\ : Sp12to4
    port map (
            O => \N__53597\,
            I => \N__53581\
        );

    \I__12989\ : Span4Mux_h
    port map (
            O => \N__53594\,
            I => \N__53578\
        );

    \I__12988\ : Span4Mux_h
    port map (
            O => \N__53591\,
            I => \N__53573\
        );

    \I__12987\ : Span4Mux_h
    port map (
            O => \N__53588\,
            I => \N__53573\
        );

    \I__12986\ : LocalMux
    port map (
            O => \N__53585\,
            I => \N__53570\
        );

    \I__12985\ : InMux
    port map (
            O => \N__53584\,
            I => \N__53567\
        );

    \I__12984\ : Odrv12
    port map (
            O => \N__53581\,
            I => comm_rx_buf_4
        );

    \I__12983\ : Odrv4
    port map (
            O => \N__53578\,
            I => comm_rx_buf_4
        );

    \I__12982\ : Odrv4
    port map (
            O => \N__53573\,
            I => comm_rx_buf_4
        );

    \I__12981\ : Odrv4
    port map (
            O => \N__53570\,
            I => comm_rx_buf_4
        );

    \I__12980\ : LocalMux
    port map (
            O => \N__53567\,
            I => comm_rx_buf_4
        );

    \I__12979\ : InMux
    port map (
            O => \N__53556\,
            I => \N__53553\
        );

    \I__12978\ : LocalMux
    port map (
            O => \N__53553\,
            I => \N__53549\
        );

    \I__12977\ : InMux
    port map (
            O => \N__53552\,
            I => \N__53546\
        );

    \I__12976\ : Span4Mux_h
    port map (
            O => \N__53549\,
            I => \N__53543\
        );

    \I__12975\ : LocalMux
    port map (
            O => \N__53546\,
            I => comm_buf_6_4
        );

    \I__12974\ : Odrv4
    port map (
            O => \N__53543\,
            I => comm_buf_6_4
        );

    \I__12973\ : InMux
    port map (
            O => \N__53538\,
            I => \N__53535\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__53535\,
            I => \N__53532\
        );

    \I__12971\ : Odrv4
    port map (
            O => \N__53532\,
            I => comm_buf_3_1
        );

    \I__12970\ : InMux
    port map (
            O => \N__53529\,
            I => \N__53526\
        );

    \I__12969\ : LocalMux
    port map (
            O => \N__53526\,
            I => \N__53523\
        );

    \I__12968\ : Span4Mux_h
    port map (
            O => \N__53523\,
            I => \N__53520\
        );

    \I__12967\ : Odrv4
    port map (
            O => \N__53520\,
            I => comm_buf_2_1
        );

    \I__12966\ : InMux
    port map (
            O => \N__53517\,
            I => \N__53514\
        );

    \I__12965\ : LocalMux
    port map (
            O => \N__53514\,
            I => n2_adj_1587
        );

    \I__12964\ : InMux
    port map (
            O => \N__53511\,
            I => \N__53507\
        );

    \I__12963\ : InMux
    port map (
            O => \N__53510\,
            I => \N__53504\
        );

    \I__12962\ : LocalMux
    port map (
            O => \N__53507\,
            I => \N__53500\
        );

    \I__12961\ : LocalMux
    port map (
            O => \N__53504\,
            I => \N__53496\
        );

    \I__12960\ : InMux
    port map (
            O => \N__53503\,
            I => \N__53493\
        );

    \I__12959\ : Span4Mux_v
    port map (
            O => \N__53500\,
            I => \N__53490\
        );

    \I__12958\ : InMux
    port map (
            O => \N__53499\,
            I => \N__53487\
        );

    \I__12957\ : Span4Mux_h
    port map (
            O => \N__53496\,
            I => \N__53482\
        );

    \I__12956\ : LocalMux
    port map (
            O => \N__53493\,
            I => \N__53482\
        );

    \I__12955\ : Sp12to4
    port map (
            O => \N__53490\,
            I => \N__53477\
        );

    \I__12954\ : LocalMux
    port map (
            O => \N__53487\,
            I => \N__53477\
        );

    \I__12953\ : Span4Mux_h
    port map (
            O => \N__53482\,
            I => \N__53474\
        );

    \I__12952\ : Span12Mux_s11_v
    port map (
            O => \N__53477\,
            I => \N__53471\
        );

    \I__12951\ : Odrv4
    port map (
            O => \N__53474\,
            I => comm_buf_1_1
        );

    \I__12950\ : Odrv12
    port map (
            O => \N__53471\,
            I => comm_buf_1_1
        );

    \I__12949\ : CascadeMux
    port map (
            O => \N__53466\,
            I => \N__53463\
        );

    \I__12948\ : InMux
    port map (
            O => \N__53463\,
            I => \N__53459\
        );

    \I__12947\ : CascadeMux
    port map (
            O => \N__53462\,
            I => \N__53455\
        );

    \I__12946\ : LocalMux
    port map (
            O => \N__53459\,
            I => \N__53452\
        );

    \I__12945\ : CascadeMux
    port map (
            O => \N__53458\,
            I => \N__53449\
        );

    \I__12944\ : InMux
    port map (
            O => \N__53455\,
            I => \N__53445\
        );

    \I__12943\ : Span4Mux_h
    port map (
            O => \N__53452\,
            I => \N__53442\
        );

    \I__12942\ : InMux
    port map (
            O => \N__53449\,
            I => \N__53439\
        );

    \I__12941\ : InMux
    port map (
            O => \N__53448\,
            I => \N__53432\
        );

    \I__12940\ : LocalMux
    port map (
            O => \N__53445\,
            I => \N__53425\
        );

    \I__12939\ : Span4Mux_h
    port map (
            O => \N__53442\,
            I => \N__53425\
        );

    \I__12938\ : LocalMux
    port map (
            O => \N__53439\,
            I => \N__53425\
        );

    \I__12937\ : InMux
    port map (
            O => \N__53438\,
            I => \N__53418\
        );

    \I__12936\ : InMux
    port map (
            O => \N__53437\,
            I => \N__53418\
        );

    \I__12935\ : InMux
    port map (
            O => \N__53436\,
            I => \N__53415\
        );

    \I__12934\ : InMux
    port map (
            O => \N__53435\,
            I => \N__53412\
        );

    \I__12933\ : LocalMux
    port map (
            O => \N__53432\,
            I => \N__53407\
        );

    \I__12932\ : Span4Mux_v
    port map (
            O => \N__53425\,
            I => \N__53407\
        );

    \I__12931\ : InMux
    port map (
            O => \N__53424\,
            I => \N__53404\
        );

    \I__12930\ : InMux
    port map (
            O => \N__53423\,
            I => \N__53401\
        );

    \I__12929\ : LocalMux
    port map (
            O => \N__53418\,
            I => \N__53398\
        );

    \I__12928\ : LocalMux
    port map (
            O => \N__53415\,
            I => \N__53393\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__53412\,
            I => \N__53393\
        );

    \I__12926\ : Span4Mux_h
    port map (
            O => \N__53407\,
            I => \N__53390\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__53404\,
            I => \N__53387\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__53401\,
            I => \N__53384\
        );

    \I__12923\ : Span4Mux_h
    port map (
            O => \N__53398\,
            I => \N__53381\
        );

    \I__12922\ : Span4Mux_v
    port map (
            O => \N__53393\,
            I => \N__53378\
        );

    \I__12921\ : Span4Mux_h
    port map (
            O => \N__53390\,
            I => \N__53375\
        );

    \I__12920\ : Span4Mux_v
    port map (
            O => \N__53387\,
            I => \N__53370\
        );

    \I__12919\ : Span4Mux_v
    port map (
            O => \N__53384\,
            I => \N__53370\
        );

    \I__12918\ : Span4Mux_v
    port map (
            O => \N__53381\,
            I => \N__53367\
        );

    \I__12917\ : Odrv4
    port map (
            O => \N__53378\,
            I => comm_buf_0_1
        );

    \I__12916\ : Odrv4
    port map (
            O => \N__53375\,
            I => comm_buf_0_1
        );

    \I__12915\ : Odrv4
    port map (
            O => \N__53370\,
            I => comm_buf_0_1
        );

    \I__12914\ : Odrv4
    port map (
            O => \N__53367\,
            I => comm_buf_0_1
        );

    \I__12913\ : InMux
    port map (
            O => \N__53358\,
            I => \N__53355\
        );

    \I__12912\ : LocalMux
    port map (
            O => \N__53355\,
            I => \N__53352\
        );

    \I__12911\ : Odrv4
    port map (
            O => \N__53352\,
            I => n1_adj_1586
        );

    \I__12910\ : CascadeMux
    port map (
            O => \N__53349\,
            I => \N__53346\
        );

    \I__12909\ : InMux
    port map (
            O => \N__53346\,
            I => \N__53339\
        );

    \I__12908\ : CascadeMux
    port map (
            O => \N__53345\,
            I => \N__53336\
        );

    \I__12907\ : CascadeMux
    port map (
            O => \N__53344\,
            I => \N__53333\
        );

    \I__12906\ : InMux
    port map (
            O => \N__53343\,
            I => \N__53328\
        );

    \I__12905\ : InMux
    port map (
            O => \N__53342\,
            I => \N__53325\
        );

    \I__12904\ : LocalMux
    port map (
            O => \N__53339\,
            I => \N__53322\
        );

    \I__12903\ : InMux
    port map (
            O => \N__53336\,
            I => \N__53319\
        );

    \I__12902\ : InMux
    port map (
            O => \N__53333\,
            I => \N__53316\
        );

    \I__12901\ : InMux
    port map (
            O => \N__53332\,
            I => \N__53313\
        );

    \I__12900\ : InMux
    port map (
            O => \N__53331\,
            I => \N__53310\
        );

    \I__12899\ : LocalMux
    port map (
            O => \N__53328\,
            I => \N__53305\
        );

    \I__12898\ : LocalMux
    port map (
            O => \N__53325\,
            I => \N__53305\
        );

    \I__12897\ : Span4Mux_h
    port map (
            O => \N__53322\,
            I => \N__53298\
        );

    \I__12896\ : LocalMux
    port map (
            O => \N__53319\,
            I => \N__53298\
        );

    \I__12895\ : LocalMux
    port map (
            O => \N__53316\,
            I => \N__53298\
        );

    \I__12894\ : LocalMux
    port map (
            O => \N__53313\,
            I => \N__53293\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__53310\,
            I => \N__53293\
        );

    \I__12892\ : Span4Mux_v
    port map (
            O => \N__53305\,
            I => \N__53288\
        );

    \I__12891\ : Span4Mux_v
    port map (
            O => \N__53298\,
            I => \N__53283\
        );

    \I__12890\ : Span4Mux_v
    port map (
            O => \N__53293\,
            I => \N__53283\
        );

    \I__12889\ : InMux
    port map (
            O => \N__53292\,
            I => \N__53280\
        );

    \I__12888\ : InMux
    port map (
            O => \N__53291\,
            I => \N__53277\
        );

    \I__12887\ : Odrv4
    port map (
            O => \N__53288\,
            I => comm_rx_buf_5
        );

    \I__12886\ : Odrv4
    port map (
            O => \N__53283\,
            I => comm_rx_buf_5
        );

    \I__12885\ : LocalMux
    port map (
            O => \N__53280\,
            I => comm_rx_buf_5
        );

    \I__12884\ : LocalMux
    port map (
            O => \N__53277\,
            I => comm_rx_buf_5
        );

    \I__12883\ : InMux
    port map (
            O => \N__53268\,
            I => \N__53264\
        );

    \I__12882\ : InMux
    port map (
            O => \N__53267\,
            I => \N__53261\
        );

    \I__12881\ : LocalMux
    port map (
            O => \N__53264\,
            I => comm_buf_6_5
        );

    \I__12880\ : LocalMux
    port map (
            O => \N__53261\,
            I => comm_buf_6_5
        );

    \I__12879\ : InMux
    port map (
            O => \N__53256\,
            I => \N__53253\
        );

    \I__12878\ : LocalMux
    port map (
            O => \N__53253\,
            I => \N__53250\
        );

    \I__12877\ : Span4Mux_h
    port map (
            O => \N__53250\,
            I => \N__53247\
        );

    \I__12876\ : Odrv4
    port map (
            O => \N__53247\,
            I => buf_data_iac_14
        );

    \I__12875\ : InMux
    port map (
            O => \N__53244\,
            I => \N__53241\
        );

    \I__12874\ : LocalMux
    port map (
            O => \N__53241\,
            I => \N__53238\
        );

    \I__12873\ : Odrv4
    port map (
            O => \N__53238\,
            I => n21547
        );

    \I__12872\ : CascadeMux
    port map (
            O => \N__53235\,
            I => \N__53231\
        );

    \I__12871\ : CascadeMux
    port map (
            O => \N__53234\,
            I => \N__53228\
        );

    \I__12870\ : InMux
    port map (
            O => \N__53231\,
            I => \N__53222\
        );

    \I__12869\ : InMux
    port map (
            O => \N__53228\,
            I => \N__53219\
        );

    \I__12868\ : InMux
    port map (
            O => \N__53227\,
            I => \N__53214\
        );

    \I__12867\ : InMux
    port map (
            O => \N__53226\,
            I => \N__53211\
        );

    \I__12866\ : InMux
    port map (
            O => \N__53225\,
            I => \N__53208\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__53222\,
            I => \N__53205\
        );

    \I__12864\ : LocalMux
    port map (
            O => \N__53219\,
            I => \N__53202\
        );

    \I__12863\ : InMux
    port map (
            O => \N__53218\,
            I => \N__53199\
        );

    \I__12862\ : InMux
    port map (
            O => \N__53217\,
            I => \N__53196\
        );

    \I__12861\ : LocalMux
    port map (
            O => \N__53214\,
            I => \N__53192\
        );

    \I__12860\ : LocalMux
    port map (
            O => \N__53211\,
            I => \N__53189\
        );

    \I__12859\ : LocalMux
    port map (
            O => \N__53208\,
            I => \N__53184\
        );

    \I__12858\ : Span4Mux_h
    port map (
            O => \N__53205\,
            I => \N__53184\
        );

    \I__12857\ : Span4Mux_v
    port map (
            O => \N__53202\,
            I => \N__53177\
        );

    \I__12856\ : LocalMux
    port map (
            O => \N__53199\,
            I => \N__53177\
        );

    \I__12855\ : LocalMux
    port map (
            O => \N__53196\,
            I => \N__53177\
        );

    \I__12854\ : InMux
    port map (
            O => \N__53195\,
            I => \N__53174\
        );

    \I__12853\ : Span4Mux_v
    port map (
            O => \N__53192\,
            I => \N__53171\
        );

    \I__12852\ : Span4Mux_h
    port map (
            O => \N__53189\,
            I => \N__53166\
        );

    \I__12851\ : Span4Mux_h
    port map (
            O => \N__53184\,
            I => \N__53166\
        );

    \I__12850\ : Span4Mux_h
    port map (
            O => \N__53177\,
            I => \N__53161\
        );

    \I__12849\ : LocalMux
    port map (
            O => \N__53174\,
            I => \N__53161\
        );

    \I__12848\ : Sp12to4
    port map (
            O => \N__53171\,
            I => \N__53157\
        );

    \I__12847\ : Sp12to4
    port map (
            O => \N__53166\,
            I => \N__53152\
        );

    \I__12846\ : Sp12to4
    port map (
            O => \N__53161\,
            I => \N__53152\
        );

    \I__12845\ : InMux
    port map (
            O => \N__53160\,
            I => \N__53149\
        );

    \I__12844\ : Odrv12
    port map (
            O => \N__53157\,
            I => comm_rx_buf_6
        );

    \I__12843\ : Odrv12
    port map (
            O => \N__53152\,
            I => comm_rx_buf_6
        );

    \I__12842\ : LocalMux
    port map (
            O => \N__53149\,
            I => comm_rx_buf_6
        );

    \I__12841\ : InMux
    port map (
            O => \N__53142\,
            I => \N__53138\
        );

    \I__12840\ : InMux
    port map (
            O => \N__53141\,
            I => \N__53135\
        );

    \I__12839\ : LocalMux
    port map (
            O => \N__53138\,
            I => \N__53132\
        );

    \I__12838\ : LocalMux
    port map (
            O => \N__53135\,
            I => \N__53123\
        );

    \I__12837\ : Span4Mux_h
    port map (
            O => \N__53132\,
            I => \N__53120\
        );

    \I__12836\ : InMux
    port map (
            O => \N__53131\,
            I => \N__53117\
        );

    \I__12835\ : InMux
    port map (
            O => \N__53130\,
            I => \N__53114\
        );

    \I__12834\ : InMux
    port map (
            O => \N__53129\,
            I => \N__53109\
        );

    \I__12833\ : InMux
    port map (
            O => \N__53128\,
            I => \N__53109\
        );

    \I__12832\ : InMux
    port map (
            O => \N__53127\,
            I => \N__53106\
        );

    \I__12831\ : InMux
    port map (
            O => \N__53126\,
            I => \N__53103\
        );

    \I__12830\ : Odrv12
    port map (
            O => \N__53123\,
            I => n12477
        );

    \I__12829\ : Odrv4
    port map (
            O => \N__53120\,
            I => n12477
        );

    \I__12828\ : LocalMux
    port map (
            O => \N__53117\,
            I => n12477
        );

    \I__12827\ : LocalMux
    port map (
            O => \N__53114\,
            I => n12477
        );

    \I__12826\ : LocalMux
    port map (
            O => \N__53109\,
            I => n12477
        );

    \I__12825\ : LocalMux
    port map (
            O => \N__53106\,
            I => n12477
        );

    \I__12824\ : LocalMux
    port map (
            O => \N__53103\,
            I => n12477
        );

    \I__12823\ : CascadeMux
    port map (
            O => \N__53088\,
            I => \N__53084\
        );

    \I__12822\ : InMux
    port map (
            O => \N__53087\,
            I => \N__53081\
        );

    \I__12821\ : InMux
    port map (
            O => \N__53084\,
            I => \N__53078\
        );

    \I__12820\ : LocalMux
    port map (
            O => \N__53081\,
            I => comm_buf_6_6
        );

    \I__12819\ : LocalMux
    port map (
            O => \N__53078\,
            I => comm_buf_6_6
        );

    \I__12818\ : InMux
    port map (
            O => \N__53073\,
            I => \N__53058\
        );

    \I__12817\ : InMux
    port map (
            O => \N__53072\,
            I => \N__53053\
        );

    \I__12816\ : InMux
    port map (
            O => \N__53071\,
            I => \N__53053\
        );

    \I__12815\ : CascadeMux
    port map (
            O => \N__53070\,
            I => \N__53043\
        );

    \I__12814\ : InMux
    port map (
            O => \N__53069\,
            I => \N__53037\
        );

    \I__12813\ : InMux
    port map (
            O => \N__53068\,
            I => \N__53037\
        );

    \I__12812\ : InMux
    port map (
            O => \N__53067\,
            I => \N__53034\
        );

    \I__12811\ : InMux
    port map (
            O => \N__53066\,
            I => \N__53025\
        );

    \I__12810\ : InMux
    port map (
            O => \N__53065\,
            I => \N__53014\
        );

    \I__12809\ : InMux
    port map (
            O => \N__53064\,
            I => \N__53014\
        );

    \I__12808\ : InMux
    port map (
            O => \N__53063\,
            I => \N__53014\
        );

    \I__12807\ : InMux
    port map (
            O => \N__53062\,
            I => \N__53014\
        );

    \I__12806\ : InMux
    port map (
            O => \N__53061\,
            I => \N__53014\
        );

    \I__12805\ : LocalMux
    port map (
            O => \N__53058\,
            I => \N__53009\
        );

    \I__12804\ : LocalMux
    port map (
            O => \N__53053\,
            I => \N__53009\
        );

    \I__12803\ : InMux
    port map (
            O => \N__53052\,
            I => \N__53002\
        );

    \I__12802\ : InMux
    port map (
            O => \N__53051\,
            I => \N__53002\
        );

    \I__12801\ : InMux
    port map (
            O => \N__53050\,
            I => \N__53002\
        );

    \I__12800\ : InMux
    port map (
            O => \N__53049\,
            I => \N__52993\
        );

    \I__12799\ : InMux
    port map (
            O => \N__53048\,
            I => \N__52993\
        );

    \I__12798\ : InMux
    port map (
            O => \N__53047\,
            I => \N__52993\
        );

    \I__12797\ : InMux
    port map (
            O => \N__53046\,
            I => \N__52993\
        );

    \I__12796\ : InMux
    port map (
            O => \N__53043\,
            I => \N__52983\
        );

    \I__12795\ : InMux
    port map (
            O => \N__53042\,
            I => \N__52980\
        );

    \I__12794\ : LocalMux
    port map (
            O => \N__53037\,
            I => \N__52975\
        );

    \I__12793\ : LocalMux
    port map (
            O => \N__53034\,
            I => \N__52975\
        );

    \I__12792\ : InMux
    port map (
            O => \N__53033\,
            I => \N__52966\
        );

    \I__12791\ : InMux
    port map (
            O => \N__53032\,
            I => \N__52966\
        );

    \I__12790\ : InMux
    port map (
            O => \N__53031\,
            I => \N__52966\
        );

    \I__12789\ : InMux
    port map (
            O => \N__53030\,
            I => \N__52966\
        );

    \I__12788\ : InMux
    port map (
            O => \N__53029\,
            I => \N__52963\
        );

    \I__12787\ : InMux
    port map (
            O => \N__53028\,
            I => \N__52960\
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__53025\,
            I => \N__52951\
        );

    \I__12785\ : LocalMux
    port map (
            O => \N__53014\,
            I => \N__52951\
        );

    \I__12784\ : Span4Mux_v
    port map (
            O => \N__53009\,
            I => \N__52951\
        );

    \I__12783\ : LocalMux
    port map (
            O => \N__53002\,
            I => \N__52951\
        );

    \I__12782\ : LocalMux
    port map (
            O => \N__52993\,
            I => \N__52948\
        );

    \I__12781\ : InMux
    port map (
            O => \N__52992\,
            I => \N__52939\
        );

    \I__12780\ : InMux
    port map (
            O => \N__52991\,
            I => \N__52939\
        );

    \I__12779\ : InMux
    port map (
            O => \N__52990\,
            I => \N__52939\
        );

    \I__12778\ : InMux
    port map (
            O => \N__52989\,
            I => \N__52939\
        );

    \I__12777\ : InMux
    port map (
            O => \N__52988\,
            I => \N__52933\
        );

    \I__12776\ : InMux
    port map (
            O => \N__52987\,
            I => \N__52933\
        );

    \I__12775\ : InMux
    port map (
            O => \N__52986\,
            I => \N__52930\
        );

    \I__12774\ : LocalMux
    port map (
            O => \N__52983\,
            I => \N__52927\
        );

    \I__12773\ : LocalMux
    port map (
            O => \N__52980\,
            I => \N__52920\
        );

    \I__12772\ : Span4Mux_v
    port map (
            O => \N__52975\,
            I => \N__52920\
        );

    \I__12771\ : LocalMux
    port map (
            O => \N__52966\,
            I => \N__52920\
        );

    \I__12770\ : LocalMux
    port map (
            O => \N__52963\,
            I => \N__52915\
        );

    \I__12769\ : LocalMux
    port map (
            O => \N__52960\,
            I => \N__52915\
        );

    \I__12768\ : Span4Mux_v
    port map (
            O => \N__52951\,
            I => \N__52908\
        );

    \I__12767\ : Span4Mux_h
    port map (
            O => \N__52948\,
            I => \N__52908\
        );

    \I__12766\ : LocalMux
    port map (
            O => \N__52939\,
            I => \N__52908\
        );

    \I__12765\ : InMux
    port map (
            O => \N__52938\,
            I => \N__52905\
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__52933\,
            I => comm_index_0
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__52930\,
            I => comm_index_0
        );

    \I__12762\ : Odrv12
    port map (
            O => \N__52927\,
            I => comm_index_0
        );

    \I__12761\ : Odrv4
    port map (
            O => \N__52920\,
            I => comm_index_0
        );

    \I__12760\ : Odrv12
    port map (
            O => \N__52915\,
            I => comm_index_0
        );

    \I__12759\ : Odrv4
    port map (
            O => \N__52908\,
            I => comm_index_0
        );

    \I__12758\ : LocalMux
    port map (
            O => \N__52905\,
            I => comm_index_0
        );

    \I__12757\ : InMux
    port map (
            O => \N__52890\,
            I => \N__52887\
        );

    \I__12756\ : LocalMux
    port map (
            O => \N__52887\,
            I => n8_adj_1456
        );

    \I__12755\ : InMux
    port map (
            O => \N__52884\,
            I => \N__52872\
        );

    \I__12754\ : InMux
    port map (
            O => \N__52883\,
            I => \N__52872\
        );

    \I__12753\ : InMux
    port map (
            O => \N__52882\,
            I => \N__52872\
        );

    \I__12752\ : InMux
    port map (
            O => \N__52881\,
            I => \N__52869\
        );

    \I__12751\ : InMux
    port map (
            O => \N__52880\,
            I => \N__52864\
        );

    \I__12750\ : InMux
    port map (
            O => \N__52879\,
            I => \N__52864\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__52872\,
            I => \N__52852\
        );

    \I__12748\ : LocalMux
    port map (
            O => \N__52869\,
            I => \N__52849\
        );

    \I__12747\ : LocalMux
    port map (
            O => \N__52864\,
            I => \N__52846\
        );

    \I__12746\ : InMux
    port map (
            O => \N__52863\,
            I => \N__52839\
        );

    \I__12745\ : InMux
    port map (
            O => \N__52862\,
            I => \N__52839\
        );

    \I__12744\ : InMux
    port map (
            O => \N__52861\,
            I => \N__52839\
        );

    \I__12743\ : InMux
    port map (
            O => \N__52860\,
            I => \N__52828\
        );

    \I__12742\ : InMux
    port map (
            O => \N__52859\,
            I => \N__52828\
        );

    \I__12741\ : InMux
    port map (
            O => \N__52858\,
            I => \N__52828\
        );

    \I__12740\ : InMux
    port map (
            O => \N__52857\,
            I => \N__52828\
        );

    \I__12739\ : InMux
    port map (
            O => \N__52856\,
            I => \N__52828\
        );

    \I__12738\ : CascadeMux
    port map (
            O => \N__52855\,
            I => \N__52825\
        );

    \I__12737\ : Span4Mux_v
    port map (
            O => \N__52852\,
            I => \N__52820\
        );

    \I__12736\ : Span4Mux_v
    port map (
            O => \N__52849\,
            I => \N__52820\
        );

    \I__12735\ : Span4Mux_v
    port map (
            O => \N__52846\,
            I => \N__52813\
        );

    \I__12734\ : LocalMux
    port map (
            O => \N__52839\,
            I => \N__52813\
        );

    \I__12733\ : LocalMux
    port map (
            O => \N__52828\,
            I => \N__52813\
        );

    \I__12732\ : InMux
    port map (
            O => \N__52825\,
            I => \N__52810\
        );

    \I__12731\ : Odrv4
    port map (
            O => \N__52820\,
            I => comm_data_vld
        );

    \I__12730\ : Odrv4
    port map (
            O => \N__52813\,
            I => comm_data_vld
        );

    \I__12729\ : LocalMux
    port map (
            O => \N__52810\,
            I => comm_data_vld
        );

    \I__12728\ : CascadeMux
    port map (
            O => \N__52803\,
            I => \N__52800\
        );

    \I__12727\ : InMux
    port map (
            O => \N__52800\,
            I => \N__52784\
        );

    \I__12726\ : InMux
    port map (
            O => \N__52799\,
            I => \N__52784\
        );

    \I__12725\ : InMux
    port map (
            O => \N__52798\,
            I => \N__52784\
        );

    \I__12724\ : InMux
    port map (
            O => \N__52797\,
            I => \N__52784\
        );

    \I__12723\ : CascadeMux
    port map (
            O => \N__52796\,
            I => \N__52778\
        );

    \I__12722\ : CascadeMux
    port map (
            O => \N__52795\,
            I => \N__52775\
        );

    \I__12721\ : CascadeMux
    port map (
            O => \N__52794\,
            I => \N__52772\
        );

    \I__12720\ : CascadeMux
    port map (
            O => \N__52793\,
            I => \N__52764\
        );

    \I__12719\ : LocalMux
    port map (
            O => \N__52784\,
            I => \N__52759\
        );

    \I__12718\ : InMux
    port map (
            O => \N__52783\,
            I => \N__52756\
        );

    \I__12717\ : InMux
    port map (
            O => \N__52782\,
            I => \N__52753\
        );

    \I__12716\ : InMux
    port map (
            O => \N__52781\,
            I => \N__52750\
        );

    \I__12715\ : InMux
    port map (
            O => \N__52778\,
            I => \N__52745\
        );

    \I__12714\ : InMux
    port map (
            O => \N__52775\,
            I => \N__52745\
        );

    \I__12713\ : InMux
    port map (
            O => \N__52772\,
            I => \N__52740\
        );

    \I__12712\ : InMux
    port map (
            O => \N__52771\,
            I => \N__52740\
        );

    \I__12711\ : InMux
    port map (
            O => \N__52770\,
            I => \N__52727\
        );

    \I__12710\ : InMux
    port map (
            O => \N__52769\,
            I => \N__52727\
        );

    \I__12709\ : InMux
    port map (
            O => \N__52768\,
            I => \N__52727\
        );

    \I__12708\ : InMux
    port map (
            O => \N__52767\,
            I => \N__52727\
        );

    \I__12707\ : InMux
    port map (
            O => \N__52764\,
            I => \N__52727\
        );

    \I__12706\ : InMux
    port map (
            O => \N__52763\,
            I => \N__52727\
        );

    \I__12705\ : InMux
    port map (
            O => \N__52762\,
            I => \N__52724\
        );

    \I__12704\ : Span4Mux_h
    port map (
            O => \N__52759\,
            I => \N__52719\
        );

    \I__12703\ : LocalMux
    port map (
            O => \N__52756\,
            I => \N__52719\
        );

    \I__12702\ : LocalMux
    port map (
            O => \N__52753\,
            I => \N__52712\
        );

    \I__12701\ : LocalMux
    port map (
            O => \N__52750\,
            I => \N__52712\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__52745\,
            I => \N__52712\
        );

    \I__12699\ : LocalMux
    port map (
            O => \N__52740\,
            I => \N__52707\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__52727\,
            I => \N__52707\
        );

    \I__12697\ : LocalMux
    port map (
            O => \N__52724\,
            I => \N__52704\
        );

    \I__12696\ : Span4Mux_v
    port map (
            O => \N__52719\,
            I => \N__52701\
        );

    \I__12695\ : Span4Mux_v
    port map (
            O => \N__52712\,
            I => \N__52698\
        );

    \I__12694\ : Span4Mux_v
    port map (
            O => \N__52707\,
            I => \N__52695\
        );

    \I__12693\ : Span4Mux_h
    port map (
            O => \N__52704\,
            I => \N__52692\
        );

    \I__12692\ : Span4Mux_h
    port map (
            O => \N__52701\,
            I => \N__52685\
        );

    \I__12691\ : Span4Mux_h
    port map (
            O => \N__52698\,
            I => \N__52685\
        );

    \I__12690\ : Sp12to4
    port map (
            O => \N__52695\,
            I => \N__52682\
        );

    \I__12689\ : Span4Mux_v
    port map (
            O => \N__52692\,
            I => \N__52679\
        );

    \I__12688\ : InMux
    port map (
            O => \N__52691\,
            I => \N__52674\
        );

    \I__12687\ : InMux
    port map (
            O => \N__52690\,
            I => \N__52674\
        );

    \I__12686\ : Sp12to4
    port map (
            O => \N__52685\,
            I => \N__52669\
        );

    \I__12685\ : Span12Mux_h
    port map (
            O => \N__52682\,
            I => \N__52669\
        );

    \I__12684\ : Sp12to4
    port map (
            O => \N__52679\,
            I => \N__52664\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__52674\,
            I => \N__52664\
        );

    \I__12682\ : Span12Mux_v
    port map (
            O => \N__52669\,
            I => \N__52661\
        );

    \I__12681\ : Span12Mux_v
    port map (
            O => \N__52664\,
            I => \N__52658\
        );

    \I__12680\ : Odrv12
    port map (
            O => \N__52661\,
            I => \ICE_SPI_CE0\
        );

    \I__12679\ : Odrv12
    port map (
            O => \N__52658\,
            I => \ICE_SPI_CE0\
        );

    \I__12678\ : InMux
    port map (
            O => \N__52653\,
            I => \N__52650\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__52650\,
            I => n6401
        );

    \I__12676\ : SRMux
    port map (
            O => \N__52647\,
            I => \N__52644\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__52644\,
            I => \N__52641\
        );

    \I__12674\ : Span4Mux_h
    port map (
            O => \N__52641\,
            I => \N__52638\
        );

    \I__12673\ : Span4Mux_h
    port map (
            O => \N__52638\,
            I => \N__52635\
        );

    \I__12672\ : Odrv4
    port map (
            O => \N__52635\,
            I => n16821
        );

    \I__12671\ : InMux
    port map (
            O => \N__52632\,
            I => \N__52628\
        );

    \I__12670\ : InMux
    port map (
            O => \N__52631\,
            I => \N__52625\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__52628\,
            I => \N__52622\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__52625\,
            I => \N__52619\
        );

    \I__12667\ : Span4Mux_h
    port map (
            O => \N__52622\,
            I => \N__52616\
        );

    \I__12666\ : Span4Mux_h
    port map (
            O => \N__52619\,
            I => \N__52613\
        );

    \I__12665\ : Span4Mux_h
    port map (
            O => \N__52616\,
            I => \N__52610\
        );

    \I__12664\ : Span4Mux_h
    port map (
            O => \N__52613\,
            I => \N__52607\
        );

    \I__12663\ : Odrv4
    port map (
            O => \N__52610\,
            I => \comm_spi.n14842\
        );

    \I__12662\ : Odrv4
    port map (
            O => \N__52607\,
            I => \comm_spi.n14842\
        );

    \I__12661\ : InMux
    port map (
            O => \N__52602\,
            I => \N__52599\
        );

    \I__12660\ : LocalMux
    port map (
            O => \N__52599\,
            I => \N__52596\
        );

    \I__12659\ : Span4Mux_h
    port map (
            O => \N__52596\,
            I => \N__52593\
        );

    \I__12658\ : Odrv4
    port map (
            O => \N__52593\,
            I => buf_data_iac_18
        );

    \I__12657\ : InMux
    port map (
            O => \N__52590\,
            I => \N__52587\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__52587\,
            I => \N__52584\
        );

    \I__12655\ : Span4Mux_h
    port map (
            O => \N__52584\,
            I => \N__52581\
        );

    \I__12654\ : Odrv4
    port map (
            O => \N__52581\,
            I => n21460
        );

    \I__12653\ : InMux
    port map (
            O => \N__52578\,
            I => \N__52575\
        );

    \I__12652\ : LocalMux
    port map (
            O => \N__52575\,
            I => \N__52572\
        );

    \I__12651\ : Span12Mux_s11_h
    port map (
            O => \N__52572\,
            I => \N__52569\
        );

    \I__12650\ : Odrv12
    port map (
            O => \N__52569\,
            I => comm_buf_2_5
        );

    \I__12649\ : InMux
    port map (
            O => \N__52566\,
            I => \N__52546\
        );

    \I__12648\ : InMux
    port map (
            O => \N__52565\,
            I => \N__52546\
        );

    \I__12647\ : InMux
    port map (
            O => \N__52564\,
            I => \N__52546\
        );

    \I__12646\ : InMux
    port map (
            O => \N__52563\,
            I => \N__52539\
        );

    \I__12645\ : InMux
    port map (
            O => \N__52562\,
            I => \N__52539\
        );

    \I__12644\ : InMux
    port map (
            O => \N__52561\,
            I => \N__52539\
        );

    \I__12643\ : InMux
    port map (
            O => \N__52560\,
            I => \N__52532\
        );

    \I__12642\ : InMux
    port map (
            O => \N__52559\,
            I => \N__52532\
        );

    \I__12641\ : InMux
    port map (
            O => \N__52558\,
            I => \N__52532\
        );

    \I__12640\ : InMux
    port map (
            O => \N__52557\,
            I => \N__52527\
        );

    \I__12639\ : InMux
    port map (
            O => \N__52556\,
            I => \N__52527\
        );

    \I__12638\ : InMux
    port map (
            O => \N__52555\,
            I => \N__52524\
        );

    \I__12637\ : CascadeMux
    port map (
            O => \N__52554\,
            I => \N__52517\
        );

    \I__12636\ : InMux
    port map (
            O => \N__52553\,
            I => \N__52514\
        );

    \I__12635\ : LocalMux
    port map (
            O => \N__52546\,
            I => \N__52503\
        );

    \I__12634\ : LocalMux
    port map (
            O => \N__52539\,
            I => \N__52503\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__52532\,
            I => \N__52503\
        );

    \I__12632\ : LocalMux
    port map (
            O => \N__52527\,
            I => \N__52503\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__52524\,
            I => \N__52500\
        );

    \I__12630\ : InMux
    port map (
            O => \N__52523\,
            I => \N__52495\
        );

    \I__12629\ : InMux
    port map (
            O => \N__52522\,
            I => \N__52495\
        );

    \I__12628\ : InMux
    port map (
            O => \N__52521\,
            I => \N__52490\
        );

    \I__12627\ : InMux
    port map (
            O => \N__52520\,
            I => \N__52490\
        );

    \I__12626\ : InMux
    port map (
            O => \N__52517\,
            I => \N__52487\
        );

    \I__12625\ : LocalMux
    port map (
            O => \N__52514\,
            I => \N__52484\
        );

    \I__12624\ : InMux
    port map (
            O => \N__52513\,
            I => \N__52481\
        );

    \I__12623\ : InMux
    port map (
            O => \N__52512\,
            I => \N__52478\
        );

    \I__12622\ : Span4Mux_v
    port map (
            O => \N__52503\,
            I => \N__52475\
        );

    \I__12621\ : Span4Mux_v
    port map (
            O => \N__52500\,
            I => \N__52468\
        );

    \I__12620\ : LocalMux
    port map (
            O => \N__52495\,
            I => \N__52468\
        );

    \I__12619\ : LocalMux
    port map (
            O => \N__52490\,
            I => \N__52468\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__52487\,
            I => \N__52463\
        );

    \I__12617\ : Span4Mux_h
    port map (
            O => \N__52484\,
            I => \N__52463\
        );

    \I__12616\ : LocalMux
    port map (
            O => \N__52481\,
            I => \N__52460\
        );

    \I__12615\ : LocalMux
    port map (
            O => \N__52478\,
            I => comm_index_2
        );

    \I__12614\ : Odrv4
    port map (
            O => \N__52475\,
            I => comm_index_2
        );

    \I__12613\ : Odrv4
    port map (
            O => \N__52468\,
            I => comm_index_2
        );

    \I__12612\ : Odrv4
    port map (
            O => \N__52463\,
            I => comm_index_2
        );

    \I__12611\ : Odrv4
    port map (
            O => \N__52460\,
            I => comm_index_2
        );

    \I__12610\ : InMux
    port map (
            O => \N__52449\,
            I => \N__52440\
        );

    \I__12609\ : CascadeMux
    port map (
            O => \N__52448\,
            I => \N__52429\
        );

    \I__12608\ : InMux
    port map (
            O => \N__52447\,
            I => \N__52426\
        );

    \I__12607\ : InMux
    port map (
            O => \N__52446\,
            I => \N__52423\
        );

    \I__12606\ : InMux
    port map (
            O => \N__52445\,
            I => \N__52420\
        );

    \I__12605\ : InMux
    port map (
            O => \N__52444\,
            I => \N__52415\
        );

    \I__12604\ : InMux
    port map (
            O => \N__52443\,
            I => \N__52415\
        );

    \I__12603\ : LocalMux
    port map (
            O => \N__52440\,
            I => \N__52412\
        );

    \I__12602\ : CascadeMux
    port map (
            O => \N__52439\,
            I => \N__52406\
        );

    \I__12601\ : InMux
    port map (
            O => \N__52438\,
            I => \N__52401\
        );

    \I__12600\ : InMux
    port map (
            O => \N__52437\,
            I => \N__52401\
        );

    \I__12599\ : InMux
    port map (
            O => \N__52436\,
            I => \N__52396\
        );

    \I__12598\ : InMux
    port map (
            O => \N__52435\,
            I => \N__52396\
        );

    \I__12597\ : InMux
    port map (
            O => \N__52434\,
            I => \N__52383\
        );

    \I__12596\ : InMux
    port map (
            O => \N__52433\,
            I => \N__52383\
        );

    \I__12595\ : InMux
    port map (
            O => \N__52432\,
            I => \N__52383\
        );

    \I__12594\ : InMux
    port map (
            O => \N__52429\,
            I => \N__52383\
        );

    \I__12593\ : LocalMux
    port map (
            O => \N__52426\,
            I => \N__52371\
        );

    \I__12592\ : LocalMux
    port map (
            O => \N__52423\,
            I => \N__52371\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__52420\,
            I => \N__52364\
        );

    \I__12590\ : LocalMux
    port map (
            O => \N__52415\,
            I => \N__52364\
        );

    \I__12589\ : Span4Mux_v
    port map (
            O => \N__52412\,
            I => \N__52364\
        );

    \I__12588\ : InMux
    port map (
            O => \N__52411\,
            I => \N__52355\
        );

    \I__12587\ : InMux
    port map (
            O => \N__52410\,
            I => \N__52355\
        );

    \I__12586\ : InMux
    port map (
            O => \N__52409\,
            I => \N__52355\
        );

    \I__12585\ : InMux
    port map (
            O => \N__52406\,
            I => \N__52355\
        );

    \I__12584\ : LocalMux
    port map (
            O => \N__52401\,
            I => \N__52350\
        );

    \I__12583\ : LocalMux
    port map (
            O => \N__52396\,
            I => \N__52350\
        );

    \I__12582\ : InMux
    port map (
            O => \N__52395\,
            I => \N__52345\
        );

    \I__12581\ : InMux
    port map (
            O => \N__52394\,
            I => \N__52345\
        );

    \I__12580\ : InMux
    port map (
            O => \N__52393\,
            I => \N__52340\
        );

    \I__12579\ : InMux
    port map (
            O => \N__52392\,
            I => \N__52340\
        );

    \I__12578\ : LocalMux
    port map (
            O => \N__52383\,
            I => \N__52337\
        );

    \I__12577\ : InMux
    port map (
            O => \N__52382\,
            I => \N__52334\
        );

    \I__12576\ : InMux
    port map (
            O => \N__52381\,
            I => \N__52325\
        );

    \I__12575\ : InMux
    port map (
            O => \N__52380\,
            I => \N__52325\
        );

    \I__12574\ : InMux
    port map (
            O => \N__52379\,
            I => \N__52325\
        );

    \I__12573\ : InMux
    port map (
            O => \N__52378\,
            I => \N__52325\
        );

    \I__12572\ : InMux
    port map (
            O => \N__52377\,
            I => \N__52320\
        );

    \I__12571\ : InMux
    port map (
            O => \N__52376\,
            I => \N__52320\
        );

    \I__12570\ : Span4Mux_v
    port map (
            O => \N__52371\,
            I => \N__52313\
        );

    \I__12569\ : Span4Mux_v
    port map (
            O => \N__52364\,
            I => \N__52313\
        );

    \I__12568\ : LocalMux
    port map (
            O => \N__52355\,
            I => \N__52313\
        );

    \I__12567\ : Span4Mux_v
    port map (
            O => \N__52350\,
            I => \N__52304\
        );

    \I__12566\ : LocalMux
    port map (
            O => \N__52345\,
            I => \N__52304\
        );

    \I__12565\ : LocalMux
    port map (
            O => \N__52340\,
            I => \N__52304\
        );

    \I__12564\ : Span4Mux_h
    port map (
            O => \N__52337\,
            I => \N__52304\
        );

    \I__12563\ : LocalMux
    port map (
            O => \N__52334\,
            I => \N__52299\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__52325\,
            I => \N__52299\
        );

    \I__12561\ : LocalMux
    port map (
            O => \N__52320\,
            I => comm_index_1
        );

    \I__12560\ : Odrv4
    port map (
            O => \N__52313\,
            I => comm_index_1
        );

    \I__12559\ : Odrv4
    port map (
            O => \N__52304\,
            I => comm_index_1
        );

    \I__12558\ : Odrv12
    port map (
            O => \N__52299\,
            I => comm_index_1
        );

    \I__12557\ : CascadeMux
    port map (
            O => \N__52290\,
            I => \N__52287\
        );

    \I__12556\ : InMux
    port map (
            O => \N__52287\,
            I => \N__52282\
        );

    \I__12555\ : CascadeMux
    port map (
            O => \N__52286\,
            I => \N__52279\
        );

    \I__12554\ : InMux
    port map (
            O => \N__52285\,
            I => \N__52272\
        );

    \I__12553\ : LocalMux
    port map (
            O => \N__52282\,
            I => \N__52269\
        );

    \I__12552\ : InMux
    port map (
            O => \N__52279\,
            I => \N__52266\
        );

    \I__12551\ : InMux
    port map (
            O => \N__52278\,
            I => \N__52263\
        );

    \I__12550\ : InMux
    port map (
            O => \N__52277\,
            I => \N__52260\
        );

    \I__12549\ : CascadeMux
    port map (
            O => \N__52276\,
            I => \N__52257\
        );

    \I__12548\ : CascadeMux
    port map (
            O => \N__52275\,
            I => \N__52254\
        );

    \I__12547\ : LocalMux
    port map (
            O => \N__52272\,
            I => \N__52251\
        );

    \I__12546\ : Span4Mux_h
    port map (
            O => \N__52269\,
            I => \N__52246\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__52266\,
            I => \N__52246\
        );

    \I__12544\ : LocalMux
    port map (
            O => \N__52263\,
            I => \N__52243\
        );

    \I__12543\ : LocalMux
    port map (
            O => \N__52260\,
            I => \N__52240\
        );

    \I__12542\ : InMux
    port map (
            O => \N__52257\,
            I => \N__52237\
        );

    \I__12541\ : InMux
    port map (
            O => \N__52254\,
            I => \N__52234\
        );

    \I__12540\ : Span12Mux_v
    port map (
            O => \N__52251\,
            I => \N__52231\
        );

    \I__12539\ : Span4Mux_h
    port map (
            O => \N__52246\,
            I => \N__52228\
        );

    \I__12538\ : Span4Mux_h
    port map (
            O => \N__52243\,
            I => \N__52225\
        );

    \I__12537\ : Span4Mux_v
    port map (
            O => \N__52240\,
            I => \N__52220\
        );

    \I__12536\ : LocalMux
    port map (
            O => \N__52237\,
            I => \N__52220\
        );

    \I__12535\ : LocalMux
    port map (
            O => \N__52234\,
            I => \N__52217\
        );

    \I__12534\ : Span12Mux_h
    port map (
            O => \N__52231\,
            I => \N__52214\
        );

    \I__12533\ : Span4Mux_v
    port map (
            O => \N__52228\,
            I => \N__52209\
        );

    \I__12532\ : Span4Mux_h
    port map (
            O => \N__52225\,
            I => \N__52209\
        );

    \I__12531\ : Odrv4
    port map (
            O => \N__52220\,
            I => comm_buf_0_5
        );

    \I__12530\ : Odrv12
    port map (
            O => \N__52217\,
            I => comm_buf_0_5
        );

    \I__12529\ : Odrv12
    port map (
            O => \N__52214\,
            I => comm_buf_0_5
        );

    \I__12528\ : Odrv4
    port map (
            O => \N__52209\,
            I => comm_buf_0_5
        );

    \I__12527\ : CascadeMux
    port map (
            O => \N__52200\,
            I => \n22503_cascade_\
        );

    \I__12526\ : InMux
    port map (
            O => \N__52197\,
            I => \N__52194\
        );

    \I__12525\ : LocalMux
    port map (
            O => \N__52194\,
            I => \N__52191\
        );

    \I__12524\ : Span4Mux_h
    port map (
            O => \N__52191\,
            I => \N__52188\
        );

    \I__12523\ : Span4Mux_v
    port map (
            O => \N__52188\,
            I => \N__52185\
        );

    \I__12522\ : Odrv4
    port map (
            O => \N__52185\,
            I => comm_buf_4_5
        );

    \I__12521\ : InMux
    port map (
            O => \N__52182\,
            I => \N__52179\
        );

    \I__12520\ : LocalMux
    port map (
            O => \N__52179\,
            I => \N__52176\
        );

    \I__12519\ : Odrv4
    port map (
            O => \N__52176\,
            I => n22506
        );

    \I__12518\ : InMux
    port map (
            O => \N__52173\,
            I => \ADC_VDC.genclk.n19902\
        );

    \I__12517\ : CEMux
    port map (
            O => \N__52170\,
            I => \N__52166\
        );

    \I__12516\ : CEMux
    port map (
            O => \N__52169\,
            I => \N__52163\
        );

    \I__12515\ : LocalMux
    port map (
            O => \N__52166\,
            I => \N__52160\
        );

    \I__12514\ : LocalMux
    port map (
            O => \N__52163\,
            I => \N__52157\
        );

    \I__12513\ : Odrv12
    port map (
            O => \N__52160\,
            I => \ADC_VDC.genclk.n11900\
        );

    \I__12512\ : Odrv4
    port map (
            O => \N__52157\,
            I => \ADC_VDC.genclk.n11900\
        );

    \I__12511\ : CascadeMux
    port map (
            O => \N__52152\,
            I => \N__52147\
        );

    \I__12510\ : InMux
    port map (
            O => \N__52151\,
            I => \N__52144\
        );

    \I__12509\ : InMux
    port map (
            O => \N__52150\,
            I => \N__52141\
        );

    \I__12508\ : InMux
    port map (
            O => \N__52147\,
            I => \N__52138\
        );

    \I__12507\ : LocalMux
    port map (
            O => \N__52144\,
            I => \N__52135\
        );

    \I__12506\ : LocalMux
    port map (
            O => \N__52141\,
            I => \N__52132\
        );

    \I__12505\ : LocalMux
    port map (
            O => \N__52138\,
            I => \N__52129\
        );

    \I__12504\ : Odrv4
    port map (
            O => \N__52135\,
            I => n14350
        );

    \I__12503\ : Odrv4
    port map (
            O => \N__52132\,
            I => n14350
        );

    \I__12502\ : Odrv4
    port map (
            O => \N__52129\,
            I => n14350
        );

    \I__12501\ : InMux
    port map (
            O => \N__52122\,
            I => \N__52119\
        );

    \I__12500\ : LocalMux
    port map (
            O => \N__52119\,
            I => n21453
        );

    \I__12499\ : CascadeMux
    port map (
            O => \N__52116\,
            I => \n21454_cascade_\
        );

    \I__12498\ : CEMux
    port map (
            O => \N__52113\,
            I => \N__52110\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__52110\,
            I => n14_adj_1638
        );

    \I__12496\ : InMux
    port map (
            O => \N__52107\,
            I => \N__52104\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__52104\,
            I => \N__52101\
        );

    \I__12494\ : Span4Mux_h
    port map (
            O => \N__52101\,
            I => \N__52098\
        );

    \I__12493\ : Odrv4
    port map (
            O => \N__52098\,
            I => n21481
        );

    \I__12492\ : CEMux
    port map (
            O => \N__52095\,
            I => \N__52091\
        );

    \I__12491\ : InMux
    port map (
            O => \N__52094\,
            I => \N__52087\
        );

    \I__12490\ : LocalMux
    port map (
            O => \N__52091\,
            I => \N__52084\
        );

    \I__12489\ : InMux
    port map (
            O => \N__52090\,
            I => \N__52081\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__52087\,
            I => \N__52078\
        );

    \I__12487\ : Span4Mux_v
    port map (
            O => \N__52084\,
            I => \N__52075\
        );

    \I__12486\ : LocalMux
    port map (
            O => \N__52081\,
            I => \N__52072\
        );

    \I__12485\ : Span4Mux_h
    port map (
            O => \N__52078\,
            I => \N__52069\
        );

    \I__12484\ : Span4Mux_h
    port map (
            O => \N__52075\,
            I => \N__52064\
        );

    \I__12483\ : Span4Mux_v
    port map (
            O => \N__52072\,
            I => \N__52064\
        );

    \I__12482\ : Span4Mux_h
    port map (
            O => \N__52069\,
            I => \N__52059\
        );

    \I__12481\ : Span4Mux_h
    port map (
            O => \N__52064\,
            I => \N__52059\
        );

    \I__12480\ : Odrv4
    port map (
            O => \N__52059\,
            I => n12089
        );

    \I__12479\ : InMux
    port map (
            O => \N__52056\,
            I => \N__52052\
        );

    \I__12478\ : InMux
    port map (
            O => \N__52055\,
            I => \N__52049\
        );

    \I__12477\ : LocalMux
    port map (
            O => \N__52052\,
            I => comm_length_2
        );

    \I__12476\ : LocalMux
    port map (
            O => \N__52049\,
            I => comm_length_2
        );

    \I__12475\ : InMux
    port map (
            O => \N__52044\,
            I => \N__52041\
        );

    \I__12474\ : LocalMux
    port map (
            O => \N__52041\,
            I => n6541
        );

    \I__12473\ : InMux
    port map (
            O => \N__52038\,
            I => \N__52035\
        );

    \I__12472\ : LocalMux
    port map (
            O => \N__52035\,
            I => n21154
        );

    \I__12471\ : InMux
    port map (
            O => \N__52032\,
            I => \ADC_VDC.genclk.n19893\
        );

    \I__12470\ : InMux
    port map (
            O => \N__52029\,
            I => \ADC_VDC.genclk.n19894\
        );

    \I__12469\ : InMux
    port map (
            O => \N__52026\,
            I => \bfn_19_8_0_\
        );

    \I__12468\ : InMux
    port map (
            O => \N__52023\,
            I => \ADC_VDC.genclk.n19896\
        );

    \I__12467\ : InMux
    port map (
            O => \N__52020\,
            I => \ADC_VDC.genclk.n19897\
        );

    \I__12466\ : InMux
    port map (
            O => \N__52017\,
            I => \ADC_VDC.genclk.n19898\
        );

    \I__12465\ : InMux
    port map (
            O => \N__52014\,
            I => \ADC_VDC.genclk.n19899\
        );

    \I__12464\ : InMux
    port map (
            O => \N__52011\,
            I => \ADC_VDC.genclk.n19900\
        );

    \I__12463\ : InMux
    port map (
            O => \N__52008\,
            I => \ADC_VDC.genclk.n19901\
        );

    \I__12462\ : InMux
    port map (
            O => \N__52005\,
            I => \N__52001\
        );

    \I__12461\ : CascadeMux
    port map (
            O => \N__52004\,
            I => \N__51997\
        );

    \I__12460\ : LocalMux
    port map (
            O => \N__52001\,
            I => \N__51994\
        );

    \I__12459\ : CascadeMux
    port map (
            O => \N__52000\,
            I => \N__51990\
        );

    \I__12458\ : InMux
    port map (
            O => \N__51997\,
            I => \N__51987\
        );

    \I__12457\ : Span4Mux_v
    port map (
            O => \N__51994\,
            I => \N__51982\
        );

    \I__12456\ : InMux
    port map (
            O => \N__51993\,
            I => \N__51979\
        );

    \I__12455\ : InMux
    port map (
            O => \N__51990\,
            I => \N__51976\
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__51987\,
            I => \N__51971\
        );

    \I__12453\ : InMux
    port map (
            O => \N__51986\,
            I => \N__51966\
        );

    \I__12452\ : InMux
    port map (
            O => \N__51985\,
            I => \N__51966\
        );

    \I__12451\ : Span4Mux_h
    port map (
            O => \N__51982\,
            I => \N__51959\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__51979\,
            I => \N__51959\
        );

    \I__12449\ : LocalMux
    port map (
            O => \N__51976\,
            I => \N__51959\
        );

    \I__12448\ : InMux
    port map (
            O => \N__51975\,
            I => \N__51954\
        );

    \I__12447\ : InMux
    port map (
            O => \N__51974\,
            I => \N__51954\
        );

    \I__12446\ : Span4Mux_v
    port map (
            O => \N__51971\,
            I => \N__51951\
        );

    \I__12445\ : LocalMux
    port map (
            O => \N__51966\,
            I => \N__51948\
        );

    \I__12444\ : Span4Mux_h
    port map (
            O => \N__51959\,
            I => \N__51943\
        );

    \I__12443\ : LocalMux
    port map (
            O => \N__51954\,
            I => \N__51943\
        );

    \I__12442\ : Span4Mux_h
    port map (
            O => \N__51951\,
            I => \N__51939\
        );

    \I__12441\ : Span4Mux_h
    port map (
            O => \N__51948\,
            I => \N__51934\
        );

    \I__12440\ : Span4Mux_h
    port map (
            O => \N__51943\,
            I => \N__51934\
        );

    \I__12439\ : InMux
    port map (
            O => \N__51942\,
            I => \N__51931\
        );

    \I__12438\ : Span4Mux_v
    port map (
            O => \N__51939\,
            I => \N__51928\
        );

    \I__12437\ : Sp12to4
    port map (
            O => \N__51934\,
            I => \N__51923\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__51931\,
            I => \N__51923\
        );

    \I__12435\ : Sp12to4
    port map (
            O => \N__51928\,
            I => \N__51918\
        );

    \I__12434\ : Span12Mux_v
    port map (
            O => \N__51923\,
            I => \N__51918\
        );

    \I__12433\ : Odrv12
    port map (
            O => \N__51918\,
            I => \VDC_SDO\
        );

    \I__12432\ : CascadeMux
    port map (
            O => \N__51915\,
            I => \N__51912\
        );

    \I__12431\ : InMux
    port map (
            O => \N__51912\,
            I => \N__51905\
        );

    \I__12430\ : InMux
    port map (
            O => \N__51911\,
            I => \N__51900\
        );

    \I__12429\ : CascadeMux
    port map (
            O => \N__51910\,
            I => \N__51897\
        );

    \I__12428\ : CascadeMux
    port map (
            O => \N__51909\,
            I => \N__51889\
        );

    \I__12427\ : InMux
    port map (
            O => \N__51908\,
            I => \N__51886\
        );

    \I__12426\ : LocalMux
    port map (
            O => \N__51905\,
            I => \N__51883\
        );

    \I__12425\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51877\
        );

    \I__12424\ : InMux
    port map (
            O => \N__51903\,
            I => \N__51874\
        );

    \I__12423\ : LocalMux
    port map (
            O => \N__51900\,
            I => \N__51871\
        );

    \I__12422\ : InMux
    port map (
            O => \N__51897\,
            I => \N__51868\
        );

    \I__12421\ : InMux
    port map (
            O => \N__51896\,
            I => \N__51864\
        );

    \I__12420\ : InMux
    port map (
            O => \N__51895\,
            I => \N__51861\
        );

    \I__12419\ : InMux
    port map (
            O => \N__51894\,
            I => \N__51853\
        );

    \I__12418\ : InMux
    port map (
            O => \N__51893\,
            I => \N__51846\
        );

    \I__12417\ : InMux
    port map (
            O => \N__51892\,
            I => \N__51846\
        );

    \I__12416\ : InMux
    port map (
            O => \N__51889\,
            I => \N__51846\
        );

    \I__12415\ : LocalMux
    port map (
            O => \N__51886\,
            I => \N__51843\
        );

    \I__12414\ : Span4Mux_h
    port map (
            O => \N__51883\,
            I => \N__51840\
        );

    \I__12413\ : InMux
    port map (
            O => \N__51882\,
            I => \N__51833\
        );

    \I__12412\ : InMux
    port map (
            O => \N__51881\,
            I => \N__51833\
        );

    \I__12411\ : InMux
    port map (
            O => \N__51880\,
            I => \N__51833\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__51877\,
            I => \N__51828\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__51874\,
            I => \N__51828\
        );

    \I__12408\ : Span4Mux_v
    port map (
            O => \N__51871\,
            I => \N__51823\
        );

    \I__12407\ : LocalMux
    port map (
            O => \N__51868\,
            I => \N__51823\
        );

    \I__12406\ : InMux
    port map (
            O => \N__51867\,
            I => \N__51820\
        );

    \I__12405\ : LocalMux
    port map (
            O => \N__51864\,
            I => \N__51817\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__51861\,
            I => \N__51814\
        );

    \I__12403\ : InMux
    port map (
            O => \N__51860\,
            I => \N__51811\
        );

    \I__12402\ : InMux
    port map (
            O => \N__51859\,
            I => \N__51806\
        );

    \I__12401\ : InMux
    port map (
            O => \N__51858\,
            I => \N__51806\
        );

    \I__12400\ : InMux
    port map (
            O => \N__51857\,
            I => \N__51803\
        );

    \I__12399\ : InMux
    port map (
            O => \N__51856\,
            I => \N__51800\
        );

    \I__12398\ : LocalMux
    port map (
            O => \N__51853\,
            I => \N__51789\
        );

    \I__12397\ : LocalMux
    port map (
            O => \N__51846\,
            I => \N__51789\
        );

    \I__12396\ : Span4Mux_v
    port map (
            O => \N__51843\,
            I => \N__51789\
        );

    \I__12395\ : Span4Mux_v
    port map (
            O => \N__51840\,
            I => \N__51789\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__51833\,
            I => \N__51789\
        );

    \I__12393\ : Span12Mux_h
    port map (
            O => \N__51828\,
            I => \N__51786\
        );

    \I__12392\ : Span4Mux_h
    port map (
            O => \N__51823\,
            I => \N__51783\
        );

    \I__12391\ : LocalMux
    port map (
            O => \N__51820\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12390\ : Odrv4
    port map (
            O => \N__51817\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12389\ : Odrv12
    port map (
            O => \N__51814\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12388\ : LocalMux
    port map (
            O => \N__51811\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12387\ : LocalMux
    port map (
            O => \N__51806\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__51803\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__51800\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12384\ : Odrv4
    port map (
            O => \N__51789\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12383\ : Odrv12
    port map (
            O => \N__51786\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12382\ : Odrv4
    port map (
            O => \N__51783\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__12381\ : CascadeMux
    port map (
            O => \N__51762\,
            I => \N__51755\
        );

    \I__12380\ : CascadeMux
    port map (
            O => \N__51761\,
            I => \N__51750\
        );

    \I__12379\ : InMux
    port map (
            O => \N__51760\,
            I => \N__51747\
        );

    \I__12378\ : CascadeMux
    port map (
            O => \N__51759\,
            I => \N__51741\
        );

    \I__12377\ : CascadeMux
    port map (
            O => \N__51758\,
            I => \N__51738\
        );

    \I__12376\ : InMux
    port map (
            O => \N__51755\,
            I => \N__51735\
        );

    \I__12375\ : CascadeMux
    port map (
            O => \N__51754\,
            I => \N__51732\
        );

    \I__12374\ : InMux
    port map (
            O => \N__51753\,
            I => \N__51729\
        );

    \I__12373\ : InMux
    port map (
            O => \N__51750\,
            I => \N__51726\
        );

    \I__12372\ : LocalMux
    port map (
            O => \N__51747\,
            I => \N__51723\
        );

    \I__12371\ : InMux
    port map (
            O => \N__51746\,
            I => \N__51717\
        );

    \I__12370\ : InMux
    port map (
            O => \N__51745\,
            I => \N__51714\
        );

    \I__12369\ : InMux
    port map (
            O => \N__51744\,
            I => \N__51691\
        );

    \I__12368\ : InMux
    port map (
            O => \N__51741\,
            I => \N__51691\
        );

    \I__12367\ : InMux
    port map (
            O => \N__51738\,
            I => \N__51687\
        );

    \I__12366\ : LocalMux
    port map (
            O => \N__51735\,
            I => \N__51684\
        );

    \I__12365\ : InMux
    port map (
            O => \N__51732\,
            I => \N__51681\
        );

    \I__12364\ : LocalMux
    port map (
            O => \N__51729\,
            I => \N__51674\
        );

    \I__12363\ : LocalMux
    port map (
            O => \N__51726\,
            I => \N__51674\
        );

    \I__12362\ : Span4Mux_v
    port map (
            O => \N__51723\,
            I => \N__51674\
        );

    \I__12361\ : InMux
    port map (
            O => \N__51722\,
            I => \N__51669\
        );

    \I__12360\ : InMux
    port map (
            O => \N__51721\,
            I => \N__51669\
        );

    \I__12359\ : InMux
    port map (
            O => \N__51720\,
            I => \N__51666\
        );

    \I__12358\ : LocalMux
    port map (
            O => \N__51717\,
            I => \N__51661\
        );

    \I__12357\ : LocalMux
    port map (
            O => \N__51714\,
            I => \N__51661\
        );

    \I__12356\ : InMux
    port map (
            O => \N__51713\,
            I => \N__51652\
        );

    \I__12355\ : InMux
    port map (
            O => \N__51712\,
            I => \N__51652\
        );

    \I__12354\ : InMux
    port map (
            O => \N__51711\,
            I => \N__51652\
        );

    \I__12353\ : InMux
    port map (
            O => \N__51710\,
            I => \N__51652\
        );

    \I__12352\ : CascadeMux
    port map (
            O => \N__51709\,
            I => \N__51649\
        );

    \I__12351\ : CascadeMux
    port map (
            O => \N__51708\,
            I => \N__51645\
        );

    \I__12350\ : CascadeMux
    port map (
            O => \N__51707\,
            I => \N__51642\
        );

    \I__12349\ : InMux
    port map (
            O => \N__51706\,
            I => \N__51625\
        );

    \I__12348\ : InMux
    port map (
            O => \N__51705\,
            I => \N__51625\
        );

    \I__12347\ : InMux
    port map (
            O => \N__51704\,
            I => \N__51625\
        );

    \I__12346\ : InMux
    port map (
            O => \N__51703\,
            I => \N__51625\
        );

    \I__12345\ : InMux
    port map (
            O => \N__51702\,
            I => \N__51616\
        );

    \I__12344\ : InMux
    port map (
            O => \N__51701\,
            I => \N__51616\
        );

    \I__12343\ : InMux
    port map (
            O => \N__51700\,
            I => \N__51616\
        );

    \I__12342\ : InMux
    port map (
            O => \N__51699\,
            I => \N__51616\
        );

    \I__12341\ : InMux
    port map (
            O => \N__51698\,
            I => \N__51609\
        );

    \I__12340\ : InMux
    port map (
            O => \N__51697\,
            I => \N__51609\
        );

    \I__12339\ : InMux
    port map (
            O => \N__51696\,
            I => \N__51609\
        );

    \I__12338\ : LocalMux
    port map (
            O => \N__51691\,
            I => \N__51606\
        );

    \I__12337\ : InMux
    port map (
            O => \N__51690\,
            I => \N__51603\
        );

    \I__12336\ : LocalMux
    port map (
            O => \N__51687\,
            I => \N__51596\
        );

    \I__12335\ : Span4Mux_v
    port map (
            O => \N__51684\,
            I => \N__51593\
        );

    \I__12334\ : LocalMux
    port map (
            O => \N__51681\,
            I => \N__51590\
        );

    \I__12333\ : Span4Mux_h
    port map (
            O => \N__51674\,
            I => \N__51587\
        );

    \I__12332\ : LocalMux
    port map (
            O => \N__51669\,
            I => \N__51578\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__51666\,
            I => \N__51578\
        );

    \I__12330\ : Span4Mux_v
    port map (
            O => \N__51661\,
            I => \N__51578\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__51652\,
            I => \N__51578\
        );

    \I__12328\ : InMux
    port map (
            O => \N__51649\,
            I => \N__51575\
        );

    \I__12327\ : InMux
    port map (
            O => \N__51648\,
            I => \N__51560\
        );

    \I__12326\ : InMux
    port map (
            O => \N__51645\,
            I => \N__51560\
        );

    \I__12325\ : InMux
    port map (
            O => \N__51642\,
            I => \N__51560\
        );

    \I__12324\ : InMux
    port map (
            O => \N__51641\,
            I => \N__51560\
        );

    \I__12323\ : InMux
    port map (
            O => \N__51640\,
            I => \N__51560\
        );

    \I__12322\ : InMux
    port map (
            O => \N__51639\,
            I => \N__51560\
        );

    \I__12321\ : InMux
    port map (
            O => \N__51638\,
            I => \N__51560\
        );

    \I__12320\ : InMux
    port map (
            O => \N__51637\,
            I => \N__51557\
        );

    \I__12319\ : InMux
    port map (
            O => \N__51636\,
            I => \N__51550\
        );

    \I__12318\ : InMux
    port map (
            O => \N__51635\,
            I => \N__51550\
        );

    \I__12317\ : InMux
    port map (
            O => \N__51634\,
            I => \N__51550\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__51625\,
            I => \N__51539\
        );

    \I__12315\ : LocalMux
    port map (
            O => \N__51616\,
            I => \N__51539\
        );

    \I__12314\ : LocalMux
    port map (
            O => \N__51609\,
            I => \N__51539\
        );

    \I__12313\ : Span4Mux_v
    port map (
            O => \N__51606\,
            I => \N__51539\
        );

    \I__12312\ : LocalMux
    port map (
            O => \N__51603\,
            I => \N__51539\
        );

    \I__12311\ : InMux
    port map (
            O => \N__51602\,
            I => \N__51530\
        );

    \I__12310\ : InMux
    port map (
            O => \N__51601\,
            I => \N__51530\
        );

    \I__12309\ : InMux
    port map (
            O => \N__51600\,
            I => \N__51530\
        );

    \I__12308\ : InMux
    port map (
            O => \N__51599\,
            I => \N__51530\
        );

    \I__12307\ : Span4Mux_v
    port map (
            O => \N__51596\,
            I => \N__51521\
        );

    \I__12306\ : Span4Mux_h
    port map (
            O => \N__51593\,
            I => \N__51521\
        );

    \I__12305\ : Span4Mux_v
    port map (
            O => \N__51590\,
            I => \N__51521\
        );

    \I__12304\ : Span4Mux_h
    port map (
            O => \N__51587\,
            I => \N__51521\
        );

    \I__12303\ : Span4Mux_h
    port map (
            O => \N__51578\,
            I => \N__51518\
        );

    \I__12302\ : LocalMux
    port map (
            O => \N__51575\,
            I => adc_state_3
        );

    \I__12301\ : LocalMux
    port map (
            O => \N__51560\,
            I => adc_state_3
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__51557\,
            I => adc_state_3
        );

    \I__12299\ : LocalMux
    port map (
            O => \N__51550\,
            I => adc_state_3
        );

    \I__12298\ : Odrv4
    port map (
            O => \N__51539\,
            I => adc_state_3
        );

    \I__12297\ : LocalMux
    port map (
            O => \N__51530\,
            I => adc_state_3
        );

    \I__12296\ : Odrv4
    port map (
            O => \N__51521\,
            I => adc_state_3
        );

    \I__12295\ : Odrv4
    port map (
            O => \N__51518\,
            I => adc_state_3
        );

    \I__12294\ : CascadeMux
    port map (
            O => \N__51501\,
            I => \N__51485\
        );

    \I__12293\ : InMux
    port map (
            O => \N__51500\,
            I => \N__51470\
        );

    \I__12292\ : InMux
    port map (
            O => \N__51499\,
            I => \N__51457\
        );

    \I__12291\ : InMux
    port map (
            O => \N__51498\,
            I => \N__51457\
        );

    \I__12290\ : InMux
    port map (
            O => \N__51497\,
            I => \N__51457\
        );

    \I__12289\ : InMux
    port map (
            O => \N__51496\,
            I => \N__51457\
        );

    \I__12288\ : InMux
    port map (
            O => \N__51495\,
            I => \N__51457\
        );

    \I__12287\ : InMux
    port map (
            O => \N__51494\,
            I => \N__51457\
        );

    \I__12286\ : InMux
    port map (
            O => \N__51493\,
            I => \N__51452\
        );

    \I__12285\ : InMux
    port map (
            O => \N__51492\,
            I => \N__51449\
        );

    \I__12284\ : CascadeMux
    port map (
            O => \N__51491\,
            I => \N__51446\
        );

    \I__12283\ : CascadeMux
    port map (
            O => \N__51490\,
            I => \N__51443\
        );

    \I__12282\ : InMux
    port map (
            O => \N__51489\,
            I => \N__51437\
        );

    \I__12281\ : InMux
    port map (
            O => \N__51488\,
            I => \N__51437\
        );

    \I__12280\ : InMux
    port map (
            O => \N__51485\,
            I => \N__51424\
        );

    \I__12279\ : InMux
    port map (
            O => \N__51484\,
            I => \N__51424\
        );

    \I__12278\ : InMux
    port map (
            O => \N__51483\,
            I => \N__51424\
        );

    \I__12277\ : InMux
    port map (
            O => \N__51482\,
            I => \N__51424\
        );

    \I__12276\ : InMux
    port map (
            O => \N__51481\,
            I => \N__51424\
        );

    \I__12275\ : InMux
    port map (
            O => \N__51480\,
            I => \N__51424\
        );

    \I__12274\ : InMux
    port map (
            O => \N__51479\,
            I => \N__51421\
        );

    \I__12273\ : InMux
    port map (
            O => \N__51478\,
            I => \N__51416\
        );

    \I__12272\ : InMux
    port map (
            O => \N__51477\,
            I => \N__51416\
        );

    \I__12271\ : InMux
    port map (
            O => \N__51476\,
            I => \N__51409\
        );

    \I__12270\ : InMux
    port map (
            O => \N__51475\,
            I => \N__51402\
        );

    \I__12269\ : InMux
    port map (
            O => \N__51474\,
            I => \N__51402\
        );

    \I__12268\ : InMux
    port map (
            O => \N__51473\,
            I => \N__51402\
        );

    \I__12267\ : LocalMux
    port map (
            O => \N__51470\,
            I => \N__51399\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__51457\,
            I => \N__51396\
        );

    \I__12265\ : InMux
    port map (
            O => \N__51456\,
            I => \N__51391\
        );

    \I__12264\ : InMux
    port map (
            O => \N__51455\,
            I => \N__51391\
        );

    \I__12263\ : LocalMux
    port map (
            O => \N__51452\,
            I => \N__51386\
        );

    \I__12262\ : LocalMux
    port map (
            O => \N__51449\,
            I => \N__51386\
        );

    \I__12261\ : InMux
    port map (
            O => \N__51446\,
            I => \N__51380\
        );

    \I__12260\ : InMux
    port map (
            O => \N__51443\,
            I => \N__51380\
        );

    \I__12259\ : InMux
    port map (
            O => \N__51442\,
            I => \N__51377\
        );

    \I__12258\ : LocalMux
    port map (
            O => \N__51437\,
            I => \N__51374\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__51424\,
            I => \N__51371\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__51421\,
            I => \N__51368\
        );

    \I__12255\ : LocalMux
    port map (
            O => \N__51416\,
            I => \N__51365\
        );

    \I__12254\ : CascadeMux
    port map (
            O => \N__51415\,
            I => \N__51358\
        );

    \I__12253\ : CascadeMux
    port map (
            O => \N__51414\,
            I => \N__51352\
        );

    \I__12252\ : InMux
    port map (
            O => \N__51413\,
            I => \N__51349\
        );

    \I__12251\ : InMux
    port map (
            O => \N__51412\,
            I => \N__51346\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__51409\,
            I => \N__51339\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__51402\,
            I => \N__51339\
        );

    \I__12248\ : Span4Mux_h
    port map (
            O => \N__51399\,
            I => \N__51332\
        );

    \I__12247\ : Span4Mux_h
    port map (
            O => \N__51396\,
            I => \N__51332\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__51391\,
            I => \N__51332\
        );

    \I__12245\ : Span4Mux_h
    port map (
            O => \N__51386\,
            I => \N__51324\
        );

    \I__12244\ : InMux
    port map (
            O => \N__51385\,
            I => \N__51321\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__51380\,
            I => \N__51312\
        );

    \I__12242\ : LocalMux
    port map (
            O => \N__51377\,
            I => \N__51312\
        );

    \I__12241\ : Span4Mux_h
    port map (
            O => \N__51374\,
            I => \N__51312\
        );

    \I__12240\ : Span4Mux_v
    port map (
            O => \N__51371\,
            I => \N__51312\
        );

    \I__12239\ : Span4Mux_v
    port map (
            O => \N__51368\,
            I => \N__51309\
        );

    \I__12238\ : Span4Mux_h
    port map (
            O => \N__51365\,
            I => \N__51306\
        );

    \I__12237\ : InMux
    port map (
            O => \N__51364\,
            I => \N__51295\
        );

    \I__12236\ : InMux
    port map (
            O => \N__51363\,
            I => \N__51295\
        );

    \I__12235\ : InMux
    port map (
            O => \N__51362\,
            I => \N__51295\
        );

    \I__12234\ : InMux
    port map (
            O => \N__51361\,
            I => \N__51295\
        );

    \I__12233\ : InMux
    port map (
            O => \N__51358\,
            I => \N__51295\
        );

    \I__12232\ : InMux
    port map (
            O => \N__51357\,
            I => \N__51286\
        );

    \I__12231\ : InMux
    port map (
            O => \N__51356\,
            I => \N__51286\
        );

    \I__12230\ : InMux
    port map (
            O => \N__51355\,
            I => \N__51286\
        );

    \I__12229\ : InMux
    port map (
            O => \N__51352\,
            I => \N__51286\
        );

    \I__12228\ : LocalMux
    port map (
            O => \N__51349\,
            I => \N__51281\
        );

    \I__12227\ : LocalMux
    port map (
            O => \N__51346\,
            I => \N__51281\
        );

    \I__12226\ : InMux
    port map (
            O => \N__51345\,
            I => \N__51278\
        );

    \I__12225\ : InMux
    port map (
            O => \N__51344\,
            I => \N__51275\
        );

    \I__12224\ : Span4Mux_v
    port map (
            O => \N__51339\,
            I => \N__51272\
        );

    \I__12223\ : Span4Mux_v
    port map (
            O => \N__51332\,
            I => \N__51269\
        );

    \I__12222\ : InMux
    port map (
            O => \N__51331\,
            I => \N__51264\
        );

    \I__12221\ : InMux
    port map (
            O => \N__51330\,
            I => \N__51264\
        );

    \I__12220\ : InMux
    port map (
            O => \N__51329\,
            I => \N__51257\
        );

    \I__12219\ : InMux
    port map (
            O => \N__51328\,
            I => \N__51257\
        );

    \I__12218\ : InMux
    port map (
            O => \N__51327\,
            I => \N__51257\
        );

    \I__12217\ : Span4Mux_h
    port map (
            O => \N__51324\,
            I => \N__51254\
        );

    \I__12216\ : LocalMux
    port map (
            O => \N__51321\,
            I => \N__51251\
        );

    \I__12215\ : Span4Mux_v
    port map (
            O => \N__51312\,
            I => \N__51246\
        );

    \I__12214\ : Span4Mux_h
    port map (
            O => \N__51309\,
            I => \N__51246\
        );

    \I__12213\ : Span4Mux_v
    port map (
            O => \N__51306\,
            I => \N__51237\
        );

    \I__12212\ : LocalMux
    port map (
            O => \N__51295\,
            I => \N__51237\
        );

    \I__12211\ : LocalMux
    port map (
            O => \N__51286\,
            I => \N__51237\
        );

    \I__12210\ : Span4Mux_h
    port map (
            O => \N__51281\,
            I => \N__51237\
        );

    \I__12209\ : LocalMux
    port map (
            O => \N__51278\,
            I => adc_state_2_adj_1500
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__51275\,
            I => adc_state_2_adj_1500
        );

    \I__12207\ : Odrv4
    port map (
            O => \N__51272\,
            I => adc_state_2_adj_1500
        );

    \I__12206\ : Odrv4
    port map (
            O => \N__51269\,
            I => adc_state_2_adj_1500
        );

    \I__12205\ : LocalMux
    port map (
            O => \N__51264\,
            I => adc_state_2_adj_1500
        );

    \I__12204\ : LocalMux
    port map (
            O => \N__51257\,
            I => adc_state_2_adj_1500
        );

    \I__12203\ : Odrv4
    port map (
            O => \N__51254\,
            I => adc_state_2_adj_1500
        );

    \I__12202\ : Odrv4
    port map (
            O => \N__51251\,
            I => adc_state_2_adj_1500
        );

    \I__12201\ : Odrv4
    port map (
            O => \N__51246\,
            I => adc_state_2_adj_1500
        );

    \I__12200\ : Odrv4
    port map (
            O => \N__51237\,
            I => adc_state_2_adj_1500
        );

    \I__12199\ : CascadeMux
    port map (
            O => \N__51216\,
            I => \ADC_VDC.n52_cascade_\
        );

    \I__12198\ : InMux
    port map (
            O => \N__51213\,
            I => \N__51205\
        );

    \I__12197\ : InMux
    port map (
            O => \N__51212\,
            I => \N__51198\
        );

    \I__12196\ : InMux
    port map (
            O => \N__51211\,
            I => \N__51198\
        );

    \I__12195\ : InMux
    port map (
            O => \N__51210\,
            I => \N__51194\
        );

    \I__12194\ : InMux
    port map (
            O => \N__51209\,
            I => \N__51191\
        );

    \I__12193\ : InMux
    port map (
            O => \N__51208\,
            I => \N__51188\
        );

    \I__12192\ : LocalMux
    port map (
            O => \N__51205\,
            I => \N__51185\
        );

    \I__12191\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51181\
        );

    \I__12190\ : InMux
    port map (
            O => \N__51203\,
            I => \N__51176\
        );

    \I__12189\ : LocalMux
    port map (
            O => \N__51198\,
            I => \N__51171\
        );

    \I__12188\ : InMux
    port map (
            O => \N__51197\,
            I => \N__51168\
        );

    \I__12187\ : LocalMux
    port map (
            O => \N__51194\,
            I => \N__51163\
        );

    \I__12186\ : LocalMux
    port map (
            O => \N__51191\,
            I => \N__51163\
        );

    \I__12185\ : LocalMux
    port map (
            O => \N__51188\,
            I => \N__51158\
        );

    \I__12184\ : Span4Mux_h
    port map (
            O => \N__51185\,
            I => \N__51158\
        );

    \I__12183\ : InMux
    port map (
            O => \N__51184\,
            I => \N__51155\
        );

    \I__12182\ : LocalMux
    port map (
            O => \N__51181\,
            I => \N__51146\
        );

    \I__12181\ : InMux
    port map (
            O => \N__51180\,
            I => \N__51142\
        );

    \I__12180\ : InMux
    port map (
            O => \N__51179\,
            I => \N__51139\
        );

    \I__12179\ : LocalMux
    port map (
            O => \N__51176\,
            I => \N__51136\
        );

    \I__12178\ : InMux
    port map (
            O => \N__51175\,
            I => \N__51133\
        );

    \I__12177\ : InMux
    port map (
            O => \N__51174\,
            I => \N__51130\
        );

    \I__12176\ : Sp12to4
    port map (
            O => \N__51171\,
            I => \N__51125\
        );

    \I__12175\ : LocalMux
    port map (
            O => \N__51168\,
            I => \N__51125\
        );

    \I__12174\ : Span4Mux_v
    port map (
            O => \N__51163\,
            I => \N__51118\
        );

    \I__12173\ : Span4Mux_h
    port map (
            O => \N__51158\,
            I => \N__51118\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__51155\,
            I => \N__51118\
        );

    \I__12171\ : InMux
    port map (
            O => \N__51154\,
            I => \N__51111\
        );

    \I__12170\ : InMux
    port map (
            O => \N__51153\,
            I => \N__51111\
        );

    \I__12169\ : InMux
    port map (
            O => \N__51152\,
            I => \N__51111\
        );

    \I__12168\ : InMux
    port map (
            O => \N__51151\,
            I => \N__51104\
        );

    \I__12167\ : InMux
    port map (
            O => \N__51150\,
            I => \N__51104\
        );

    \I__12166\ : InMux
    port map (
            O => \N__51149\,
            I => \N__51104\
        );

    \I__12165\ : Span12Mux_h
    port map (
            O => \N__51146\,
            I => \N__51101\
        );

    \I__12164\ : InMux
    port map (
            O => \N__51145\,
            I => \N__51098\
        );

    \I__12163\ : LocalMux
    port map (
            O => \N__51142\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12162\ : LocalMux
    port map (
            O => \N__51139\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12161\ : Odrv4
    port map (
            O => \N__51136\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__51133\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12159\ : LocalMux
    port map (
            O => \N__51130\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12158\ : Odrv12
    port map (
            O => \N__51125\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12157\ : Odrv4
    port map (
            O => \N__51118\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__51111\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12155\ : LocalMux
    port map (
            O => \N__51104\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12154\ : Odrv12
    port map (
            O => \N__51101\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__51098\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__12152\ : CEMux
    port map (
            O => \N__51075\,
            I => \N__51072\
        );

    \I__12151\ : LocalMux
    port map (
            O => \N__51072\,
            I => \N__51069\
        );

    \I__12150\ : Span4Mux_h
    port map (
            O => \N__51069\,
            I => \N__51066\
        );

    \I__12149\ : Odrv4
    port map (
            O => \N__51066\,
            I => \ADC_VDC.n11905\
        );

    \I__12148\ : InMux
    port map (
            O => \N__51063\,
            I => \bfn_19_7_0_\
        );

    \I__12147\ : InMux
    port map (
            O => \N__51060\,
            I => \ADC_VDC.genclk.n19888\
        );

    \I__12146\ : InMux
    port map (
            O => \N__51057\,
            I => \ADC_VDC.genclk.n19889\
        );

    \I__12145\ : InMux
    port map (
            O => \N__51054\,
            I => \ADC_VDC.genclk.n19890\
        );

    \I__12144\ : InMux
    port map (
            O => \N__51051\,
            I => \ADC_VDC.genclk.n19891\
        );

    \I__12143\ : InMux
    port map (
            O => \N__51048\,
            I => \ADC_VDC.genclk.n19892\
        );

    \I__12142\ : InMux
    port map (
            O => \N__51045\,
            I => \N__51041\
        );

    \I__12141\ : InMux
    port map (
            O => \N__51044\,
            I => \N__51038\
        );

    \I__12140\ : LocalMux
    port map (
            O => \N__51041\,
            I => dds0_mclkcnt_5
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__51038\,
            I => dds0_mclkcnt_5
        );

    \I__12138\ : InMux
    port map (
            O => \N__51033\,
            I => n19929
        );

    \I__12137\ : InMux
    port map (
            O => \N__51030\,
            I => \N__51027\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__51027\,
            I => n10_adj_1528
        );

    \I__12135\ : CascadeMux
    port map (
            O => \N__51024\,
            I => \N__51021\
        );

    \I__12134\ : InMux
    port map (
            O => \N__51021\,
            I => \N__51015\
        );

    \I__12133\ : InMux
    port map (
            O => \N__51020\,
            I => \N__51015\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__51015\,
            I => dds0_mclkcnt_6
        );

    \I__12131\ : InMux
    port map (
            O => \N__51012\,
            I => n19930
        );

    \I__12130\ : InMux
    port map (
            O => \N__51009\,
            I => n19931
        );

    \I__12129\ : InMux
    port map (
            O => \N__51006\,
            I => \N__51002\
        );

    \I__12128\ : InMux
    port map (
            O => \N__51005\,
            I => \N__50999\
        );

    \I__12127\ : LocalMux
    port map (
            O => \N__51002\,
            I => dds0_mclkcnt_7
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__50999\,
            I => dds0_mclkcnt_7
        );

    \I__12125\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50991\
        );

    \I__12124\ : LocalMux
    port map (
            O => \N__50991\,
            I => \N__50987\
        );

    \I__12123\ : CascadeMux
    port map (
            O => \N__50990\,
            I => \N__50984\
        );

    \I__12122\ : Span4Mux_v
    port map (
            O => \N__50987\,
            I => \N__50977\
        );

    \I__12121\ : InMux
    port map (
            O => \N__50984\,
            I => \N__50972\
        );

    \I__12120\ : InMux
    port map (
            O => \N__50983\,
            I => \N__50972\
        );

    \I__12119\ : InMux
    port map (
            O => \N__50982\,
            I => \N__50969\
        );

    \I__12118\ : InMux
    port map (
            O => \N__50981\,
            I => \N__50966\
        );

    \I__12117\ : CascadeMux
    port map (
            O => \N__50980\,
            I => \N__50963\
        );

    \I__12116\ : Span4Mux_h
    port map (
            O => \N__50977\,
            I => \N__50960\
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__50972\,
            I => \N__50957\
        );

    \I__12114\ : LocalMux
    port map (
            O => \N__50969\,
            I => \N__50954\
        );

    \I__12113\ : LocalMux
    port map (
            O => \N__50966\,
            I => \N__50949\
        );

    \I__12112\ : InMux
    port map (
            O => \N__50963\,
            I => \N__50946\
        );

    \I__12111\ : Span4Mux_h
    port map (
            O => \N__50960\,
            I => \N__50941\
        );

    \I__12110\ : Span4Mux_v
    port map (
            O => \N__50957\,
            I => \N__50941\
        );

    \I__12109\ : Span4Mux_v
    port map (
            O => \N__50954\,
            I => \N__50938\
        );

    \I__12108\ : InMux
    port map (
            O => \N__50953\,
            I => \N__50933\
        );

    \I__12107\ : InMux
    port map (
            O => \N__50952\,
            I => \N__50933\
        );

    \I__12106\ : Span4Mux_h
    port map (
            O => \N__50949\,
            I => \N__50928\
        );

    \I__12105\ : LocalMux
    port map (
            O => \N__50946\,
            I => \N__50928\
        );

    \I__12104\ : Span4Mux_h
    port map (
            O => \N__50941\,
            I => \N__50925\
        );

    \I__12103\ : Span4Mux_h
    port map (
            O => \N__50938\,
            I => \N__50922\
        );

    \I__12102\ : LocalMux
    port map (
            O => \N__50933\,
            I => \N__50919\
        );

    \I__12101\ : Sp12to4
    port map (
            O => \N__50928\,
            I => \N__50916\
        );

    \I__12100\ : Span4Mux_v
    port map (
            O => \N__50925\,
            I => \N__50913\
        );

    \I__12099\ : Span4Mux_h
    port map (
            O => \N__50922\,
            I => \N__50908\
        );

    \I__12098\ : Span4Mux_v
    port map (
            O => \N__50919\,
            I => \N__50908\
        );

    \I__12097\ : Span12Mux_v
    port map (
            O => \N__50916\,
            I => \N__50905\
        );

    \I__12096\ : Span4Mux_h
    port map (
            O => \N__50913\,
            I => \N__50902\
        );

    \I__12095\ : Span4Mux_h
    port map (
            O => \N__50908\,
            I => \N__50899\
        );

    \I__12094\ : Odrv12
    port map (
            O => \N__50905\,
            I => n14716
        );

    \I__12093\ : Odrv4
    port map (
            O => \N__50902\,
            I => n14716
        );

    \I__12092\ : Odrv4
    port map (
            O => \N__50899\,
            I => n14716
        );

    \I__12091\ : InMux
    port map (
            O => \N__50892\,
            I => \N__50888\
        );

    \I__12090\ : InMux
    port map (
            O => \N__50891\,
            I => \N__50885\
        );

    \I__12089\ : LocalMux
    port map (
            O => \N__50888\,
            I => \N__50879\
        );

    \I__12088\ : LocalMux
    port map (
            O => \N__50885\,
            I => \N__50879\
        );

    \I__12087\ : InMux
    port map (
            O => \N__50884\,
            I => \N__50876\
        );

    \I__12086\ : Span4Mux_v
    port map (
            O => \N__50879\,
            I => \N__50870\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__50876\,
            I => \N__50870\
        );

    \I__12084\ : InMux
    port map (
            O => \N__50875\,
            I => \N__50866\
        );

    \I__12083\ : Span4Mux_v
    port map (
            O => \N__50870\,
            I => \N__50863\
        );

    \I__12082\ : InMux
    port map (
            O => \N__50869\,
            I => \N__50860\
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__50866\,
            I => \N__50857\
        );

    \I__12080\ : Span4Mux_h
    port map (
            O => \N__50863\,
            I => \N__50852\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__50860\,
            I => \N__50852\
        );

    \I__12078\ : Span4Mux_h
    port map (
            O => \N__50857\,
            I => \N__50849\
        );

    \I__12077\ : Sp12to4
    port map (
            O => \N__50852\,
            I => \N__50846\
        );

    \I__12076\ : Sp12to4
    port map (
            O => \N__50849\,
            I => \N__50843\
        );

    \I__12075\ : Span12Mux_v
    port map (
            O => \N__50846\,
            I => \N__50840\
        );

    \I__12074\ : Span12Mux_v
    port map (
            O => \N__50843\,
            I => \N__50837\
        );

    \I__12073\ : Odrv12
    port map (
            O => \N__50840\,
            I => \ICE_SPI_MOSI\
        );

    \I__12072\ : Odrv12
    port map (
            O => \N__50837\,
            I => \ICE_SPI_MOSI\
        );

    \I__12071\ : SRMux
    port map (
            O => \N__50832\,
            I => \N__50829\
        );

    \I__12070\ : LocalMux
    port map (
            O => \N__50829\,
            I => \N__50826\
        );

    \I__12069\ : Span12Mux_h
    port map (
            O => \N__50826\,
            I => \N__50823\
        );

    \I__12068\ : Odrv12
    port map (
            O => \N__50823\,
            I => \comm_spi.imosi_N_793\
        );

    \I__12067\ : SRMux
    port map (
            O => \N__50820\,
            I => \N__50817\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__50817\,
            I => \N__50814\
        );

    \I__12065\ : Odrv12
    port map (
            O => \N__50814\,
            I => \comm_spi.data_tx_7__N_810\
        );

    \I__12064\ : InMux
    port map (
            O => \N__50811\,
            I => \N__50807\
        );

    \I__12063\ : InMux
    port map (
            O => \N__50810\,
            I => \N__50804\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__50807\,
            I => \N__50800\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__50804\,
            I => \N__50778\
        );

    \I__12060\ : ClkMux
    port map (
            O => \N__50803\,
            I => \N__50733\
        );

    \I__12059\ : Glb2LocalMux
    port map (
            O => \N__50800\,
            I => \N__50733\
        );

    \I__12058\ : ClkMux
    port map (
            O => \N__50799\,
            I => \N__50733\
        );

    \I__12057\ : ClkMux
    port map (
            O => \N__50798\,
            I => \N__50733\
        );

    \I__12056\ : ClkMux
    port map (
            O => \N__50797\,
            I => \N__50733\
        );

    \I__12055\ : ClkMux
    port map (
            O => \N__50796\,
            I => \N__50733\
        );

    \I__12054\ : ClkMux
    port map (
            O => \N__50795\,
            I => \N__50733\
        );

    \I__12053\ : ClkMux
    port map (
            O => \N__50794\,
            I => \N__50733\
        );

    \I__12052\ : ClkMux
    port map (
            O => \N__50793\,
            I => \N__50733\
        );

    \I__12051\ : ClkMux
    port map (
            O => \N__50792\,
            I => \N__50733\
        );

    \I__12050\ : ClkMux
    port map (
            O => \N__50791\,
            I => \N__50733\
        );

    \I__12049\ : ClkMux
    port map (
            O => \N__50790\,
            I => \N__50733\
        );

    \I__12048\ : ClkMux
    port map (
            O => \N__50789\,
            I => \N__50733\
        );

    \I__12047\ : ClkMux
    port map (
            O => \N__50788\,
            I => \N__50733\
        );

    \I__12046\ : ClkMux
    port map (
            O => \N__50787\,
            I => \N__50733\
        );

    \I__12045\ : ClkMux
    port map (
            O => \N__50786\,
            I => \N__50733\
        );

    \I__12044\ : ClkMux
    port map (
            O => \N__50785\,
            I => \N__50733\
        );

    \I__12043\ : ClkMux
    port map (
            O => \N__50784\,
            I => \N__50733\
        );

    \I__12042\ : ClkMux
    port map (
            O => \N__50783\,
            I => \N__50733\
        );

    \I__12041\ : ClkMux
    port map (
            O => \N__50782\,
            I => \N__50733\
        );

    \I__12040\ : ClkMux
    port map (
            O => \N__50781\,
            I => \N__50733\
        );

    \I__12039\ : Glb2LocalMux
    port map (
            O => \N__50778\,
            I => \N__50733\
        );

    \I__12038\ : GlobalMux
    port map (
            O => \N__50733\,
            I => \clk_16MHz\
        );

    \I__12037\ : InMux
    port map (
            O => \N__50730\,
            I => \N__50724\
        );

    \I__12036\ : InMux
    port map (
            O => \N__50729\,
            I => \N__50724\
        );

    \I__12035\ : LocalMux
    port map (
            O => \N__50724\,
            I => dds0_mclk
        );

    \I__12034\ : InMux
    port map (
            O => \N__50721\,
            I => \N__50717\
        );

    \I__12033\ : InMux
    port map (
            O => \N__50720\,
            I => \N__50714\
        );

    \I__12032\ : LocalMux
    port map (
            O => \N__50717\,
            I => \N__50711\
        );

    \I__12031\ : LocalMux
    port map (
            O => \N__50714\,
            I => \N__50707\
        );

    \I__12030\ : Span4Mux_v
    port map (
            O => \N__50711\,
            I => \N__50704\
        );

    \I__12029\ : InMux
    port map (
            O => \N__50710\,
            I => \N__50701\
        );

    \I__12028\ : Span12Mux_v
    port map (
            O => \N__50707\,
            I => \N__50698\
        );

    \I__12027\ : Odrv4
    port map (
            O => \N__50704\,
            I => buf_control_6
        );

    \I__12026\ : LocalMux
    port map (
            O => \N__50701\,
            I => buf_control_6
        );

    \I__12025\ : Odrv12
    port map (
            O => \N__50698\,
            I => buf_control_6
        );

    \I__12024\ : IoInMux
    port map (
            O => \N__50691\,
            I => \N__50688\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__50688\,
            I => \N__50685\
        );

    \I__12022\ : Span4Mux_s3_v
    port map (
            O => \N__50685\,
            I => \N__50682\
        );

    \I__12021\ : Span4Mux_h
    port map (
            O => \N__50682\,
            I => \N__50679\
        );

    \I__12020\ : Span4Mux_v
    port map (
            O => \N__50679\,
            I => \N__50676\
        );

    \I__12019\ : Span4Mux_v
    port map (
            O => \N__50676\,
            I => \N__50673\
        );

    \I__12018\ : Odrv4
    port map (
            O => \N__50673\,
            I => \DDS_MCLK\
        );

    \I__12017\ : InMux
    port map (
            O => \N__50670\,
            I => \N__50667\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__50667\,
            I => \N__50664\
        );

    \I__12015\ : Span4Mux_v
    port map (
            O => \N__50664\,
            I => \N__50660\
        );

    \I__12014\ : InMux
    port map (
            O => \N__50663\,
            I => \N__50657\
        );

    \I__12013\ : Span4Mux_h
    port map (
            O => \N__50660\,
            I => \N__50654\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__50657\,
            I => acadc_skipcnt_10
        );

    \I__12011\ : Odrv4
    port map (
            O => \N__50654\,
            I => acadc_skipcnt_10
        );

    \I__12010\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50645\
        );

    \I__12009\ : InMux
    port map (
            O => \N__50648\,
            I => \N__50641\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__50645\,
            I => \N__50638\
        );

    \I__12007\ : InMux
    port map (
            O => \N__50644\,
            I => \N__50635\
        );

    \I__12006\ : LocalMux
    port map (
            O => \N__50641\,
            I => \acadc_skipCount_12\
        );

    \I__12005\ : Odrv4
    port map (
            O => \N__50638\,
            I => \acadc_skipCount_12\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__50635\,
            I => \acadc_skipCount_12\
        );

    \I__12003\ : CascadeMux
    port map (
            O => \N__50628\,
            I => \N__50625\
        );

    \I__12002\ : InMux
    port map (
            O => \N__50625\,
            I => \N__50622\
        );

    \I__12001\ : LocalMux
    port map (
            O => \N__50622\,
            I => \N__50618\
        );

    \I__12000\ : InMux
    port map (
            O => \N__50621\,
            I => \N__50615\
        );

    \I__11999\ : Span12Mux_v
    port map (
            O => \N__50618\,
            I => \N__50612\
        );

    \I__11998\ : LocalMux
    port map (
            O => \N__50615\,
            I => acadc_skipcnt_12
        );

    \I__11997\ : Odrv12
    port map (
            O => \N__50612\,
            I => acadc_skipcnt_12
        );

    \I__11996\ : InMux
    port map (
            O => \N__50607\,
            I => \N__50600\
        );

    \I__11995\ : InMux
    port map (
            O => \N__50606\,
            I => \N__50600\
        );

    \I__11994\ : InMux
    port map (
            O => \N__50605\,
            I => \N__50597\
        );

    \I__11993\ : LocalMux
    port map (
            O => \N__50600\,
            I => \acadc_skipCount_10\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__50597\,
            I => \acadc_skipCount_10\
        );

    \I__11991\ : InMux
    port map (
            O => \N__50592\,
            I => \N__50589\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__50589\,
            I => \N__50586\
        );

    \I__11989\ : Span4Mux_h
    port map (
            O => \N__50586\,
            I => \N__50583\
        );

    \I__11988\ : Odrv4
    port map (
            O => \N__50583\,
            I => n21
        );

    \I__11987\ : CEMux
    port map (
            O => \N__50580\,
            I => \N__50577\
        );

    \I__11986\ : LocalMux
    port map (
            O => \N__50577\,
            I => \N__50574\
        );

    \I__11985\ : Span4Mux_v
    port map (
            O => \N__50574\,
            I => \N__50571\
        );

    \I__11984\ : Odrv4
    port map (
            O => \N__50571\,
            I => n11590
        );

    \I__11983\ : InMux
    port map (
            O => \N__50568\,
            I => \N__50564\
        );

    \I__11982\ : InMux
    port map (
            O => \N__50567\,
            I => \N__50561\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__50564\,
            I => dds0_mclkcnt_0
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__50561\,
            I => dds0_mclkcnt_0
        );

    \I__11979\ : InMux
    port map (
            O => \N__50556\,
            I => \bfn_18_16_0_\
        );

    \I__11978\ : CascadeMux
    port map (
            O => \N__50553\,
            I => \N__50549\
        );

    \I__11977\ : InMux
    port map (
            O => \N__50552\,
            I => \N__50546\
        );

    \I__11976\ : InMux
    port map (
            O => \N__50549\,
            I => \N__50543\
        );

    \I__11975\ : LocalMux
    port map (
            O => \N__50546\,
            I => dds0_mclkcnt_1
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__50543\,
            I => dds0_mclkcnt_1
        );

    \I__11973\ : InMux
    port map (
            O => \N__50538\,
            I => n19925
        );

    \I__11972\ : CascadeMux
    port map (
            O => \N__50535\,
            I => \N__50531\
        );

    \I__11971\ : InMux
    port map (
            O => \N__50534\,
            I => \N__50528\
        );

    \I__11970\ : InMux
    port map (
            O => \N__50531\,
            I => \N__50525\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__50528\,
            I => dds0_mclkcnt_2
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__50525\,
            I => dds0_mclkcnt_2
        );

    \I__11967\ : InMux
    port map (
            O => \N__50520\,
            I => n19926
        );

    \I__11966\ : InMux
    port map (
            O => \N__50517\,
            I => \N__50513\
        );

    \I__11965\ : InMux
    port map (
            O => \N__50516\,
            I => \N__50510\
        );

    \I__11964\ : LocalMux
    port map (
            O => \N__50513\,
            I => dds0_mclkcnt_3
        );

    \I__11963\ : LocalMux
    port map (
            O => \N__50510\,
            I => dds0_mclkcnt_3
        );

    \I__11962\ : InMux
    port map (
            O => \N__50505\,
            I => n19927
        );

    \I__11961\ : InMux
    port map (
            O => \N__50502\,
            I => \N__50498\
        );

    \I__11960\ : InMux
    port map (
            O => \N__50501\,
            I => \N__50495\
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__50498\,
            I => dds0_mclkcnt_4
        );

    \I__11958\ : LocalMux
    port map (
            O => \N__50495\,
            I => dds0_mclkcnt_4
        );

    \I__11957\ : InMux
    port map (
            O => \N__50490\,
            I => n19928
        );

    \I__11956\ : InMux
    port map (
            O => \N__50487\,
            I => \N__50484\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__50484\,
            I => \N__50481\
        );

    \I__11954\ : Odrv4
    port map (
            O => \N__50481\,
            I => n4_adj_1581
        );

    \I__11953\ : CascadeMux
    port map (
            O => \N__50478\,
            I => \n21282_cascade_\
        );

    \I__11952\ : InMux
    port map (
            O => \N__50475\,
            I => \N__50472\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__50472\,
            I => \N__50469\
        );

    \I__11950\ : Odrv4
    port map (
            O => \N__50469\,
            I => n22548
        );

    \I__11949\ : InMux
    port map (
            O => \N__50466\,
            I => \N__50463\
        );

    \I__11948\ : LocalMux
    port map (
            O => \N__50463\,
            I => \N__50459\
        );

    \I__11947\ : InMux
    port map (
            O => \N__50462\,
            I => \N__50456\
        );

    \I__11946\ : Span4Mux_v
    port map (
            O => \N__50459\,
            I => \N__50450\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__50456\,
            I => \N__50450\
        );

    \I__11944\ : InMux
    port map (
            O => \N__50455\,
            I => \N__50447\
        );

    \I__11943\ : Span4Mux_v
    port map (
            O => \N__50450\,
            I => \N__50442\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__50447\,
            I => \N__50442\
        );

    \I__11941\ : Span4Mux_v
    port map (
            O => \N__50442\,
            I => \N__50439\
        );

    \I__11940\ : Span4Mux_h
    port map (
            O => \N__50439\,
            I => \N__50436\
        );

    \I__11939\ : Odrv4
    port map (
            O => \N__50436\,
            I => comm_tx_buf_6
        );

    \I__11938\ : InMux
    port map (
            O => \N__50433\,
            I => \N__50430\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__50430\,
            I => \N__50427\
        );

    \I__11936\ : Odrv12
    port map (
            O => \N__50427\,
            I => comm_buf_5_5
        );

    \I__11935\ : CascadeMux
    port map (
            O => \N__50424\,
            I => \N__50419\
        );

    \I__11934\ : InMux
    port map (
            O => \N__50423\,
            I => \N__50415\
        );

    \I__11933\ : InMux
    port map (
            O => \N__50422\,
            I => \N__50411\
        );

    \I__11932\ : InMux
    port map (
            O => \N__50419\,
            I => \N__50406\
        );

    \I__11931\ : InMux
    port map (
            O => \N__50418\,
            I => \N__50406\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__50415\,
            I => \N__50403\
        );

    \I__11929\ : InMux
    port map (
            O => \N__50414\,
            I => \N__50400\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__50411\,
            I => \N__50397\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__50406\,
            I => \N__50394\
        );

    \I__11926\ : Span4Mux_v
    port map (
            O => \N__50403\,
            I => \N__50391\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__50400\,
            I => \N__50388\
        );

    \I__11924\ : Span4Mux_h
    port map (
            O => \N__50397\,
            I => \N__50385\
        );

    \I__11923\ : Span4Mux_v
    port map (
            O => \N__50394\,
            I => \N__50382\
        );

    \I__11922\ : Span4Mux_h
    port map (
            O => \N__50391\,
            I => \N__50375\
        );

    \I__11921\ : Span4Mux_v
    port map (
            O => \N__50388\,
            I => \N__50375\
        );

    \I__11920\ : Span4Mux_v
    port map (
            O => \N__50385\,
            I => \N__50375\
        );

    \I__11919\ : Odrv4
    port map (
            O => \N__50382\,
            I => comm_buf_1_5
        );

    \I__11918\ : Odrv4
    port map (
            O => \N__50375\,
            I => comm_buf_1_5
        );

    \I__11917\ : InMux
    port map (
            O => \N__50370\,
            I => \N__50367\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__50367\,
            I => \N__50364\
        );

    \I__11915\ : Odrv4
    port map (
            O => \N__50364\,
            I => comm_buf_3_5
        );

    \I__11914\ : CascadeMux
    port map (
            O => \N__50361\,
            I => \n17698_cascade_\
        );

    \I__11913\ : CascadeMux
    port map (
            O => \N__50358\,
            I => \n21270_cascade_\
        );

    \I__11912\ : CEMux
    port map (
            O => \N__50355\,
            I => \N__50351\
        );

    \I__11911\ : CEMux
    port map (
            O => \N__50354\,
            I => \N__50348\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__50351\,
            I => \N__50343\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__50348\,
            I => \N__50343\
        );

    \I__11908\ : Span4Mux_v
    port map (
            O => \N__50343\,
            I => \N__50338\
        );

    \I__11907\ : CEMux
    port map (
            O => \N__50342\,
            I => \N__50335\
        );

    \I__11906\ : CEMux
    port map (
            O => \N__50341\,
            I => \N__50330\
        );

    \I__11905\ : Span4Mux_h
    port map (
            O => \N__50338\,
            I => \N__50325\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__50335\,
            I => \N__50325\
        );

    \I__11903\ : CEMux
    port map (
            O => \N__50334\,
            I => \N__50322\
        );

    \I__11902\ : CEMux
    port map (
            O => \N__50333\,
            I => \N__50318\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__50330\,
            I => \N__50315\
        );

    \I__11900\ : Span4Mux_h
    port map (
            O => \N__50325\,
            I => \N__50312\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__50322\,
            I => \N__50309\
        );

    \I__11898\ : InMux
    port map (
            O => \N__50321\,
            I => \N__50306\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__50318\,
            I => \N__50302\
        );

    \I__11896\ : Span4Mux_h
    port map (
            O => \N__50315\,
            I => \N__50299\
        );

    \I__11895\ : Sp12to4
    port map (
            O => \N__50312\,
            I => \N__50296\
        );

    \I__11894\ : Span4Mux_v
    port map (
            O => \N__50309\,
            I => \N__50291\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__50306\,
            I => \N__50291\
        );

    \I__11892\ : CEMux
    port map (
            O => \N__50305\,
            I => \N__50288\
        );

    \I__11891\ : Span12Mux_h
    port map (
            O => \N__50302\,
            I => \N__50285\
        );

    \I__11890\ : Span4Mux_v
    port map (
            O => \N__50299\,
            I => \N__50282\
        );

    \I__11889\ : Span12Mux_v
    port map (
            O => \N__50296\,
            I => \N__50279\
        );

    \I__11888\ : Span4Mux_h
    port map (
            O => \N__50291\,
            I => \N__50276\
        );

    \I__11887\ : LocalMux
    port map (
            O => \N__50288\,
            I => n12541
        );

    \I__11886\ : Odrv12
    port map (
            O => \N__50285\,
            I => n12541
        );

    \I__11885\ : Odrv4
    port map (
            O => \N__50282\,
            I => n12541
        );

    \I__11884\ : Odrv12
    port map (
            O => \N__50279\,
            I => n12541
        );

    \I__11883\ : Odrv4
    port map (
            O => \N__50276\,
            I => n12541
        );

    \I__11882\ : SRMux
    port map (
            O => \N__50265\,
            I => \N__50262\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__50262\,
            I => \N__50258\
        );

    \I__11880\ : SRMux
    port map (
            O => \N__50261\,
            I => \N__50255\
        );

    \I__11879\ : Span4Mux_h
    port map (
            O => \N__50258\,
            I => \N__50251\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__50255\,
            I => \N__50247\
        );

    \I__11877\ : SRMux
    port map (
            O => \N__50254\,
            I => \N__50244\
        );

    \I__11876\ : Span4Mux_h
    port map (
            O => \N__50251\,
            I => \N__50240\
        );

    \I__11875\ : SRMux
    port map (
            O => \N__50250\,
            I => \N__50237\
        );

    \I__11874\ : Span4Mux_h
    port map (
            O => \N__50247\,
            I => \N__50232\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__50244\,
            I => \N__50232\
        );

    \I__11872\ : SRMux
    port map (
            O => \N__50243\,
            I => \N__50228\
        );

    \I__11871\ : Span4Mux_v
    port map (
            O => \N__50240\,
            I => \N__50224\
        );

    \I__11870\ : LocalMux
    port map (
            O => \N__50237\,
            I => \N__50219\
        );

    \I__11869\ : Span4Mux_v
    port map (
            O => \N__50232\,
            I => \N__50219\
        );

    \I__11868\ : SRMux
    port map (
            O => \N__50231\,
            I => \N__50216\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__50228\,
            I => \N__50213\
        );

    \I__11866\ : SRMux
    port map (
            O => \N__50227\,
            I => \N__50210\
        );

    \I__11865\ : Sp12to4
    port map (
            O => \N__50224\,
            I => \N__50207\
        );

    \I__11864\ : Span4Mux_v
    port map (
            O => \N__50219\,
            I => \N__50204\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__50216\,
            I => \N__50201\
        );

    \I__11862\ : Span4Mux_h
    port map (
            O => \N__50213\,
            I => \N__50198\
        );

    \I__11861\ : LocalMux
    port map (
            O => \N__50210\,
            I => \N__50191\
        );

    \I__11860\ : Span12Mux_s10_h
    port map (
            O => \N__50207\,
            I => \N__50191\
        );

    \I__11859\ : Sp12to4
    port map (
            O => \N__50204\,
            I => \N__50191\
        );

    \I__11858\ : Odrv12
    port map (
            O => \N__50201\,
            I => n15007
        );

    \I__11857\ : Odrv4
    port map (
            O => \N__50198\,
            I => n15007
        );

    \I__11856\ : Odrv12
    port map (
            O => \N__50191\,
            I => n15007
        );

    \I__11855\ : CascadeMux
    port map (
            O => \N__50184\,
            I => \n20996_cascade_\
        );

    \I__11854\ : InMux
    port map (
            O => \N__50181\,
            I => \N__50178\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__50178\,
            I => n12_adj_1663
        );

    \I__11852\ : InMux
    port map (
            O => \N__50175\,
            I => \N__50172\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__50172\,
            I => n20996
        );

    \I__11850\ : CascadeMux
    port map (
            O => \N__50169\,
            I => \N__50166\
        );

    \I__11849\ : InMux
    port map (
            O => \N__50166\,
            I => \N__50162\
        );

    \I__11848\ : InMux
    port map (
            O => \N__50165\,
            I => \N__50159\
        );

    \I__11847\ : LocalMux
    port map (
            O => \N__50162\,
            I => \N__50153\
        );

    \I__11846\ : LocalMux
    port map (
            O => \N__50159\,
            I => \N__50150\
        );

    \I__11845\ : InMux
    port map (
            O => \N__50158\,
            I => \N__50147\
        );

    \I__11844\ : InMux
    port map (
            O => \N__50157\,
            I => \N__50142\
        );

    \I__11843\ : InMux
    port map (
            O => \N__50156\,
            I => \N__50139\
        );

    \I__11842\ : Span4Mux_v
    port map (
            O => \N__50153\,
            I => \N__50136\
        );

    \I__11841\ : Span4Mux_h
    port map (
            O => \N__50150\,
            I => \N__50131\
        );

    \I__11840\ : LocalMux
    port map (
            O => \N__50147\,
            I => \N__50131\
        );

    \I__11839\ : InMux
    port map (
            O => \N__50146\,
            I => \N__50128\
        );

    \I__11838\ : InMux
    port map (
            O => \N__50145\,
            I => \N__50125\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__50142\,
            I => \N__50122\
        );

    \I__11836\ : LocalMux
    port map (
            O => \N__50139\,
            I => \N__50119\
        );

    \I__11835\ : Span4Mux_h
    port map (
            O => \N__50136\,
            I => \N__50114\
        );

    \I__11834\ : Span4Mux_v
    port map (
            O => \N__50131\,
            I => \N__50114\
        );

    \I__11833\ : LocalMux
    port map (
            O => \N__50128\,
            I => \N__50109\
        );

    \I__11832\ : LocalMux
    port map (
            O => \N__50125\,
            I => \N__50109\
        );

    \I__11831\ : Span4Mux_v
    port map (
            O => \N__50122\,
            I => \N__50105\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__50119\,
            I => \N__50098\
        );

    \I__11829\ : Span4Mux_h
    port map (
            O => \N__50114\,
            I => \N__50098\
        );

    \I__11828\ : Span4Mux_v
    port map (
            O => \N__50109\,
            I => \N__50098\
        );

    \I__11827\ : InMux
    port map (
            O => \N__50108\,
            I => \N__50095\
        );

    \I__11826\ : Span4Mux_h
    port map (
            O => \N__50105\,
            I => \N__50091\
        );

    \I__11825\ : Sp12to4
    port map (
            O => \N__50098\,
            I => \N__50088\
        );

    \I__11824\ : LocalMux
    port map (
            O => \N__50095\,
            I => \N__50085\
        );

    \I__11823\ : InMux
    port map (
            O => \N__50094\,
            I => \N__50082\
        );

    \I__11822\ : Odrv4
    port map (
            O => \N__50091\,
            I => comm_rx_buf_2
        );

    \I__11821\ : Odrv12
    port map (
            O => \N__50088\,
            I => comm_rx_buf_2
        );

    \I__11820\ : Odrv12
    port map (
            O => \N__50085\,
            I => comm_rx_buf_2
        );

    \I__11819\ : LocalMux
    port map (
            O => \N__50082\,
            I => comm_rx_buf_2
        );

    \I__11818\ : InMux
    port map (
            O => \N__50073\,
            I => \N__50069\
        );

    \I__11817\ : InMux
    port map (
            O => \N__50072\,
            I => \N__50066\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__50069\,
            I => comm_buf_6_2
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__50066\,
            I => comm_buf_6_2
        );

    \I__11814\ : InMux
    port map (
            O => \N__50061\,
            I => \N__50058\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__50058\,
            I => \N__50055\
        );

    \I__11812\ : Span4Mux_v
    port map (
            O => \N__50055\,
            I => \N__50052\
        );

    \I__11811\ : Odrv4
    port map (
            O => \N__50052\,
            I => comm_buf_5_0
        );

    \I__11810\ : InMux
    port map (
            O => \N__50049\,
            I => \N__50046\
        );

    \I__11809\ : LocalMux
    port map (
            O => \N__50046\,
            I => \N__50043\
        );

    \I__11808\ : Span4Mux_v
    port map (
            O => \N__50043\,
            I => \N__50040\
        );

    \I__11807\ : Odrv4
    port map (
            O => \N__50040\,
            I => comm_buf_4_0
        );

    \I__11806\ : InMux
    port map (
            O => \N__50037\,
            I => \N__50034\
        );

    \I__11805\ : LocalMux
    port map (
            O => \N__50034\,
            I => n4_adj_1457
        );

    \I__11804\ : InMux
    port map (
            O => \N__50031\,
            I => \N__50028\
        );

    \I__11803\ : LocalMux
    port map (
            O => \N__50028\,
            I => \N__50025\
        );

    \I__11802\ : Span4Mux_v
    port map (
            O => \N__50025\,
            I => \N__50022\
        );

    \I__11801\ : Odrv4
    port map (
            O => \N__50022\,
            I => comm_buf_5_1
        );

    \I__11800\ : InMux
    port map (
            O => \N__50019\,
            I => \N__50016\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__50016\,
            I => \N__50013\
        );

    \I__11798\ : Span4Mux_v
    port map (
            O => \N__50013\,
            I => \N__50010\
        );

    \I__11797\ : Odrv4
    port map (
            O => \N__50010\,
            I => comm_buf_4_1
        );

    \I__11796\ : InMux
    port map (
            O => \N__50007\,
            I => \N__50004\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__50004\,
            I => \N__49999\
        );

    \I__11794\ : InMux
    port map (
            O => \N__50003\,
            I => \N__49994\
        );

    \I__11793\ : InMux
    port map (
            O => \N__50002\,
            I => \N__49994\
        );

    \I__11792\ : Span4Mux_v
    port map (
            O => \N__49999\,
            I => \N__49988\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__49994\,
            I => \N__49988\
        );

    \I__11790\ : InMux
    port map (
            O => \N__49993\,
            I => \N__49985\
        );

    \I__11789\ : Span4Mux_h
    port map (
            O => \N__49988\,
            I => \N__49982\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__49985\,
            I => comm_cmd_7
        );

    \I__11787\ : Odrv4
    port map (
            O => \N__49982\,
            I => comm_cmd_7
        );

    \I__11786\ : InMux
    port map (
            O => \N__49977\,
            I => \N__49974\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__49974\,
            I => \N__49970\
        );

    \I__11784\ : InMux
    port map (
            O => \N__49973\,
            I => \N__49967\
        );

    \I__11783\ : Span12Mux_h
    port map (
            O => \N__49970\,
            I => \N__49964\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__49967\,
            I => comm_buf_6_1
        );

    \I__11781\ : Odrv12
    port map (
            O => \N__49964\,
            I => comm_buf_6_1
        );

    \I__11780\ : InMux
    port map (
            O => \N__49959\,
            I => \N__49956\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__49956\,
            I => n4_adj_1588
        );

    \I__11778\ : CascadeMux
    port map (
            O => \N__49953\,
            I => \n21433_cascade_\
        );

    \I__11777\ : CascadeMux
    port map (
            O => \N__49950\,
            I => \n22419_cascade_\
        );

    \I__11776\ : InMux
    port map (
            O => \N__49947\,
            I => \N__49944\
        );

    \I__11775\ : LocalMux
    port map (
            O => \N__49944\,
            I => \N__49939\
        );

    \I__11774\ : InMux
    port map (
            O => \N__49943\,
            I => \N__49936\
        );

    \I__11773\ : InMux
    port map (
            O => \N__49942\,
            I => \N__49933\
        );

    \I__11772\ : Span4Mux_v
    port map (
            O => \N__49939\,
            I => \N__49928\
        );

    \I__11771\ : LocalMux
    port map (
            O => \N__49936\,
            I => \N__49923\
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__49933\,
            I => \N__49923\
        );

    \I__11769\ : InMux
    port map (
            O => \N__49932\,
            I => \N__49920\
        );

    \I__11768\ : InMux
    port map (
            O => \N__49931\,
            I => \N__49917\
        );

    \I__11767\ : Odrv4
    port map (
            O => \N__49928\,
            I => n21085
        );

    \I__11766\ : Odrv4
    port map (
            O => \N__49923\,
            I => n21085
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__49920\,
            I => n21085
        );

    \I__11764\ : LocalMux
    port map (
            O => \N__49917\,
            I => n21085
        );

    \I__11763\ : CascadeMux
    port map (
            O => \N__49908\,
            I => \n7_adj_1458_cascade_\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49905\,
            I => \N__49902\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__49902\,
            I => \N__49899\
        );

    \I__11760\ : Span4Mux_h
    port map (
            O => \N__49899\,
            I => \N__49896\
        );

    \I__11759\ : Span4Mux_v
    port map (
            O => \N__49896\,
            I => \N__49893\
        );

    \I__11758\ : Odrv4
    port map (
            O => \N__49893\,
            I => buf_data_vac_20
        );

    \I__11757\ : InMux
    port map (
            O => \N__49890\,
            I => \N__49887\
        );

    \I__11756\ : LocalMux
    port map (
            O => \N__49887\,
            I => \N__49884\
        );

    \I__11755\ : Span4Mux_h
    port map (
            O => \N__49884\,
            I => \N__49881\
        );

    \I__11754\ : Odrv4
    port map (
            O => \N__49881\,
            I => comm_buf_3_4
        );

    \I__11753\ : InMux
    port map (
            O => \N__49878\,
            I => \N__49872\
        );

    \I__11752\ : InMux
    port map (
            O => \N__49877\,
            I => \N__49869\
        );

    \I__11751\ : InMux
    port map (
            O => \N__49876\,
            I => \N__49864\
        );

    \I__11750\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49861\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__49872\,
            I => \N__49857\
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__49869\,
            I => \N__49853\
        );

    \I__11747\ : InMux
    port map (
            O => \N__49868\,
            I => \N__49850\
        );

    \I__11746\ : InMux
    port map (
            O => \N__49867\,
            I => \N__49847\
        );

    \I__11745\ : LocalMux
    port map (
            O => \N__49864\,
            I => \N__49844\
        );

    \I__11744\ : LocalMux
    port map (
            O => \N__49861\,
            I => \N__49841\
        );

    \I__11743\ : InMux
    port map (
            O => \N__49860\,
            I => \N__49838\
        );

    \I__11742\ : Span4Mux_v
    port map (
            O => \N__49857\,
            I => \N__49835\
        );

    \I__11741\ : InMux
    port map (
            O => \N__49856\,
            I => \N__49832\
        );

    \I__11740\ : Span4Mux_v
    port map (
            O => \N__49853\,
            I => \N__49827\
        );

    \I__11739\ : LocalMux
    port map (
            O => \N__49850\,
            I => \N__49827\
        );

    \I__11738\ : LocalMux
    port map (
            O => \N__49847\,
            I => \N__49824\
        );

    \I__11737\ : Span4Mux_h
    port map (
            O => \N__49844\,
            I => \N__49821\
        );

    \I__11736\ : Span4Mux_h
    port map (
            O => \N__49841\,
            I => \N__49816\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__49838\,
            I => \N__49816\
        );

    \I__11734\ : Span4Mux_h
    port map (
            O => \N__49835\,
            I => \N__49811\
        );

    \I__11733\ : LocalMux
    port map (
            O => \N__49832\,
            I => \N__49811\
        );

    \I__11732\ : Span4Mux_v
    port map (
            O => \N__49827\,
            I => \N__49805\
        );

    \I__11731\ : Span4Mux_v
    port map (
            O => \N__49824\,
            I => \N__49805\
        );

    \I__11730\ : Span4Mux_h
    port map (
            O => \N__49821\,
            I => \N__49798\
        );

    \I__11729\ : Span4Mux_v
    port map (
            O => \N__49816\,
            I => \N__49798\
        );

    \I__11728\ : Span4Mux_h
    port map (
            O => \N__49811\,
            I => \N__49798\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49810\,
            I => \N__49795\
        );

    \I__11726\ : Odrv4
    port map (
            O => \N__49805\,
            I => comm_rx_buf_3
        );

    \I__11725\ : Odrv4
    port map (
            O => \N__49798\,
            I => comm_rx_buf_3
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__49795\,
            I => comm_rx_buf_3
        );

    \I__11723\ : InMux
    port map (
            O => \N__49788\,
            I => \N__49785\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__49785\,
            I => \N__49782\
        );

    \I__11721\ : Span4Mux_v
    port map (
            O => \N__49782\,
            I => \N__49779\
        );

    \I__11720\ : Odrv4
    port map (
            O => \N__49779\,
            I => buf_data_vac_19
        );

    \I__11719\ : CascadeMux
    port map (
            O => \N__49776\,
            I => \N__49773\
        );

    \I__11718\ : InMux
    port map (
            O => \N__49773\,
            I => \N__49770\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__49770\,
            I => comm_buf_3_3
        );

    \I__11716\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49764\
        );

    \I__11715\ : LocalMux
    port map (
            O => \N__49764\,
            I => \N__49761\
        );

    \I__11714\ : Span4Mux_h
    port map (
            O => \N__49761\,
            I => \N__49758\
        );

    \I__11713\ : Odrv4
    port map (
            O => \N__49758\,
            I => buf_data_vac_18
        );

    \I__11712\ : CascadeMux
    port map (
            O => \N__49755\,
            I => \N__49752\
        );

    \I__11711\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49749\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__49749\,
            I => comm_buf_3_2
        );

    \I__11709\ : CascadeMux
    port map (
            O => \N__49746\,
            I => \N__49742\
        );

    \I__11708\ : CascadeMux
    port map (
            O => \N__49745\,
            I => \N__49739\
        );

    \I__11707\ : InMux
    port map (
            O => \N__49742\,
            I => \N__49736\
        );

    \I__11706\ : InMux
    port map (
            O => \N__49739\,
            I => \N__49733\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__49736\,
            I => \N__49730\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__49733\,
            I => \N__49727\
        );

    \I__11703\ : Span4Mux_h
    port map (
            O => \N__49730\,
            I => \N__49724\
        );

    \I__11702\ : Span4Mux_v
    port map (
            O => \N__49727\,
            I => \N__49718\
        );

    \I__11701\ : Span4Mux_h
    port map (
            O => \N__49724\,
            I => \N__49714\
        );

    \I__11700\ : InMux
    port map (
            O => \N__49723\,
            I => \N__49711\
        );

    \I__11699\ : InMux
    port map (
            O => \N__49722\,
            I => \N__49708\
        );

    \I__11698\ : InMux
    port map (
            O => \N__49721\,
            I => \N__49705\
        );

    \I__11697\ : Span4Mux_h
    port map (
            O => \N__49718\,
            I => \N__49701\
        );

    \I__11696\ : InMux
    port map (
            O => \N__49717\,
            I => \N__49698\
        );

    \I__11695\ : Span4Mux_h
    port map (
            O => \N__49714\,
            I => \N__49693\
        );

    \I__11694\ : LocalMux
    port map (
            O => \N__49711\,
            I => \N__49693\
        );

    \I__11693\ : LocalMux
    port map (
            O => \N__49708\,
            I => \N__49690\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__49705\,
            I => \N__49687\
        );

    \I__11691\ : InMux
    port map (
            O => \N__49704\,
            I => \N__49684\
        );

    \I__11690\ : Span4Mux_h
    port map (
            O => \N__49701\,
            I => \N__49679\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__49698\,
            I => \N__49679\
        );

    \I__11688\ : Span4Mux_v
    port map (
            O => \N__49693\,
            I => \N__49675\
        );

    \I__11687\ : Span4Mux_h
    port map (
            O => \N__49690\,
            I => \N__49672\
        );

    \I__11686\ : Span4Mux_h
    port map (
            O => \N__49687\,
            I => \N__49669\
        );

    \I__11685\ : LocalMux
    port map (
            O => \N__49684\,
            I => \N__49666\
        );

    \I__11684\ : Span4Mux_h
    port map (
            O => \N__49679\,
            I => \N__49663\
        );

    \I__11683\ : InMux
    port map (
            O => \N__49678\,
            I => \N__49660\
        );

    \I__11682\ : Sp12to4
    port map (
            O => \N__49675\,
            I => \N__49656\
        );

    \I__11681\ : Span4Mux_v
    port map (
            O => \N__49672\,
            I => \N__49649\
        );

    \I__11680\ : Span4Mux_h
    port map (
            O => \N__49669\,
            I => \N__49649\
        );

    \I__11679\ : Span4Mux_h
    port map (
            O => \N__49666\,
            I => \N__49649\
        );

    \I__11678\ : Span4Mux_v
    port map (
            O => \N__49663\,
            I => \N__49644\
        );

    \I__11677\ : LocalMux
    port map (
            O => \N__49660\,
            I => \N__49644\
        );

    \I__11676\ : InMux
    port map (
            O => \N__49659\,
            I => \N__49641\
        );

    \I__11675\ : Odrv12
    port map (
            O => \N__49656\,
            I => comm_rx_buf_1
        );

    \I__11674\ : Odrv4
    port map (
            O => \N__49649\,
            I => comm_rx_buf_1
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__49644\,
            I => comm_rx_buf_1
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__49641\,
            I => comm_rx_buf_1
        );

    \I__11671\ : InMux
    port map (
            O => \N__49632\,
            I => \N__49629\
        );

    \I__11670\ : LocalMux
    port map (
            O => \N__49629\,
            I => \N__49626\
        );

    \I__11669\ : Odrv12
    port map (
            O => \N__49626\,
            I => buf_data_vac_17
        );

    \I__11668\ : InMux
    port map (
            O => \N__49623\,
            I => \N__49620\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__49620\,
            I => \N__49617\
        );

    \I__11666\ : Odrv12
    port map (
            O => \N__49617\,
            I => comm_buf_5_6
        );

    \I__11665\ : InMux
    port map (
            O => \N__49614\,
            I => \N__49611\
        );

    \I__11664\ : LocalMux
    port map (
            O => \N__49611\,
            I => \N__49608\
        );

    \I__11663\ : Span4Mux_v
    port map (
            O => \N__49608\,
            I => \N__49605\
        );

    \I__11662\ : Odrv4
    port map (
            O => \N__49605\,
            I => comm_buf_4_6
        );

    \I__11661\ : InMux
    port map (
            O => \N__49602\,
            I => \N__49599\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__49599\,
            I => comm_buf_2_6
        );

    \I__11659\ : CascadeMux
    port map (
            O => \N__49596\,
            I => \N__49593\
        );

    \I__11658\ : InMux
    port map (
            O => \N__49593\,
            I => \N__49590\
        );

    \I__11657\ : LocalMux
    port map (
            O => \N__49590\,
            I => comm_buf_3_6
        );

    \I__11656\ : CascadeMux
    port map (
            O => \N__49587\,
            I => \N__49582\
        );

    \I__11655\ : CascadeMux
    port map (
            O => \N__49586\,
            I => \N__49579\
        );

    \I__11654\ : CascadeMux
    port map (
            O => \N__49585\,
            I => \N__49576\
        );

    \I__11653\ : InMux
    port map (
            O => \N__49582\,
            I => \N__49573\
        );

    \I__11652\ : InMux
    port map (
            O => \N__49579\,
            I => \N__49570\
        );

    \I__11651\ : InMux
    port map (
            O => \N__49576\,
            I => \N__49564\
        );

    \I__11650\ : LocalMux
    port map (
            O => \N__49573\,
            I => \N__49561\
        );

    \I__11649\ : LocalMux
    port map (
            O => \N__49570\,
            I => \N__49558\
        );

    \I__11648\ : CascadeMux
    port map (
            O => \N__49569\,
            I => \N__49554\
        );

    \I__11647\ : InMux
    port map (
            O => \N__49568\,
            I => \N__49549\
        );

    \I__11646\ : InMux
    port map (
            O => \N__49567\,
            I => \N__49549\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__49564\,
            I => \N__49546\
        );

    \I__11644\ : Span4Mux_v
    port map (
            O => \N__49561\,
            I => \N__49541\
        );

    \I__11643\ : Span4Mux_v
    port map (
            O => \N__49558\,
            I => \N__49541\
        );

    \I__11642\ : InMux
    port map (
            O => \N__49557\,
            I => \N__49538\
        );

    \I__11641\ : InMux
    port map (
            O => \N__49554\,
            I => \N__49534\
        );

    \I__11640\ : LocalMux
    port map (
            O => \N__49549\,
            I => \N__49531\
        );

    \I__11639\ : Span4Mux_v
    port map (
            O => \N__49546\,
            I => \N__49524\
        );

    \I__11638\ : Span4Mux_h
    port map (
            O => \N__49541\,
            I => \N__49524\
        );

    \I__11637\ : LocalMux
    port map (
            O => \N__49538\,
            I => \N__49524\
        );

    \I__11636\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49521\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__49534\,
            I => \N__49518\
        );

    \I__11634\ : Span4Mux_h
    port map (
            O => \N__49531\,
            I => \N__49515\
        );

    \I__11633\ : Span4Mux_h
    port map (
            O => \N__49524\,
            I => \N__49512\
        );

    \I__11632\ : LocalMux
    port map (
            O => \N__49521\,
            I => \N__49505\
        );

    \I__11631\ : Span4Mux_h
    port map (
            O => \N__49518\,
            I => \N__49505\
        );

    \I__11630\ : Span4Mux_h
    port map (
            O => \N__49515\,
            I => \N__49505\
        );

    \I__11629\ : Odrv4
    port map (
            O => \N__49512\,
            I => comm_buf_0_6
        );

    \I__11628\ : Odrv4
    port map (
            O => \N__49505\,
            I => comm_buf_0_6
        );

    \I__11627\ : CascadeMux
    port map (
            O => \N__49500\,
            I => \n22545_cascade_\
        );

    \I__11626\ : CascadeMux
    port map (
            O => \N__49497\,
            I => \N__49491\
        );

    \I__11625\ : InMux
    port map (
            O => \N__49496\,
            I => \N__49488\
        );

    \I__11624\ : CascadeMux
    port map (
            O => \N__49495\,
            I => \N__49483\
        );

    \I__11623\ : InMux
    port map (
            O => \N__49494\,
            I => \N__49480\
        );

    \I__11622\ : InMux
    port map (
            O => \N__49491\,
            I => \N__49477\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__49488\,
            I => \N__49474\
        );

    \I__11620\ : CascadeMux
    port map (
            O => \N__49487\,
            I => \N__49471\
        );

    \I__11619\ : InMux
    port map (
            O => \N__49486\,
            I => \N__49468\
        );

    \I__11618\ : InMux
    port map (
            O => \N__49483\,
            I => \N__49465\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__49480\,
            I => \N__49462\
        );

    \I__11616\ : LocalMux
    port map (
            O => \N__49477\,
            I => \N__49459\
        );

    \I__11615\ : Span4Mux_v
    port map (
            O => \N__49474\,
            I => \N__49456\
        );

    \I__11614\ : InMux
    port map (
            O => \N__49471\,
            I => \N__49453\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__49468\,
            I => \N__49450\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__49465\,
            I => \N__49445\
        );

    \I__11611\ : Span4Mux_h
    port map (
            O => \N__49462\,
            I => \N__49445\
        );

    \I__11610\ : Span4Mux_h
    port map (
            O => \N__49459\,
            I => \N__49440\
        );

    \I__11609\ : Span4Mux_h
    port map (
            O => \N__49456\,
            I => \N__49440\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__49453\,
            I => \N__49433\
        );

    \I__11607\ : Span4Mux_h
    port map (
            O => \N__49450\,
            I => \N__49433\
        );

    \I__11606\ : Span4Mux_h
    port map (
            O => \N__49445\,
            I => \N__49433\
        );

    \I__11605\ : Odrv4
    port map (
            O => \N__49440\,
            I => comm_buf_1_6
        );

    \I__11604\ : Odrv4
    port map (
            O => \N__49433\,
            I => comm_buf_1_6
        );

    \I__11603\ : CEMux
    port map (
            O => \N__49428\,
            I => \N__49425\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__49425\,
            I => \N__49421\
        );

    \I__11601\ : InMux
    port map (
            O => \N__49424\,
            I => \N__49418\
        );

    \I__11600\ : Odrv4
    port map (
            O => \N__49421\,
            I => n12353
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__49418\,
            I => n12353
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49413\,
            I => \N__49410\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__49410\,
            I => \N__49407\
        );

    \I__11596\ : Span4Mux_h
    port map (
            O => \N__49407\,
            I => \N__49404\
        );

    \I__11595\ : Odrv4
    port map (
            O => \N__49404\,
            I => n14979
        );

    \I__11594\ : InMux
    port map (
            O => \N__49401\,
            I => \N__49398\
        );

    \I__11593\ : LocalMux
    port map (
            O => \N__49398\,
            I => \N__49395\
        );

    \I__11592\ : Odrv12
    port map (
            O => \N__49395\,
            I => n21588
        );

    \I__11591\ : CascadeMux
    port map (
            O => \N__49392\,
            I => \N__49379\
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__49391\,
            I => \N__49371\
        );

    \I__11589\ : CascadeMux
    port map (
            O => \N__49390\,
            I => \N__49366\
        );

    \I__11588\ : CascadeMux
    port map (
            O => \N__49389\,
            I => \N__49362\
        );

    \I__11587\ : InMux
    port map (
            O => \N__49388\,
            I => \N__49356\
        );

    \I__11586\ : InMux
    port map (
            O => \N__49387\,
            I => \N__49356\
        );

    \I__11585\ : CascadeMux
    port map (
            O => \N__49386\,
            I => \N__49352\
        );

    \I__11584\ : InMux
    port map (
            O => \N__49385\,
            I => \N__49347\
        );

    \I__11583\ : InMux
    port map (
            O => \N__49384\,
            I => \N__49342\
        );

    \I__11582\ : InMux
    port map (
            O => \N__49383\,
            I => \N__49342\
        );

    \I__11581\ : CascadeMux
    port map (
            O => \N__49382\,
            I => \N__49338\
        );

    \I__11580\ : InMux
    port map (
            O => \N__49379\,
            I => \N__49332\
        );

    \I__11579\ : InMux
    port map (
            O => \N__49378\,
            I => \N__49326\
        );

    \I__11578\ : InMux
    port map (
            O => \N__49377\,
            I => \N__49326\
        );

    \I__11577\ : CascadeMux
    port map (
            O => \N__49376\,
            I => \N__49319\
        );

    \I__11576\ : CascadeMux
    port map (
            O => \N__49375\,
            I => \N__49313\
        );

    \I__11575\ : InMux
    port map (
            O => \N__49374\,
            I => \N__49306\
        );

    \I__11574\ : InMux
    port map (
            O => \N__49371\,
            I => \N__49298\
        );

    \I__11573\ : CascadeMux
    port map (
            O => \N__49370\,
            I => \N__49294\
        );

    \I__11572\ : InMux
    port map (
            O => \N__49369\,
            I => \N__49291\
        );

    \I__11571\ : InMux
    port map (
            O => \N__49366\,
            I => \N__49284\
        );

    \I__11570\ : InMux
    port map (
            O => \N__49365\,
            I => \N__49284\
        );

    \I__11569\ : InMux
    port map (
            O => \N__49362\,
            I => \N__49284\
        );

    \I__11568\ : CascadeMux
    port map (
            O => \N__49361\,
            I => \N__49281\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__49356\,
            I => \N__49276\
        );

    \I__11566\ : CascadeMux
    port map (
            O => \N__49355\,
            I => \N__49273\
        );

    \I__11565\ : InMux
    port map (
            O => \N__49352\,
            I => \N__49269\
        );

    \I__11564\ : InMux
    port map (
            O => \N__49351\,
            I => \N__49264\
        );

    \I__11563\ : InMux
    port map (
            O => \N__49350\,
            I => \N__49264\
        );

    \I__11562\ : LocalMux
    port map (
            O => \N__49347\,
            I => \N__49259\
        );

    \I__11561\ : LocalMux
    port map (
            O => \N__49342\,
            I => \N__49259\
        );

    \I__11560\ : CascadeMux
    port map (
            O => \N__49341\,
            I => \N__49255\
        );

    \I__11559\ : InMux
    port map (
            O => \N__49338\,
            I => \N__49252\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49337\,
            I => \N__49249\
        );

    \I__11557\ : InMux
    port map (
            O => \N__49336\,
            I => \N__49244\
        );

    \I__11556\ : InMux
    port map (
            O => \N__49335\,
            I => \N__49244\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__49332\,
            I => \N__49239\
        );

    \I__11554\ : CascadeMux
    port map (
            O => \N__49331\,
            I => \N__49236\
        );

    \I__11553\ : LocalMux
    port map (
            O => \N__49326\,
            I => \N__49231\
        );

    \I__11552\ : InMux
    port map (
            O => \N__49325\,
            I => \N__49224\
        );

    \I__11551\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49224\
        );

    \I__11550\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49224\
        );

    \I__11549\ : InMux
    port map (
            O => \N__49322\,
            I => \N__49221\
        );

    \I__11548\ : InMux
    port map (
            O => \N__49319\,
            I => \N__49216\
        );

    \I__11547\ : InMux
    port map (
            O => \N__49318\,
            I => \N__49216\
        );

    \I__11546\ : CascadeMux
    port map (
            O => \N__49317\,
            I => \N__49211\
        );

    \I__11545\ : CascadeMux
    port map (
            O => \N__49316\,
            I => \N__49204\
        );

    \I__11544\ : InMux
    port map (
            O => \N__49313\,
            I => \N__49200\
        );

    \I__11543\ : InMux
    port map (
            O => \N__49312\,
            I => \N__49197\
        );

    \I__11542\ : InMux
    port map (
            O => \N__49311\,
            I => \N__49194\
        );

    \I__11541\ : InMux
    port map (
            O => \N__49310\,
            I => \N__49191\
        );

    \I__11540\ : InMux
    port map (
            O => \N__49309\,
            I => \N__49188\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__49306\,
            I => \N__49185\
        );

    \I__11538\ : InMux
    port map (
            O => \N__49305\,
            I => \N__49180\
        );

    \I__11537\ : InMux
    port map (
            O => \N__49304\,
            I => \N__49180\
        );

    \I__11536\ : InMux
    port map (
            O => \N__49303\,
            I => \N__49173\
        );

    \I__11535\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49173\
        );

    \I__11534\ : InMux
    port map (
            O => \N__49301\,
            I => \N__49173\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__49298\,
            I => \N__49170\
        );

    \I__11532\ : InMux
    port map (
            O => \N__49297\,
            I => \N__49167\
        );

    \I__11531\ : InMux
    port map (
            O => \N__49294\,
            I => \N__49164\
        );

    \I__11530\ : LocalMux
    port map (
            O => \N__49291\,
            I => \N__49159\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__49284\,
            I => \N__49159\
        );

    \I__11528\ : InMux
    port map (
            O => \N__49281\,
            I => \N__49156\
        );

    \I__11527\ : InMux
    port map (
            O => \N__49280\,
            I => \N__49151\
        );

    \I__11526\ : InMux
    port map (
            O => \N__49279\,
            I => \N__49151\
        );

    \I__11525\ : Span4Mux_h
    port map (
            O => \N__49276\,
            I => \N__49148\
        );

    \I__11524\ : InMux
    port map (
            O => \N__49273\,
            I => \N__49143\
        );

    \I__11523\ : InMux
    port map (
            O => \N__49272\,
            I => \N__49143\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__49269\,
            I => \N__49140\
        );

    \I__11521\ : LocalMux
    port map (
            O => \N__49264\,
            I => \N__49135\
        );

    \I__11520\ : Span4Mux_h
    port map (
            O => \N__49259\,
            I => \N__49135\
        );

    \I__11519\ : CascadeMux
    port map (
            O => \N__49258\,
            I => \N__49128\
        );

    \I__11518\ : InMux
    port map (
            O => \N__49255\,
            I => \N__49120\
        );

    \I__11517\ : LocalMux
    port map (
            O => \N__49252\,
            I => \N__49113\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__49249\,
            I => \N__49113\
        );

    \I__11515\ : LocalMux
    port map (
            O => \N__49244\,
            I => \N__49113\
        );

    \I__11514\ : CascadeMux
    port map (
            O => \N__49243\,
            I => \N__49109\
        );

    \I__11513\ : CascadeMux
    port map (
            O => \N__49242\,
            I => \N__49105\
        );

    \I__11512\ : Span4Mux_h
    port map (
            O => \N__49239\,
            I => \N__49100\
        );

    \I__11511\ : InMux
    port map (
            O => \N__49236\,
            I => \N__49093\
        );

    \I__11510\ : InMux
    port map (
            O => \N__49235\,
            I => \N__49093\
        );

    \I__11509\ : InMux
    port map (
            O => \N__49234\,
            I => \N__49093\
        );

    \I__11508\ : Span4Mux_v
    port map (
            O => \N__49231\,
            I => \N__49088\
        );

    \I__11507\ : LocalMux
    port map (
            O => \N__49224\,
            I => \N__49088\
        );

    \I__11506\ : LocalMux
    port map (
            O => \N__49221\,
            I => \N__49083\
        );

    \I__11505\ : LocalMux
    port map (
            O => \N__49216\,
            I => \N__49083\
        );

    \I__11504\ : InMux
    port map (
            O => \N__49215\,
            I => \N__49070\
        );

    \I__11503\ : InMux
    port map (
            O => \N__49214\,
            I => \N__49070\
        );

    \I__11502\ : InMux
    port map (
            O => \N__49211\,
            I => \N__49070\
        );

    \I__11501\ : InMux
    port map (
            O => \N__49210\,
            I => \N__49070\
        );

    \I__11500\ : InMux
    port map (
            O => \N__49209\,
            I => \N__49070\
        );

    \I__11499\ : InMux
    port map (
            O => \N__49208\,
            I => \N__49070\
        );

    \I__11498\ : InMux
    port map (
            O => \N__49207\,
            I => \N__49063\
        );

    \I__11497\ : InMux
    port map (
            O => \N__49204\,
            I => \N__49063\
        );

    \I__11496\ : InMux
    port map (
            O => \N__49203\,
            I => \N__49063\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__49200\,
            I => \N__49056\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__49197\,
            I => \N__49053\
        );

    \I__11493\ : LocalMux
    port map (
            O => \N__49194\,
            I => \N__49050\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__49191\,
            I => \N__49043\
        );

    \I__11491\ : LocalMux
    port map (
            O => \N__49188\,
            I => \N__49043\
        );

    \I__11490\ : Span4Mux_v
    port map (
            O => \N__49185\,
            I => \N__49043\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__49180\,
            I => \N__49030\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__49173\,
            I => \N__49030\
        );

    \I__11487\ : Span4Mux_v
    port map (
            O => \N__49170\,
            I => \N__49030\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__49167\,
            I => \N__49030\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__49164\,
            I => \N__49030\
        );

    \I__11484\ : Span4Mux_v
    port map (
            O => \N__49159\,
            I => \N__49030\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__49156\,
            I => \N__49021\
        );

    \I__11482\ : LocalMux
    port map (
            O => \N__49151\,
            I => \N__49021\
        );

    \I__11481\ : Span4Mux_v
    port map (
            O => \N__49148\,
            I => \N__49021\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__49143\,
            I => \N__49021\
        );

    \I__11479\ : Span4Mux_h
    port map (
            O => \N__49140\,
            I => \N__49016\
        );

    \I__11478\ : Span4Mux_h
    port map (
            O => \N__49135\,
            I => \N__49016\
        );

    \I__11477\ : InMux
    port map (
            O => \N__49134\,
            I => \N__49013\
        );

    \I__11476\ : InMux
    port map (
            O => \N__49133\,
            I => \N__49008\
        );

    \I__11475\ : InMux
    port map (
            O => \N__49132\,
            I => \N__49008\
        );

    \I__11474\ : InMux
    port map (
            O => \N__49131\,
            I => \N__48999\
        );

    \I__11473\ : InMux
    port map (
            O => \N__49128\,
            I => \N__48999\
        );

    \I__11472\ : InMux
    port map (
            O => \N__49127\,
            I => \N__48999\
        );

    \I__11471\ : InMux
    port map (
            O => \N__49126\,
            I => \N__48999\
        );

    \I__11470\ : InMux
    port map (
            O => \N__49125\,
            I => \N__48992\
        );

    \I__11469\ : InMux
    port map (
            O => \N__49124\,
            I => \N__48992\
        );

    \I__11468\ : InMux
    port map (
            O => \N__49123\,
            I => \N__48992\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__49120\,
            I => \N__48987\
        );

    \I__11466\ : Span4Mux_v
    port map (
            O => \N__49113\,
            I => \N__48987\
        );

    \I__11465\ : InMux
    port map (
            O => \N__49112\,
            I => \N__48984\
        );

    \I__11464\ : InMux
    port map (
            O => \N__49109\,
            I => \N__48973\
        );

    \I__11463\ : InMux
    port map (
            O => \N__49108\,
            I => \N__48973\
        );

    \I__11462\ : InMux
    port map (
            O => \N__49105\,
            I => \N__48973\
        );

    \I__11461\ : InMux
    port map (
            O => \N__49104\,
            I => \N__48973\
        );

    \I__11460\ : InMux
    port map (
            O => \N__49103\,
            I => \N__48973\
        );

    \I__11459\ : Span4Mux_v
    port map (
            O => \N__49100\,
            I => \N__48966\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__49093\,
            I => \N__48966\
        );

    \I__11457\ : Span4Mux_h
    port map (
            O => \N__49088\,
            I => \N__48966\
        );

    \I__11456\ : Span4Mux_v
    port map (
            O => \N__49083\,
            I => \N__48959\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__49070\,
            I => \N__48959\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__49063\,
            I => \N__48959\
        );

    \I__11453\ : InMux
    port map (
            O => \N__49062\,
            I => \N__48956\
        );

    \I__11452\ : InMux
    port map (
            O => \N__49061\,
            I => \N__48949\
        );

    \I__11451\ : InMux
    port map (
            O => \N__49060\,
            I => \N__48949\
        );

    \I__11450\ : InMux
    port map (
            O => \N__49059\,
            I => \N__48949\
        );

    \I__11449\ : Span12Mux_h
    port map (
            O => \N__49056\,
            I => \N__48946\
        );

    \I__11448\ : Span12Mux_v
    port map (
            O => \N__49053\,
            I => \N__48943\
        );

    \I__11447\ : Span4Mux_v
    port map (
            O => \N__49050\,
            I => \N__48936\
        );

    \I__11446\ : Span4Mux_v
    port map (
            O => \N__49043\,
            I => \N__48936\
        );

    \I__11445\ : Span4Mux_h
    port map (
            O => \N__49030\,
            I => \N__48936\
        );

    \I__11444\ : Span4Mux_h
    port map (
            O => \N__49021\,
            I => \N__48931\
        );

    \I__11443\ : Span4Mux_v
    port map (
            O => \N__49016\,
            I => \N__48931\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__49013\,
            I => \N__48926\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__49008\,
            I => \N__48926\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48999\,
            I => \N__48913\
        );

    \I__11439\ : LocalMux
    port map (
            O => \N__48992\,
            I => \N__48913\
        );

    \I__11438\ : Span4Mux_h
    port map (
            O => \N__48987\,
            I => \N__48913\
        );

    \I__11437\ : LocalMux
    port map (
            O => \N__48984\,
            I => \N__48913\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48973\,
            I => \N__48913\
        );

    \I__11435\ : Span4Mux_v
    port map (
            O => \N__48966\,
            I => \N__48913\
        );

    \I__11434\ : Span4Mux_h
    port map (
            O => \N__48959\,
            I => \N__48910\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__48956\,
            I => n9342
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__48949\,
            I => n9342
        );

    \I__11431\ : Odrv12
    port map (
            O => \N__48946\,
            I => n9342
        );

    \I__11430\ : Odrv12
    port map (
            O => \N__48943\,
            I => n9342
        );

    \I__11429\ : Odrv4
    port map (
            O => \N__48936\,
            I => n9342
        );

    \I__11428\ : Odrv4
    port map (
            O => \N__48931\,
            I => n9342
        );

    \I__11427\ : Odrv4
    port map (
            O => \N__48926\,
            I => n9342
        );

    \I__11426\ : Odrv4
    port map (
            O => \N__48913\,
            I => n9342
        );

    \I__11425\ : Odrv4
    port map (
            O => \N__48910\,
            I => n9342
        );

    \I__11424\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48888\
        );

    \I__11423\ : LocalMux
    port map (
            O => \N__48888\,
            I => \N__48885\
        );

    \I__11422\ : Span4Mux_h
    port map (
            O => \N__48885\,
            I => \N__48882\
        );

    \I__11421\ : Odrv4
    port map (
            O => \N__48882\,
            I => n18070
        );

    \I__11420\ : CEMux
    port map (
            O => \N__48879\,
            I => \N__48876\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48876\,
            I => \N__48873\
        );

    \I__11418\ : Odrv12
    port map (
            O => \N__48873\,
            I => n21033
        );

    \I__11417\ : InMux
    port map (
            O => \N__48870\,
            I => \N__48867\
        );

    \I__11416\ : LocalMux
    port map (
            O => \N__48867\,
            I => \N__48864\
        );

    \I__11415\ : Span12Mux_v
    port map (
            O => \N__48864\,
            I => \N__48861\
        );

    \I__11414\ : Odrv12
    port map (
            O => \N__48861\,
            I => n7_adj_1650
        );

    \I__11413\ : InMux
    port map (
            O => \N__48858\,
            I => \N__48855\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48855\,
            I => \N__48852\
        );

    \I__11411\ : Span4Mux_h
    port map (
            O => \N__48852\,
            I => \N__48848\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48851\,
            I => \N__48844\
        );

    \I__11409\ : Span4Mux_h
    port map (
            O => \N__48848\,
            I => \N__48841\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48847\,
            I => \N__48838\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__48844\,
            I => comm_cmd_6
        );

    \I__11406\ : Odrv4
    port map (
            O => \N__48841\,
            I => comm_cmd_6
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48838\,
            I => comm_cmd_6
        );

    \I__11404\ : InMux
    port map (
            O => \N__48831\,
            I => \N__48828\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__48828\,
            I => \N__48825\
        );

    \I__11402\ : Span4Mux_h
    port map (
            O => \N__48825\,
            I => \N__48822\
        );

    \I__11401\ : Span4Mux_h
    port map (
            O => \N__48822\,
            I => \N__48817\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48821\,
            I => \N__48812\
        );

    \I__11399\ : InMux
    port map (
            O => \N__48820\,
            I => \N__48812\
        );

    \I__11398\ : Odrv4
    port map (
            O => \N__48817\,
            I => comm_cmd_5
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48812\,
            I => comm_cmd_5
        );

    \I__11396\ : InMux
    port map (
            O => \N__48807\,
            I => \N__48804\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48804\,
            I => \N__48801\
        );

    \I__11394\ : Span4Mux_h
    port map (
            O => \N__48801\,
            I => \N__48798\
        );

    \I__11393\ : Span4Mux_h
    port map (
            O => \N__48798\,
            I => \N__48795\
        );

    \I__11392\ : Odrv4
    port map (
            O => \N__48795\,
            I => n4_adj_1455
        );

    \I__11391\ : InMux
    port map (
            O => \N__48792\,
            I => \N__48788\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48791\,
            I => \N__48785\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48788\,
            I => \N__48782\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__48785\,
            I => \N__48779\
        );

    \I__11387\ : Span4Mux_h
    port map (
            O => \N__48782\,
            I => \N__48776\
        );

    \I__11386\ : Span4Mux_h
    port map (
            O => \N__48779\,
            I => \N__48773\
        );

    \I__11385\ : Odrv4
    port map (
            O => \N__48776\,
            I => n21147
        );

    \I__11384\ : Odrv4
    port map (
            O => \N__48773\,
            I => n21147
        );

    \I__11383\ : CascadeMux
    port map (
            O => \N__48768\,
            I => \n21219_cascade_\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48765\,
            I => \N__48758\
        );

    \I__11381\ : InMux
    port map (
            O => \N__48764\,
            I => \N__48758\
        );

    \I__11380\ : InMux
    port map (
            O => \N__48763\,
            I => \N__48755\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__48758\,
            I => n21089
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__48755\,
            I => n21089
        );

    \I__11377\ : InMux
    port map (
            O => \N__48750\,
            I => \N__48746\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48749\,
            I => \N__48743\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__48746\,
            I => \N__48738\
        );

    \I__11374\ : LocalMux
    port map (
            O => \N__48743\,
            I => \N__48735\
        );

    \I__11373\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48732\
        );

    \I__11372\ : InMux
    port map (
            O => \N__48741\,
            I => \N__48729\
        );

    \I__11371\ : Odrv4
    port map (
            O => \N__48738\,
            I => n21043
        );

    \I__11370\ : Odrv4
    port map (
            O => \N__48735\,
            I => n21043
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__48732\,
            I => n21043
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__48729\,
            I => n21043
        );

    \I__11367\ : InMux
    port map (
            O => \N__48720\,
            I => \N__48717\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__48717\,
            I => \N__48714\
        );

    \I__11365\ : Span4Mux_h
    port map (
            O => \N__48714\,
            I => \N__48711\
        );

    \I__11364\ : Odrv4
    port map (
            O => \N__48711\,
            I => buf_data_vac_16
        );

    \I__11363\ : InMux
    port map (
            O => \N__48708\,
            I => \N__48704\
        );

    \I__11362\ : InMux
    port map (
            O => \N__48707\,
            I => \N__48700\
        );

    \I__11361\ : LocalMux
    port map (
            O => \N__48704\,
            I => \N__48693\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48703\,
            I => \N__48690\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__48700\,
            I => \N__48687\
        );

    \I__11358\ : InMux
    port map (
            O => \N__48699\,
            I => \N__48684\
        );

    \I__11357\ : InMux
    port map (
            O => \N__48698\,
            I => \N__48681\
        );

    \I__11356\ : InMux
    port map (
            O => \N__48697\,
            I => \N__48678\
        );

    \I__11355\ : InMux
    port map (
            O => \N__48696\,
            I => \N__48673\
        );

    \I__11354\ : Span4Mux_h
    port map (
            O => \N__48693\,
            I => \N__48668\
        );

    \I__11353\ : LocalMux
    port map (
            O => \N__48690\,
            I => \N__48668\
        );

    \I__11352\ : Span4Mux_h
    port map (
            O => \N__48687\,
            I => \N__48659\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__48684\,
            I => \N__48659\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__48681\,
            I => \N__48659\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48659\
        );

    \I__11348\ : InMux
    port map (
            O => \N__48677\,
            I => \N__48656\
        );

    \I__11347\ : InMux
    port map (
            O => \N__48676\,
            I => \N__48653\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__48673\,
            I => \N__48650\
        );

    \I__11345\ : Span4Mux_v
    port map (
            O => \N__48668\,
            I => \N__48645\
        );

    \I__11344\ : Span4Mux_v
    port map (
            O => \N__48659\,
            I => \N__48645\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__48656\,
            I => \N__48640\
        );

    \I__11342\ : LocalMux
    port map (
            O => \N__48653\,
            I => \N__48640\
        );

    \I__11341\ : Span4Mux_h
    port map (
            O => \N__48650\,
            I => \N__48635\
        );

    \I__11340\ : Span4Mux_h
    port map (
            O => \N__48645\,
            I => \N__48635\
        );

    \I__11339\ : Span12Mux_v
    port map (
            O => \N__48640\,
            I => \N__48632\
        );

    \I__11338\ : Span4Mux_v
    port map (
            O => \N__48635\,
            I => \N__48629\
        );

    \I__11337\ : Odrv12
    port map (
            O => \N__48632\,
            I => comm_rx_buf_0
        );

    \I__11336\ : Odrv4
    port map (
            O => \N__48629\,
            I => comm_rx_buf_0
        );

    \I__11335\ : CascadeMux
    port map (
            O => \N__48624\,
            I => \N__48621\
        );

    \I__11334\ : InMux
    port map (
            O => \N__48621\,
            I => \N__48618\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__48618\,
            I => comm_buf_3_0
        );

    \I__11332\ : InMux
    port map (
            O => \N__48615\,
            I => \N__48612\
        );

    \I__11331\ : LocalMux
    port map (
            O => \N__48612\,
            I => \N__48609\
        );

    \I__11330\ : Sp12to4
    port map (
            O => \N__48609\,
            I => \N__48606\
        );

    \I__11329\ : Span12Mux_v
    port map (
            O => \N__48606\,
            I => \N__48603\
        );

    \I__11328\ : Odrv12
    port map (
            O => \N__48603\,
            I => buf_data_vac_23
        );

    \I__11327\ : InMux
    port map (
            O => \N__48600\,
            I => \N__48592\
        );

    \I__11326\ : InMux
    port map (
            O => \N__48599\,
            I => \N__48589\
        );

    \I__11325\ : CascadeMux
    port map (
            O => \N__48598\,
            I => \N__48585\
        );

    \I__11324\ : CascadeMux
    port map (
            O => \N__48597\,
            I => \N__48582\
        );

    \I__11323\ : CascadeMux
    port map (
            O => \N__48596\,
            I => \N__48579\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48595\,
            I => \N__48576\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__48592\,
            I => \N__48573\
        );

    \I__11320\ : LocalMux
    port map (
            O => \N__48589\,
            I => \N__48569\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48588\,
            I => \N__48566\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48585\,
            I => \N__48563\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48560\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48579\,
            I => \N__48557\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__48576\,
            I => \N__48554\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__48573\,
            I => \N__48551\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48572\,
            I => \N__48548\
        );

    \I__11312\ : Span4Mux_v
    port map (
            O => \N__48569\,
            I => \N__48543\
        );

    \I__11311\ : LocalMux
    port map (
            O => \N__48566\,
            I => \N__48543\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__48563\,
            I => \N__48540\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__48560\,
            I => \N__48535\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__48557\,
            I => \N__48535\
        );

    \I__11307\ : Span4Mux_h
    port map (
            O => \N__48554\,
            I => \N__48528\
        );

    \I__11306\ : Span4Mux_h
    port map (
            O => \N__48551\,
            I => \N__48528\
        );

    \I__11305\ : LocalMux
    port map (
            O => \N__48548\,
            I => \N__48528\
        );

    \I__11304\ : Span4Mux_v
    port map (
            O => \N__48543\,
            I => \N__48525\
        );

    \I__11303\ : Span4Mux_v
    port map (
            O => \N__48540\,
            I => \N__48520\
        );

    \I__11302\ : Span4Mux_v
    port map (
            O => \N__48535\,
            I => \N__48520\
        );

    \I__11301\ : Span4Mux_v
    port map (
            O => \N__48528\,
            I => \N__48517\
        );

    \I__11300\ : Odrv4
    port map (
            O => \N__48525\,
            I => comm_rx_buf_7
        );

    \I__11299\ : Odrv4
    port map (
            O => \N__48520\,
            I => comm_rx_buf_7
        );

    \I__11298\ : Odrv4
    port map (
            O => \N__48517\,
            I => comm_rx_buf_7
        );

    \I__11297\ : CascadeMux
    port map (
            O => \N__48510\,
            I => \N__48507\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48507\,
            I => \N__48504\
        );

    \I__11295\ : LocalMux
    port map (
            O => \N__48504\,
            I => \N__48501\
        );

    \I__11294\ : Span4Mux_h
    port map (
            O => \N__48501\,
            I => \N__48498\
        );

    \I__11293\ : Span4Mux_h
    port map (
            O => \N__48498\,
            I => \N__48495\
        );

    \I__11292\ : Odrv4
    port map (
            O => \N__48495\,
            I => comm_buf_3_7
        );

    \I__11291\ : InMux
    port map (
            O => \N__48492\,
            I => \N__48489\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__48489\,
            I => \N__48486\
        );

    \I__11289\ : Sp12to4
    port map (
            O => \N__48486\,
            I => \N__48483\
        );

    \I__11288\ : Span12Mux_v
    port map (
            O => \N__48483\,
            I => \N__48480\
        );

    \I__11287\ : Odrv12
    port map (
            O => \N__48480\,
            I => buf_data_vac_22
        );

    \I__11286\ : InMux
    port map (
            O => \N__48477\,
            I => \N__48474\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__48474\,
            I => \N__48471\
        );

    \I__11284\ : Span4Mux_v
    port map (
            O => \N__48471\,
            I => \N__48468\
        );

    \I__11283\ : Span4Mux_v
    port map (
            O => \N__48468\,
            I => \N__48465\
        );

    \I__11282\ : Odrv4
    port map (
            O => \N__48465\,
            I => buf_data_vac_21
        );

    \I__11281\ : InMux
    port map (
            O => \N__48462\,
            I => \N__48459\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__48459\,
            I => n4
        );

    \I__11279\ : CascadeMux
    port map (
            O => \N__48456\,
            I => \n21013_cascade_\
        );

    \I__11278\ : CEMux
    port map (
            O => \N__48453\,
            I => \N__48450\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__48450\,
            I => \N__48447\
        );

    \I__11276\ : Odrv4
    port map (
            O => \N__48447\,
            I => n21035
        );

    \I__11275\ : CascadeMux
    port map (
            O => \N__48444\,
            I => \N__48441\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48441\,
            I => \N__48438\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__48438\,
            I => \N__48435\
        );

    \I__11272\ : Span4Mux_v
    port map (
            O => \N__48435\,
            I => \N__48432\
        );

    \I__11271\ : Odrv4
    port map (
            O => \N__48432\,
            I => comm_length_0
        );

    \I__11270\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48426\
        );

    \I__11269\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48423\
        );

    \I__11268\ : Span4Mux_v
    port map (
            O => \N__48423\,
            I => \N__48420\
        );

    \I__11267\ : Odrv4
    port map (
            O => \N__48420\,
            I => n4_adj_1623
        );

    \I__11266\ : InMux
    port map (
            O => \N__48417\,
            I => \N__48414\
        );

    \I__11265\ : LocalMux
    port map (
            O => \N__48414\,
            I => n3
        );

    \I__11264\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48404\
        );

    \I__11263\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48401\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48398\
        );

    \I__11261\ : CascadeMux
    port map (
            O => \N__48408\,
            I => \N__48395\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48407\,
            I => \N__48392\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__48404\,
            I => \N__48389\
        );

    \I__11258\ : LocalMux
    port map (
            O => \N__48401\,
            I => \N__48384\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__48398\,
            I => \N__48384\
        );

    \I__11256\ : InMux
    port map (
            O => \N__48395\,
            I => \N__48381\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__48392\,
            I => \N__48378\
        );

    \I__11254\ : Span4Mux_v
    port map (
            O => \N__48389\,
            I => \N__48375\
        );

    \I__11253\ : Span4Mux_v
    port map (
            O => \N__48384\,
            I => \N__48370\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__48381\,
            I => \N__48370\
        );

    \I__11251\ : Odrv12
    port map (
            O => \N__48378\,
            I => n21110
        );

    \I__11250\ : Odrv4
    port map (
            O => \N__48375\,
            I => n21110
        );

    \I__11249\ : Odrv4
    port map (
            O => \N__48370\,
            I => n21110
        );

    \I__11248\ : CascadeMux
    port map (
            O => \N__48363\,
            I => \n3_cascade_\
        );

    \I__11247\ : InMux
    port map (
            O => \N__48360\,
            I => \N__48355\
        );

    \I__11246\ : InMux
    port map (
            O => \N__48359\,
            I => \N__48350\
        );

    \I__11245\ : InMux
    port map (
            O => \N__48358\,
            I => \N__48350\
        );

    \I__11244\ : LocalMux
    port map (
            O => \N__48355\,
            I => \N__48345\
        );

    \I__11243\ : LocalMux
    port map (
            O => \N__48350\,
            I => \N__48345\
        );

    \I__11242\ : Span4Mux_h
    port map (
            O => \N__48345\,
            I => \N__48342\
        );

    \I__11241\ : Span4Mux_h
    port map (
            O => \N__48342\,
            I => \N__48338\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48341\,
            I => \N__48335\
        );

    \I__11239\ : Odrv4
    port map (
            O => \N__48338\,
            I => n12442
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__48335\,
            I => n12442
        );

    \I__11237\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48327\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48327\,
            I => n4_adj_1589
        );

    \I__11235\ : CascadeMux
    port map (
            O => \N__48324\,
            I => \n20095_cascade_\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48321\,
            I => \N__48318\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__48318\,
            I => n21013
        );

    \I__11232\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48312\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48312\,
            I => n11619
        );

    \I__11230\ : CascadeMux
    port map (
            O => \N__48309\,
            I => \N__48306\
        );

    \I__11229\ : InMux
    port map (
            O => \N__48306\,
            I => \N__48303\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__48303\,
            I => \N__48300\
        );

    \I__11227\ : Odrv4
    port map (
            O => \N__48300\,
            I => buf_data_vac_1
        );

    \I__11226\ : CEMux
    port map (
            O => \N__48297\,
            I => \N__48294\
        );

    \I__11225\ : LocalMux
    port map (
            O => \N__48294\,
            I => \N__48290\
        );

    \I__11224\ : InMux
    port map (
            O => \N__48293\,
            I => \N__48287\
        );

    \I__11223\ : Span4Mux_h
    port map (
            O => \N__48290\,
            I => \N__48284\
        );

    \I__11222\ : LocalMux
    port map (
            O => \N__48287\,
            I => \N__48281\
        );

    \I__11221\ : Odrv4
    port map (
            O => \N__48284\,
            I => n12431
        );

    \I__11220\ : Odrv4
    port map (
            O => \N__48281\,
            I => n12431
        );

    \I__11219\ : SRMux
    port map (
            O => \N__48276\,
            I => \N__48273\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__48273\,
            I => \N__48270\
        );

    \I__11217\ : Odrv4
    port map (
            O => \N__48270\,
            I => n14993
        );

    \I__11216\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48263\
        );

    \I__11215\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48260\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__48263\,
            I => \N__48254\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__48260\,
            I => \N__48251\
        );

    \I__11212\ : InMux
    port map (
            O => \N__48259\,
            I => \N__48248\
        );

    \I__11211\ : InMux
    port map (
            O => \N__48258\,
            I => \N__48245\
        );

    \I__11210\ : InMux
    port map (
            O => \N__48257\,
            I => \N__48242\
        );

    \I__11209\ : Span4Mux_h
    port map (
            O => \N__48254\,
            I => \N__48238\
        );

    \I__11208\ : Span4Mux_h
    port map (
            O => \N__48251\,
            I => \N__48232\
        );

    \I__11207\ : LocalMux
    port map (
            O => \N__48248\,
            I => \N__48232\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__48245\,
            I => \N__48229\
        );

    \I__11205\ : LocalMux
    port map (
            O => \N__48242\,
            I => \N__48226\
        );

    \I__11204\ : InMux
    port map (
            O => \N__48241\,
            I => \N__48223\
        );

    \I__11203\ : Span4Mux_h
    port map (
            O => \N__48238\,
            I => \N__48220\
        );

    \I__11202\ : InMux
    port map (
            O => \N__48237\,
            I => \N__48217\
        );

    \I__11201\ : Span4Mux_v
    port map (
            O => \N__48232\,
            I => \N__48208\
        );

    \I__11200\ : Span4Mux_v
    port map (
            O => \N__48229\,
            I => \N__48208\
        );

    \I__11199\ : Span4Mux_h
    port map (
            O => \N__48226\,
            I => \N__48208\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__48223\,
            I => \N__48208\
        );

    \I__11197\ : Odrv4
    port map (
            O => \N__48220\,
            I => n11652
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__48217\,
            I => n11652
        );

    \I__11195\ : Odrv4
    port map (
            O => \N__48208\,
            I => n11652
        );

    \I__11194\ : CascadeMux
    port map (
            O => \N__48201\,
            I => \n2_adj_1576_cascade_\
        );

    \I__11193\ : InMux
    port map (
            O => \N__48198\,
            I => \N__48195\
        );

    \I__11192\ : LocalMux
    port map (
            O => \N__48195\,
            I => n22611
        );

    \I__11191\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48189\
        );

    \I__11190\ : LocalMux
    port map (
            O => \N__48189\,
            I => \N__48185\
        );

    \I__11189\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48182\
        );

    \I__11188\ : Span4Mux_v
    port map (
            O => \N__48185\,
            I => \N__48177\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__48182\,
            I => \N__48177\
        );

    \I__11186\ : Span4Mux_h
    port map (
            O => \N__48177\,
            I => \N__48174\
        );

    \I__11185\ : Span4Mux_h
    port map (
            O => \N__48174\,
            I => \N__48171\
        );

    \I__11184\ : Odrv4
    port map (
            O => \N__48171\,
            I => \comm_state_3_N_460_3\
        );

    \I__11183\ : CascadeMux
    port map (
            O => \N__48168\,
            I => \n1348_cascade_\
        );

    \I__11182\ : CascadeMux
    port map (
            O => \N__48165\,
            I => \n21139_cascade_\
        );

    \I__11181\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48156\
        );

    \I__11180\ : InMux
    port map (
            O => \N__48161\,
            I => \N__48156\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__48156\,
            I => n1348
        );

    \I__11178\ : InMux
    port map (
            O => \N__48153\,
            I => \N__48150\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__48150\,
            I => n8_adj_1577
        );

    \I__11176\ : InMux
    port map (
            O => \N__48147\,
            I => \N__48144\
        );

    \I__11175\ : LocalMux
    port map (
            O => \N__48144\,
            I => n22614
        );

    \I__11174\ : InMux
    port map (
            O => \N__48141\,
            I => \N__48134\
        );

    \I__11173\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48131\
        );

    \I__11172\ : InMux
    port map (
            O => \N__48139\,
            I => \N__48128\
        );

    \I__11171\ : InMux
    port map (
            O => \N__48138\,
            I => \N__48125\
        );

    \I__11170\ : InMux
    port map (
            O => \N__48137\,
            I => \N__48122\
        );

    \I__11169\ : LocalMux
    port map (
            O => \N__48134\,
            I => \N__48117\
        );

    \I__11168\ : LocalMux
    port map (
            O => \N__48131\,
            I => \N__48117\
        );

    \I__11167\ : LocalMux
    port map (
            O => \N__48128\,
            I => \N__48110\
        );

    \I__11166\ : LocalMux
    port map (
            O => \N__48125\,
            I => \N__48110\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__48122\,
            I => \N__48110\
        );

    \I__11164\ : Span4Mux_v
    port map (
            O => \N__48117\,
            I => \N__48107\
        );

    \I__11163\ : Span4Mux_v
    port map (
            O => \N__48110\,
            I => \N__48104\
        );

    \I__11162\ : Sp12to4
    port map (
            O => \N__48107\,
            I => \N__48099\
        );

    \I__11161\ : Sp12to4
    port map (
            O => \N__48104\,
            I => \N__48099\
        );

    \I__11160\ : Span12Mux_h
    port map (
            O => \N__48099\,
            I => \N__48096\
        );

    \I__11159\ : Span12Mux_v
    port map (
            O => \N__48096\,
            I => \N__48093\
        );

    \I__11158\ : Odrv12
    port map (
            O => \N__48093\,
            I => \ICE_SPI_SCLK\
        );

    \I__11157\ : SRMux
    port map (
            O => \N__48090\,
            I => \N__48087\
        );

    \I__11156\ : LocalMux
    port map (
            O => \N__48087\,
            I => \N__48084\
        );

    \I__11155\ : Span4Mux_v
    port map (
            O => \N__48084\,
            I => \N__48081\
        );

    \I__11154\ : Odrv4
    port map (
            O => \N__48081\,
            I => \comm_spi.iclk_N_803\
        );

    \I__11153\ : InMux
    port map (
            O => \N__48078\,
            I => \N__48075\
        );

    \I__11152\ : LocalMux
    port map (
            O => \N__48075\,
            I => \N__48072\
        );

    \I__11151\ : Span4Mux_h
    port map (
            O => \N__48072\,
            I => \N__48069\
        );

    \I__11150\ : Odrv4
    port map (
            O => \N__48069\,
            I => buf_data_vac_0
        );

    \I__11149\ : InMux
    port map (
            O => \N__48066\,
            I => \N__48063\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__48063\,
            I => \N__48060\
        );

    \I__11147\ : Span4Mux_v
    port map (
            O => \N__48060\,
            I => \N__48057\
        );

    \I__11146\ : Span4Mux_h
    port map (
            O => \N__48057\,
            I => \N__48054\
        );

    \I__11145\ : Sp12to4
    port map (
            O => \N__48054\,
            I => \N__48051\
        );

    \I__11144\ : Odrv12
    port map (
            O => \N__48051\,
            I => buf_data_vac_7
        );

    \I__11143\ : InMux
    port map (
            O => \N__48048\,
            I => \N__48045\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__48045\,
            I => \N__48042\
        );

    \I__11141\ : Span4Mux_h
    port map (
            O => \N__48042\,
            I => \N__48039\
        );

    \I__11140\ : Odrv4
    port map (
            O => \N__48039\,
            I => comm_buf_5_7
        );

    \I__11139\ : InMux
    port map (
            O => \N__48036\,
            I => \N__48033\
        );

    \I__11138\ : LocalMux
    port map (
            O => \N__48033\,
            I => \N__48030\
        );

    \I__11137\ : Span12Mux_v
    port map (
            O => \N__48030\,
            I => \N__48027\
        );

    \I__11136\ : Span12Mux_h
    port map (
            O => \N__48027\,
            I => \N__48024\
        );

    \I__11135\ : Odrv12
    port map (
            O => \N__48024\,
            I => buf_data_vac_6
        );

    \I__11134\ : InMux
    port map (
            O => \N__48021\,
            I => \N__48018\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__48018\,
            I => \N__48015\
        );

    \I__11132\ : Span4Mux_h
    port map (
            O => \N__48015\,
            I => \N__48012\
        );

    \I__11131\ : Span4Mux_h
    port map (
            O => \N__48012\,
            I => \N__48009\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__48009\,
            I => \N__48006\
        );

    \I__11129\ : Odrv4
    port map (
            O => \N__48006\,
            I => buf_data_vac_5
        );

    \I__11128\ : InMux
    port map (
            O => \N__48003\,
            I => \N__48000\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__48000\,
            I => \N__47997\
        );

    \I__11126\ : Span4Mux_v
    port map (
            O => \N__47997\,
            I => \N__47994\
        );

    \I__11125\ : Span4Mux_h
    port map (
            O => \N__47994\,
            I => \N__47991\
        );

    \I__11124\ : Sp12to4
    port map (
            O => \N__47991\,
            I => \N__47988\
        );

    \I__11123\ : Odrv12
    port map (
            O => \N__47988\,
            I => buf_data_vac_4
        );

    \I__11122\ : InMux
    port map (
            O => \N__47985\,
            I => \N__47982\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__47982\,
            I => \N__47979\
        );

    \I__11120\ : Span4Mux_h
    port map (
            O => \N__47979\,
            I => \N__47976\
        );

    \I__11119\ : Odrv4
    port map (
            O => \N__47976\,
            I => comm_buf_5_4
        );

    \I__11118\ : InMux
    port map (
            O => \N__47973\,
            I => \N__47970\
        );

    \I__11117\ : LocalMux
    port map (
            O => \N__47970\,
            I => \N__47967\
        );

    \I__11116\ : Span4Mux_h
    port map (
            O => \N__47967\,
            I => \N__47964\
        );

    \I__11115\ : Odrv4
    port map (
            O => \N__47964\,
            I => buf_data_vac_3
        );

    \I__11114\ : CascadeMux
    port map (
            O => \N__47961\,
            I => \N__47958\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47958\,
            I => \N__47955\
        );

    \I__11112\ : LocalMux
    port map (
            O => \N__47955\,
            I => \N__47952\
        );

    \I__11111\ : Odrv4
    port map (
            O => \N__47952\,
            I => comm_buf_5_3
        );

    \I__11110\ : InMux
    port map (
            O => \N__47949\,
            I => \N__47946\
        );

    \I__11109\ : LocalMux
    port map (
            O => \N__47946\,
            I => \N__47943\
        );

    \I__11108\ : Span4Mux_v
    port map (
            O => \N__47943\,
            I => \N__47940\
        );

    \I__11107\ : Odrv4
    port map (
            O => \N__47940\,
            I => buf_data_vac_2
        );

    \I__11106\ : InMux
    port map (
            O => \N__47937\,
            I => \N__47934\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47934\,
            I => \N__47931\
        );

    \I__11104\ : Span4Mux_v
    port map (
            O => \N__47931\,
            I => \N__47928\
        );

    \I__11103\ : Odrv4
    port map (
            O => \N__47928\,
            I => comm_buf_5_2
        );

    \I__11102\ : InMux
    port map (
            O => \N__47925\,
            I => \N__47917\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47924\,
            I => \N__47911\
        );

    \I__11100\ : InMux
    port map (
            O => \N__47923\,
            I => \N__47911\
        );

    \I__11099\ : CascadeMux
    port map (
            O => \N__47922\,
            I => \N__47902\
        );

    \I__11098\ : CascadeMux
    port map (
            O => \N__47921\,
            I => \N__47899\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47920\,
            I => \N__47896\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__47917\,
            I => \N__47893\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47916\,
            I => \N__47890\
        );

    \I__11094\ : LocalMux
    port map (
            O => \N__47911\,
            I => \N__47887\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47910\,
            I => \N__47882\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47909\,
            I => \N__47882\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47908\,
            I => \N__47873\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47907\,
            I => \N__47873\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47906\,
            I => \N__47873\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47905\,
            I => \N__47873\
        );

    \I__11087\ : InMux
    port map (
            O => \N__47902\,
            I => \N__47868\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47899\,
            I => \N__47868\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47896\,
            I => \N__47865\
        );

    \I__11084\ : Span4Mux_h
    port map (
            O => \N__47893\,
            I => \N__47859\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__47890\,
            I => \N__47856\
        );

    \I__11082\ : Span4Mux_v
    port map (
            O => \N__47887\,
            I => \N__47847\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__47882\,
            I => \N__47847\
        );

    \I__11080\ : LocalMux
    port map (
            O => \N__47873\,
            I => \N__47847\
        );

    \I__11079\ : LocalMux
    port map (
            O => \N__47868\,
            I => \N__47847\
        );

    \I__11078\ : Span12Mux_v
    port map (
            O => \N__47865\,
            I => \N__47844\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47864\,
            I => \N__47841\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47863\,
            I => \N__47836\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47862\,
            I => \N__47836\
        );

    \I__11074\ : Span4Mux_h
    port map (
            O => \N__47859\,
            I => \N__47829\
        );

    \I__11073\ : Span4Mux_v
    port map (
            O => \N__47856\,
            I => \N__47829\
        );

    \I__11072\ : Span4Mux_v
    port map (
            O => \N__47847\,
            I => \N__47829\
        );

    \I__11071\ : Odrv12
    port map (
            O => \N__47844\,
            I => n12654
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__47841\,
            I => n12654
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__47836\,
            I => n12654
        );

    \I__11068\ : Odrv4
    port map (
            O => \N__47829\,
            I => n12654
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__47820\,
            I => \N__47816\
        );

    \I__11066\ : CascadeMux
    port map (
            O => \N__47819\,
            I => \N__47812\
        );

    \I__11065\ : InMux
    port map (
            O => \N__47816\,
            I => \N__47809\
        );

    \I__11064\ : CascadeMux
    port map (
            O => \N__47815\,
            I => \N__47806\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47812\,
            I => \N__47803\
        );

    \I__11062\ : LocalMux
    port map (
            O => \N__47809\,
            I => \N__47800\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47806\,
            I => \N__47796\
        );

    \I__11060\ : LocalMux
    port map (
            O => \N__47803\,
            I => \N__47791\
        );

    \I__11059\ : Span4Mux_v
    port map (
            O => \N__47800\,
            I => \N__47791\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47799\,
            I => \N__47788\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47796\,
            I => \N__47783\
        );

    \I__11056\ : Span4Mux_v
    port map (
            O => \N__47791\,
            I => \N__47778\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47778\
        );

    \I__11054\ : InMux
    port map (
            O => \N__47787\,
            I => \N__47775\
        );

    \I__11053\ : InMux
    port map (
            O => \N__47786\,
            I => \N__47771\
        );

    \I__11052\ : Span4Mux_v
    port map (
            O => \N__47783\,
            I => \N__47768\
        );

    \I__11051\ : Span4Mux_v
    port map (
            O => \N__47778\,
            I => \N__47763\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47775\,
            I => \N__47763\
        );

    \I__11049\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47760\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47771\,
            I => \N__47756\
        );

    \I__11047\ : Span4Mux_v
    port map (
            O => \N__47768\,
            I => \N__47751\
        );

    \I__11046\ : Span4Mux_h
    port map (
            O => \N__47763\,
            I => \N__47751\
        );

    \I__11045\ : LocalMux
    port map (
            O => \N__47760\,
            I => \N__47748\
        );

    \I__11044\ : InMux
    port map (
            O => \N__47759\,
            I => \N__47745\
        );

    \I__11043\ : Span4Mux_h
    port map (
            O => \N__47756\,
            I => \N__47742\
        );

    \I__11042\ : Odrv4
    port map (
            O => \N__47751\,
            I => comm_buf_0_4
        );

    \I__11041\ : Odrv12
    port map (
            O => \N__47748\,
            I => comm_buf_0_4
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__47745\,
            I => comm_buf_0_4
        );

    \I__11039\ : Odrv4
    port map (
            O => \N__47742\,
            I => comm_buf_0_4
        );

    \I__11038\ : InMux
    port map (
            O => \N__47733\,
            I => \N__47730\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__47730\,
            I => \N__47725\
        );

    \I__11036\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47718\
        );

    \I__11035\ : CascadeMux
    port map (
            O => \N__47728\,
            I => \N__47713\
        );

    \I__11034\ : Span4Mux_h
    port map (
            O => \N__47725\,
            I => \N__47688\
        );

    \I__11033\ : InMux
    port map (
            O => \N__47724\,
            I => \N__47679\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47723\,
            I => \N__47679\
        );

    \I__11031\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47679\
        );

    \I__11030\ : InMux
    port map (
            O => \N__47721\,
            I => \N__47679\
        );

    \I__11029\ : LocalMux
    port map (
            O => \N__47718\,
            I => \N__47668\
        );

    \I__11028\ : InMux
    port map (
            O => \N__47717\,
            I => \N__47658\
        );

    \I__11027\ : InMux
    port map (
            O => \N__47716\,
            I => \N__47649\
        );

    \I__11026\ : InMux
    port map (
            O => \N__47713\,
            I => \N__47649\
        );

    \I__11025\ : InMux
    port map (
            O => \N__47712\,
            I => \N__47649\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47711\,
            I => \N__47649\
        );

    \I__11023\ : InMux
    port map (
            O => \N__47710\,
            I => \N__47644\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47709\,
            I => \N__47644\
        );

    \I__11021\ : CascadeMux
    port map (
            O => \N__47708\,
            I => \N__47639\
        );

    \I__11020\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47628\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47628\
        );

    \I__11018\ : InMux
    port map (
            O => \N__47705\,
            I => \N__47628\
        );

    \I__11017\ : InMux
    port map (
            O => \N__47704\,
            I => \N__47628\
        );

    \I__11016\ : InMux
    port map (
            O => \N__47703\,
            I => \N__47625\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47702\,
            I => \N__47622\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47613\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47613\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47699\,
            I => \N__47613\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47613\
        );

    \I__11010\ : InMux
    port map (
            O => \N__47697\,
            I => \N__47608\
        );

    \I__11009\ : InMux
    port map (
            O => \N__47696\,
            I => \N__47608\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47695\,
            I => \N__47605\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47694\,
            I => \N__47602\
        );

    \I__11006\ : InMux
    port map (
            O => \N__47693\,
            I => \N__47594\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47692\,
            I => \N__47594\
        );

    \I__11004\ : InMux
    port map (
            O => \N__47691\,
            I => \N__47594\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__47688\,
            I => \N__47589\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__47679\,
            I => \N__47589\
        );

    \I__11001\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47578\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47578\
        );

    \I__10999\ : InMux
    port map (
            O => \N__47676\,
            I => \N__47578\
        );

    \I__10998\ : InMux
    port map (
            O => \N__47675\,
            I => \N__47578\
        );

    \I__10997\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47578\
        );

    \I__10996\ : InMux
    port map (
            O => \N__47673\,
            I => \N__47571\
        );

    \I__10995\ : InMux
    port map (
            O => \N__47672\,
            I => \N__47571\
        );

    \I__10994\ : InMux
    port map (
            O => \N__47671\,
            I => \N__47571\
        );

    \I__10993\ : Span4Mux_h
    port map (
            O => \N__47668\,
            I => \N__47568\
        );

    \I__10992\ : InMux
    port map (
            O => \N__47667\,
            I => \N__47565\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47666\,
            I => \N__47560\
        );

    \I__10990\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47557\
        );

    \I__10989\ : InMux
    port map (
            O => \N__47664\,
            I => \N__47548\
        );

    \I__10988\ : InMux
    port map (
            O => \N__47663\,
            I => \N__47548\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47662\,
            I => \N__47548\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47548\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47658\,
            I => \N__47541\
        );

    \I__10984\ : LocalMux
    port map (
            O => \N__47649\,
            I => \N__47541\
        );

    \I__10983\ : LocalMux
    port map (
            O => \N__47644\,
            I => \N__47541\
        );

    \I__10982\ : InMux
    port map (
            O => \N__47643\,
            I => \N__47538\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47533\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47639\,
            I => \N__47524\
        );

    \I__10979\ : InMux
    port map (
            O => \N__47638\,
            I => \N__47524\
        );

    \I__10978\ : InMux
    port map (
            O => \N__47637\,
            I => \N__47521\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__47628\,
            I => \N__47510\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__47625\,
            I => \N__47510\
        );

    \I__10975\ : LocalMux
    port map (
            O => \N__47622\,
            I => \N__47507\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__47613\,
            I => \N__47502\
        );

    \I__10973\ : LocalMux
    port map (
            O => \N__47608\,
            I => \N__47502\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__47605\,
            I => \N__47495\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__47602\,
            I => \N__47495\
        );

    \I__10970\ : InMux
    port map (
            O => \N__47601\,
            I => \N__47492\
        );

    \I__10969\ : LocalMux
    port map (
            O => \N__47594\,
            I => \N__47485\
        );

    \I__10968\ : Span4Mux_v
    port map (
            O => \N__47589\,
            I => \N__47485\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__47578\,
            I => \N__47485\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__47571\,
            I => \N__47478\
        );

    \I__10965\ : Span4Mux_h
    port map (
            O => \N__47568\,
            I => \N__47478\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__47565\,
            I => \N__47478\
        );

    \I__10963\ : InMux
    port map (
            O => \N__47564\,
            I => \N__47473\
        );

    \I__10962\ : InMux
    port map (
            O => \N__47563\,
            I => \N__47473\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__47560\,
            I => \N__47468\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__47557\,
            I => \N__47468\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__47548\,
            I => \N__47461\
        );

    \I__10958\ : Span4Mux_v
    port map (
            O => \N__47541\,
            I => \N__47461\
        );

    \I__10957\ : LocalMux
    port map (
            O => \N__47538\,
            I => \N__47461\
        );

    \I__10956\ : CascadeMux
    port map (
            O => \N__47537\,
            I => \N__47458\
        );

    \I__10955\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47454\
        );

    \I__10954\ : LocalMux
    port map (
            O => \N__47533\,
            I => \N__47446\
        );

    \I__10953\ : InMux
    port map (
            O => \N__47532\,
            I => \N__47443\
        );

    \I__10952\ : InMux
    port map (
            O => \N__47531\,
            I => \N__47436\
        );

    \I__10951\ : InMux
    port map (
            O => \N__47530\,
            I => \N__47436\
        );

    \I__10950\ : InMux
    port map (
            O => \N__47529\,
            I => \N__47436\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__47524\,
            I => \N__47431\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__47521\,
            I => \N__47431\
        );

    \I__10947\ : InMux
    port map (
            O => \N__47520\,
            I => \N__47424\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47519\,
            I => \N__47424\
        );

    \I__10945\ : InMux
    port map (
            O => \N__47518\,
            I => \N__47424\
        );

    \I__10944\ : InMux
    port map (
            O => \N__47517\,
            I => \N__47419\
        );

    \I__10943\ : InMux
    port map (
            O => \N__47516\,
            I => \N__47419\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47515\,
            I => \N__47416\
        );

    \I__10941\ : Span4Mux_v
    port map (
            O => \N__47510\,
            I => \N__47409\
        );

    \I__10940\ : Span4Mux_v
    port map (
            O => \N__47507\,
            I => \N__47409\
        );

    \I__10939\ : Span4Mux_v
    port map (
            O => \N__47502\,
            I => \N__47409\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47404\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47500\,
            I => \N__47404\
        );

    \I__10936\ : Span4Mux_h
    port map (
            O => \N__47495\,
            I => \N__47397\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__47492\,
            I => \N__47397\
        );

    \I__10934\ : Span4Mux_h
    port map (
            O => \N__47485\,
            I => \N__47397\
        );

    \I__10933\ : Span4Mux_v
    port map (
            O => \N__47478\,
            I => \N__47394\
        );

    \I__10932\ : LocalMux
    port map (
            O => \N__47473\,
            I => \N__47387\
        );

    \I__10931\ : Span4Mux_v
    port map (
            O => \N__47468\,
            I => \N__47387\
        );

    \I__10930\ : Span4Mux_h
    port map (
            O => \N__47461\,
            I => \N__47387\
        );

    \I__10929\ : InMux
    port map (
            O => \N__47458\,
            I => \N__47384\
        );

    \I__10928\ : InMux
    port map (
            O => \N__47457\,
            I => \N__47381\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__47454\,
            I => \N__47378\
        );

    \I__10926\ : InMux
    port map (
            O => \N__47453\,
            I => \N__47375\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47452\,
            I => \N__47370\
        );

    \I__10924\ : InMux
    port map (
            O => \N__47451\,
            I => \N__47370\
        );

    \I__10923\ : InMux
    port map (
            O => \N__47450\,
            I => \N__47365\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47449\,
            I => \N__47365\
        );

    \I__10921\ : Span12Mux_h
    port map (
            O => \N__47446\,
            I => \N__47360\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__47443\,
            I => \N__47360\
        );

    \I__10919\ : LocalMux
    port map (
            O => \N__47436\,
            I => \N__47347\
        );

    \I__10918\ : Span12Mux_v
    port map (
            O => \N__47431\,
            I => \N__47347\
        );

    \I__10917\ : LocalMux
    port map (
            O => \N__47424\,
            I => \N__47347\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__47419\,
            I => \N__47347\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__47416\,
            I => \N__47347\
        );

    \I__10914\ : Sp12to4
    port map (
            O => \N__47409\,
            I => \N__47347\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47342\
        );

    \I__10912\ : Span4Mux_h
    port map (
            O => \N__47397\,
            I => \N__47342\
        );

    \I__10911\ : Span4Mux_h
    port map (
            O => \N__47394\,
            I => \N__47337\
        );

    \I__10910\ : Span4Mux_h
    port map (
            O => \N__47387\,
            I => \N__47337\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__47384\,
            I => comm_cmd_2
        );

    \I__10908\ : LocalMux
    port map (
            O => \N__47381\,
            I => comm_cmd_2
        );

    \I__10907\ : Odrv4
    port map (
            O => \N__47378\,
            I => comm_cmd_2
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__47375\,
            I => comm_cmd_2
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__47370\,
            I => comm_cmd_2
        );

    \I__10904\ : LocalMux
    port map (
            O => \N__47365\,
            I => comm_cmd_2
        );

    \I__10903\ : Odrv12
    port map (
            O => \N__47360\,
            I => comm_cmd_2
        );

    \I__10902\ : Odrv12
    port map (
            O => \N__47347\,
            I => comm_cmd_2
        );

    \I__10901\ : Odrv4
    port map (
            O => \N__47342\,
            I => comm_cmd_2
        );

    \I__10900\ : Odrv4
    port map (
            O => \N__47337\,
            I => comm_cmd_2
        );

    \I__10899\ : CascadeMux
    port map (
            O => \N__47316\,
            I => \N__47313\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47313\,
            I => \N__47310\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__47310\,
            I => n21368
        );

    \I__10896\ : InMux
    port map (
            O => \N__47307\,
            I => \N__47304\
        );

    \I__10895\ : LocalMux
    port map (
            O => \N__47304\,
            I => n21369
        );

    \I__10894\ : InMux
    port map (
            O => \N__47301\,
            I => \N__47298\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__47298\,
            I => \N__47295\
        );

    \I__10892\ : Odrv4
    port map (
            O => \N__47295\,
            I => n21362
        );

    \I__10891\ : InMux
    port map (
            O => \N__47292\,
            I => \N__47289\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__47289\,
            I => \N__47286\
        );

    \I__10889\ : Span4Mux_h
    port map (
            O => \N__47286\,
            I => \N__47283\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__47283\,
            I => \N__47280\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__47280\,
            I => \N__47277\
        );

    \I__10886\ : Odrv4
    port map (
            O => \N__47277\,
            I => n21363
        );

    \I__10885\ : CascadeMux
    port map (
            O => \N__47274\,
            I => \n22599_cascade_\
        );

    \I__10884\ : InMux
    port map (
            O => \N__47271\,
            I => \N__47264\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47270\,
            I => \N__47259\
        );

    \I__10882\ : InMux
    port map (
            O => \N__47269\,
            I => \N__47246\
        );

    \I__10881\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47240\
        );

    \I__10880\ : InMux
    port map (
            O => \N__47267\,
            I => \N__47237\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47264\,
            I => \N__47234\
        );

    \I__10878\ : InMux
    port map (
            O => \N__47263\,
            I => \N__47227\
        );

    \I__10877\ : InMux
    port map (
            O => \N__47262\,
            I => \N__47227\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__47259\,
            I => \N__47224\
        );

    \I__10875\ : InMux
    port map (
            O => \N__47258\,
            I => \N__47221\
        );

    \I__10874\ : InMux
    port map (
            O => \N__47257\,
            I => \N__47218\
        );

    \I__10873\ : InMux
    port map (
            O => \N__47256\,
            I => \N__47215\
        );

    \I__10872\ : InMux
    port map (
            O => \N__47255\,
            I => \N__47212\
        );

    \I__10871\ : InMux
    port map (
            O => \N__47254\,
            I => \N__47209\
        );

    \I__10870\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47204\
        );

    \I__10869\ : InMux
    port map (
            O => \N__47252\,
            I => \N__47204\
        );

    \I__10868\ : InMux
    port map (
            O => \N__47251\,
            I => \N__47197\
        );

    \I__10867\ : InMux
    port map (
            O => \N__47250\,
            I => \N__47197\
        );

    \I__10866\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47197\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__47246\,
            I => \N__47187\
        );

    \I__10864\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47182\
        );

    \I__10863\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47182\
        );

    \I__10862\ : InMux
    port map (
            O => \N__47243\,
            I => \N__47179\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__47240\,
            I => \N__47176\
        );

    \I__10860\ : LocalMux
    port map (
            O => \N__47237\,
            I => \N__47171\
        );

    \I__10859\ : Span4Mux_v
    port map (
            O => \N__47234\,
            I => \N__47171\
        );

    \I__10858\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47166\
        );

    \I__10857\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47166\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__47227\,
            I => \N__47160\
        );

    \I__10855\ : Span4Mux_v
    port map (
            O => \N__47224\,
            I => \N__47155\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__47221\,
            I => \N__47150\
        );

    \I__10853\ : LocalMux
    port map (
            O => \N__47218\,
            I => \N__47137\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__47215\,
            I => \N__47137\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__47212\,
            I => \N__47137\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__47209\,
            I => \N__47137\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__47204\,
            I => \N__47137\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__47197\,
            I => \N__47137\
        );

    \I__10847\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47128\
        );

    \I__10846\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47123\
        );

    \I__10845\ : InMux
    port map (
            O => \N__47194\,
            I => \N__47123\
        );

    \I__10844\ : InMux
    port map (
            O => \N__47193\,
            I => \N__47120\
        );

    \I__10843\ : InMux
    port map (
            O => \N__47192\,
            I => \N__47117\
        );

    \I__10842\ : InMux
    port map (
            O => \N__47191\,
            I => \N__47112\
        );

    \I__10841\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47112\
        );

    \I__10840\ : Span4Mux_h
    port map (
            O => \N__47187\,
            I => \N__47107\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__47182\,
            I => \N__47107\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__47179\,
            I => \N__47098\
        );

    \I__10837\ : Span4Mux_h
    port map (
            O => \N__47176\,
            I => \N__47098\
        );

    \I__10836\ : Span4Mux_v
    port map (
            O => \N__47171\,
            I => \N__47098\
        );

    \I__10835\ : LocalMux
    port map (
            O => \N__47166\,
            I => \N__47098\
        );

    \I__10834\ : InMux
    port map (
            O => \N__47165\,
            I => \N__47095\
        );

    \I__10833\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47092\
        );

    \I__10832\ : InMux
    port map (
            O => \N__47163\,
            I => \N__47088\
        );

    \I__10831\ : Sp12to4
    port map (
            O => \N__47160\,
            I => \N__47085\
        );

    \I__10830\ : InMux
    port map (
            O => \N__47159\,
            I => \N__47080\
        );

    \I__10829\ : InMux
    port map (
            O => \N__47158\,
            I => \N__47080\
        );

    \I__10828\ : Span4Mux_v
    port map (
            O => \N__47155\,
            I => \N__47077\
        );

    \I__10827\ : InMux
    port map (
            O => \N__47154\,
            I => \N__47072\
        );

    \I__10826\ : InMux
    port map (
            O => \N__47153\,
            I => \N__47072\
        );

    \I__10825\ : Span4Mux_v
    port map (
            O => \N__47150\,
            I => \N__47067\
        );

    \I__10824\ : Span4Mux_v
    port map (
            O => \N__47137\,
            I => \N__47067\
        );

    \I__10823\ : InMux
    port map (
            O => \N__47136\,
            I => \N__47058\
        );

    \I__10822\ : InMux
    port map (
            O => \N__47135\,
            I => \N__47058\
        );

    \I__10821\ : InMux
    port map (
            O => \N__47134\,
            I => \N__47058\
        );

    \I__10820\ : InMux
    port map (
            O => \N__47133\,
            I => \N__47058\
        );

    \I__10819\ : InMux
    port map (
            O => \N__47132\,
            I => \N__47055\
        );

    \I__10818\ : CascadeMux
    port map (
            O => \N__47131\,
            I => \N__47052\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__47128\,
            I => \N__47049\
        );

    \I__10816\ : LocalMux
    port map (
            O => \N__47123\,
            I => \N__47041\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__47120\,
            I => \N__47041\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__47117\,
            I => \N__47041\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47034\
        );

    \I__10812\ : Span4Mux_v
    port map (
            O => \N__47107\,
            I => \N__47034\
        );

    \I__10811\ : Span4Mux_h
    port map (
            O => \N__47098\,
            I => \N__47034\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__47095\,
            I => \N__47029\
        );

    \I__10809\ : LocalMux
    port map (
            O => \N__47092\,
            I => \N__47029\
        );

    \I__10808\ : InMux
    port map (
            O => \N__47091\,
            I => \N__47026\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__47088\,
            I => \N__47009\
        );

    \I__10806\ : Span12Mux_v
    port map (
            O => \N__47085\,
            I => \N__47009\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__47080\,
            I => \N__47009\
        );

    \I__10804\ : Sp12to4
    port map (
            O => \N__47077\,
            I => \N__47009\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__47072\,
            I => \N__47009\
        );

    \I__10802\ : Sp12to4
    port map (
            O => \N__47067\,
            I => \N__47009\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__47058\,
            I => \N__47009\
        );

    \I__10800\ : LocalMux
    port map (
            O => \N__47055\,
            I => \N__47009\
        );

    \I__10799\ : InMux
    port map (
            O => \N__47052\,
            I => \N__47006\
        );

    \I__10798\ : Span12Mux_h
    port map (
            O => \N__47049\,
            I => \N__47003\
        );

    \I__10797\ : InMux
    port map (
            O => \N__47048\,
            I => \N__47000\
        );

    \I__10796\ : Span12Mux_h
    port map (
            O => \N__47041\,
            I => \N__46997\
        );

    \I__10795\ : Span4Mux_h
    port map (
            O => \N__47034\,
            I => \N__46994\
        );

    \I__10794\ : Span4Mux_h
    port map (
            O => \N__47029\,
            I => \N__46991\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__47026\,
            I => \N__46986\
        );

    \I__10792\ : Span12Mux_h
    port map (
            O => \N__47009\,
            I => \N__46986\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__47006\,
            I => comm_cmd_3
        );

    \I__10790\ : Odrv12
    port map (
            O => \N__47003\,
            I => comm_cmd_3
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__47000\,
            I => comm_cmd_3
        );

    \I__10788\ : Odrv12
    port map (
            O => \N__46997\,
            I => comm_cmd_3
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__46994\,
            I => comm_cmd_3
        );

    \I__10786\ : Odrv4
    port map (
            O => \N__46991\,
            I => comm_cmd_3
        );

    \I__10785\ : Odrv12
    port map (
            O => \N__46986\,
            I => comm_cmd_3
        );

    \I__10784\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46968\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__46968\,
            I => n22602
        );

    \I__10782\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46962\
        );

    \I__10781\ : LocalMux
    port map (
            O => \N__46962\,
            I => \N__46959\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__46959\,
            I => \N__46954\
        );

    \I__10779\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46951\
        );

    \I__10778\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46948\
        );

    \I__10777\ : Sp12to4
    port map (
            O => \N__46954\,
            I => \N__46943\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__46951\,
            I => \N__46943\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46948\,
            I => buf_dds1_6
        );

    \I__10774\ : Odrv12
    port map (
            O => \N__46943\,
            I => buf_dds1_6
        );

    \I__10773\ : InMux
    port map (
            O => \N__46938\,
            I => \N__46935\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__46935\,
            I => \N__46931\
        );

    \I__10771\ : CascadeMux
    port map (
            O => \N__46934\,
            I => \N__46928\
        );

    \I__10770\ : Span4Mux_h
    port map (
            O => \N__46931\,
            I => \N__46925\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46922\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__46925\,
            I => n68
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__46922\,
            I => n68
        );

    \I__10766\ : CascadeMux
    port map (
            O => \N__46917\,
            I => \N__46911\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46906\
        );

    \I__10764\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46903\
        );

    \I__10763\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46900\
        );

    \I__10762\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46895\
        );

    \I__10761\ : CascadeMux
    port map (
            O => \N__46910\,
            I => \N__46891\
        );

    \I__10760\ : InMux
    port map (
            O => \N__46909\,
            I => \N__46886\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__46906\,
            I => \N__46878\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__46903\,
            I => \N__46878\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__46900\,
            I => \N__46878\
        );

    \I__10756\ : CascadeMux
    port map (
            O => \N__46899\,
            I => \N__46875\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46898\,
            I => \N__46869\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__46895\,
            I => \N__46866\
        );

    \I__10753\ : InMux
    port map (
            O => \N__46894\,
            I => \N__46859\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46859\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46890\,
            I => \N__46859\
        );

    \I__10750\ : InMux
    port map (
            O => \N__46889\,
            I => \N__46856\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__46886\,
            I => \N__46853\
        );

    \I__10748\ : InMux
    port map (
            O => \N__46885\,
            I => \N__46850\
        );

    \I__10747\ : Span4Mux_v
    port map (
            O => \N__46878\,
            I => \N__46847\
        );

    \I__10746\ : InMux
    port map (
            O => \N__46875\,
            I => \N__46842\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46842\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46873\,
            I => \N__46839\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46872\,
            I => \N__46836\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__46869\,
            I => \N__46833\
        );

    \I__10741\ : Span4Mux_h
    port map (
            O => \N__46866\,
            I => \N__46828\
        );

    \I__10740\ : LocalMux
    port map (
            O => \N__46859\,
            I => \N__46828\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46856\,
            I => \N__46823\
        );

    \I__10738\ : Span4Mux_h
    port map (
            O => \N__46853\,
            I => \N__46823\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__46850\,
            I => \N__46818\
        );

    \I__10736\ : Span4Mux_h
    port map (
            O => \N__46847\,
            I => \N__46818\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__46842\,
            I => \N__46811\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__46839\,
            I => \N__46811\
        );

    \I__10733\ : LocalMux
    port map (
            O => \N__46836\,
            I => \N__46811\
        );

    \I__10732\ : Span4Mux_h
    port map (
            O => \N__46833\,
            I => \N__46807\
        );

    \I__10731\ : Span4Mux_v
    port map (
            O => \N__46828\,
            I => \N__46804\
        );

    \I__10730\ : Span4Mux_h
    port map (
            O => \N__46823\,
            I => \N__46801\
        );

    \I__10729\ : Span4Mux_h
    port map (
            O => \N__46818\,
            I => \N__46796\
        );

    \I__10728\ : Span4Mux_v
    port map (
            O => \N__46811\,
            I => \N__46796\
        );

    \I__10727\ : InMux
    port map (
            O => \N__46810\,
            I => \N__46793\
        );

    \I__10726\ : Span4Mux_v
    port map (
            O => \N__46807\,
            I => \N__46790\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__46804\,
            I => \N__46787\
        );

    \I__10724\ : Span4Mux_h
    port map (
            O => \N__46801\,
            I => \N__46784\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__46796\,
            I => \N__46781\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__46793\,
            I => n12048
        );

    \I__10721\ : Odrv4
    port map (
            O => \N__46790\,
            I => n12048
        );

    \I__10720\ : Odrv4
    port map (
            O => \N__46787\,
            I => n12048
        );

    \I__10719\ : Odrv4
    port map (
            O => \N__46784\,
            I => n12048
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__46781\,
            I => n12048
        );

    \I__10717\ : CascadeMux
    port map (
            O => \N__46770\,
            I => \n12048_cascade_\
        );

    \I__10716\ : CascadeMux
    port map (
            O => \N__46767\,
            I => \N__46760\
        );

    \I__10715\ : InMux
    port map (
            O => \N__46766\,
            I => \N__46757\
        );

    \I__10714\ : InMux
    port map (
            O => \N__46765\,
            I => \N__46747\
        );

    \I__10713\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46747\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46763\,
            I => \N__46747\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46760\,
            I => \N__46742\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__46757\,
            I => \N__46739\
        );

    \I__10709\ : InMux
    port map (
            O => \N__46756\,
            I => \N__46734\
        );

    \I__10708\ : InMux
    port map (
            O => \N__46755\,
            I => \N__46734\
        );

    \I__10707\ : InMux
    port map (
            O => \N__46754\,
            I => \N__46729\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46747\,
            I => \N__46726\
        );

    \I__10705\ : InMux
    port map (
            O => \N__46746\,
            I => \N__46723\
        );

    \I__10704\ : InMux
    port map (
            O => \N__46745\,
            I => \N__46720\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__46742\,
            I => \N__46717\
        );

    \I__10702\ : Span4Mux_v
    port map (
            O => \N__46739\,
            I => \N__46712\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__46734\,
            I => \N__46712\
        );

    \I__10700\ : InMux
    port map (
            O => \N__46733\,
            I => \N__46709\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46732\,
            I => \N__46706\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__46729\,
            I => \N__46703\
        );

    \I__10697\ : Span4Mux_v
    port map (
            O => \N__46726\,
            I => \N__46700\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__46723\,
            I => \N__46697\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__46720\,
            I => \N__46689\
        );

    \I__10694\ : Span4Mux_v
    port map (
            O => \N__46717\,
            I => \N__46689\
        );

    \I__10693\ : Span4Mux_h
    port map (
            O => \N__46712\,
            I => \N__46689\
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__46709\,
            I => \N__46686\
        );

    \I__10691\ : LocalMux
    port map (
            O => \N__46706\,
            I => \N__46681\
        );

    \I__10690\ : Span4Mux_v
    port map (
            O => \N__46703\,
            I => \N__46681\
        );

    \I__10689\ : Span4Mux_h
    port map (
            O => \N__46700\,
            I => \N__46676\
        );

    \I__10688\ : Span4Mux_h
    port map (
            O => \N__46697\,
            I => \N__46676\
        );

    \I__10687\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46673\
        );

    \I__10686\ : Span4Mux_h
    port map (
            O => \N__46689\,
            I => \N__46670\
        );

    \I__10685\ : Span12Mux_v
    port map (
            O => \N__46686\,
            I => \N__46665\
        );

    \I__10684\ : Sp12to4
    port map (
            O => \N__46681\,
            I => \N__46665\
        );

    \I__10683\ : Span4Mux_v
    port map (
            O => \N__46676\,
            I => \N__46662\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__46673\,
            I => n16971
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__46670\,
            I => n16971
        );

    \I__10680\ : Odrv12
    port map (
            O => \N__46665\,
            I => n16971
        );

    \I__10679\ : Odrv4
    port map (
            O => \N__46662\,
            I => n16971
        );

    \I__10678\ : InMux
    port map (
            O => \N__46653\,
            I => \N__46650\
        );

    \I__10677\ : LocalMux
    port map (
            O => \N__46650\,
            I => \comm_spi.n14805\
        );

    \I__10676\ : SRMux
    port map (
            O => \N__46647\,
            I => \N__46644\
        );

    \I__10675\ : LocalMux
    port map (
            O => \N__46644\,
            I => \comm_spi.iclk_N_802\
        );

    \I__10674\ : CascadeMux
    port map (
            O => \N__46641\,
            I => \N__46637\
        );

    \I__10673\ : CascadeMux
    port map (
            O => \N__46640\,
            I => \N__46634\
        );

    \I__10672\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46631\
        );

    \I__10671\ : InMux
    port map (
            O => \N__46634\,
            I => \N__46628\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__46631\,
            I => \N__46625\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__46628\,
            I => comm_buf_6_0
        );

    \I__10668\ : Odrv4
    port map (
            O => \N__46625\,
            I => comm_buf_6_0
        );

    \I__10667\ : InMux
    port map (
            O => \N__46620\,
            I => \N__46617\
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__46617\,
            I => \N__46613\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46616\,
            I => \N__46610\
        );

    \I__10664\ : Span4Mux_v
    port map (
            O => \N__46613\,
            I => \N__46607\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__46610\,
            I => comm_buf_6_3
        );

    \I__10662\ : Odrv4
    port map (
            O => \N__46607\,
            I => comm_buf_6_3
        );

    \I__10661\ : InMux
    port map (
            O => \N__46602\,
            I => \N__46599\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46599\,
            I => \N__46595\
        );

    \I__10659\ : InMux
    port map (
            O => \N__46598\,
            I => \N__46591\
        );

    \I__10658\ : Span4Mux_h
    port map (
            O => \N__46595\,
            I => \N__46588\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46594\,
            I => \N__46585\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46591\,
            I => \acadc_skipCount_7\
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__46588\,
            I => \acadc_skipCount_7\
        );

    \I__10654\ : LocalMux
    port map (
            O => \N__46585\,
            I => \acadc_skipCount_7\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46575\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__46575\,
            I => \N__46572\
        );

    \I__10651\ : Span4Mux_v
    port map (
            O => \N__46572\,
            I => \N__46568\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46571\,
            I => \N__46564\
        );

    \I__10649\ : Span4Mux_h
    port map (
            O => \N__46568\,
            I => \N__46561\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46567\,
            I => \N__46558\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__46564\,
            I => req_data_cnt_7
        );

    \I__10646\ : Odrv4
    port map (
            O => \N__46561\,
            I => req_data_cnt_7
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__46558\,
            I => req_data_cnt_7
        );

    \I__10644\ : InMux
    port map (
            O => \N__46551\,
            I => \N__46548\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46548\,
            I => \N__46545\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__46545\,
            I => \N__46541\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46544\,
            I => \N__46538\
        );

    \I__10640\ : Span4Mux_h
    port map (
            O => \N__46541\,
            I => \N__46535\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46538\,
            I => \N__46530\
        );

    \I__10638\ : Span4Mux_v
    port map (
            O => \N__46535\,
            I => \N__46530\
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__46530\,
            I => data_idxvec_7
        );

    \I__10636\ : InMux
    port map (
            O => \N__46527\,
            I => \N__46523\
        );

    \I__10635\ : InMux
    port map (
            O => \N__46526\,
            I => \N__46520\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__46523\,
            I => \N__46516\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__46520\,
            I => \N__46513\
        );

    \I__10632\ : InMux
    port map (
            O => \N__46519\,
            I => \N__46510\
        );

    \I__10631\ : Span4Mux_v
    port map (
            O => \N__46516\,
            I => \N__46505\
        );

    \I__10630\ : Span4Mux_h
    port map (
            O => \N__46513\,
            I => \N__46505\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__46510\,
            I => data_cntvec_7
        );

    \I__10628\ : Odrv4
    port map (
            O => \N__46505\,
            I => data_cntvec_7
        );

    \I__10627\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46497\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__46497\,
            I => \N__46494\
        );

    \I__10625\ : Span4Mux_v
    port map (
            O => \N__46494\,
            I => \N__46491\
        );

    \I__10624\ : Odrv4
    port map (
            O => \N__46491\,
            I => buf_data_iac_15
        );

    \I__10623\ : CascadeMux
    port map (
            O => \N__46488\,
            I => \n26_adj_1622_cascade_\
        );

    \I__10622\ : InMux
    port map (
            O => \N__46485\,
            I => \N__46450\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46484\,
            I => \N__46445\
        );

    \I__10620\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46445\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46482\,
            I => \N__46438\
        );

    \I__10618\ : InMux
    port map (
            O => \N__46481\,
            I => \N__46438\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46480\,
            I => \N__46438\
        );

    \I__10616\ : InMux
    port map (
            O => \N__46479\,
            I => \N__46433\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46478\,
            I => \N__46433\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46477\,
            I => \N__46430\
        );

    \I__10613\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46425\
        );

    \I__10612\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46425\
        );

    \I__10611\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46418\
        );

    \I__10610\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46418\
        );

    \I__10609\ : InMux
    port map (
            O => \N__46472\,
            I => \N__46418\
        );

    \I__10608\ : InMux
    port map (
            O => \N__46471\,
            I => \N__46415\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46470\,
            I => \N__46412\
        );

    \I__10606\ : CascadeMux
    port map (
            O => \N__46469\,
            I => \N__46403\
        );

    \I__10605\ : InMux
    port map (
            O => \N__46468\,
            I => \N__46397\
        );

    \I__10604\ : InMux
    port map (
            O => \N__46467\,
            I => \N__46397\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46392\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46465\,
            I => \N__46392\
        );

    \I__10601\ : InMux
    port map (
            O => \N__46464\,
            I => \N__46387\
        );

    \I__10600\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46387\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46462\,
            I => \N__46384\
        );

    \I__10598\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46381\
        );

    \I__10597\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46378\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46360\
        );

    \I__10595\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46360\
        );

    \I__10594\ : InMux
    port map (
            O => \N__46457\,
            I => \N__46360\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46456\,
            I => \N__46360\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46455\,
            I => \N__46357\
        );

    \I__10591\ : InMux
    port map (
            O => \N__46454\,
            I => \N__46354\
        );

    \I__10590\ : InMux
    port map (
            O => \N__46453\,
            I => \N__46351\
        );

    \I__10589\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46346\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__46445\,
            I => \N__46346\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__46438\,
            I => \N__46339\
        );

    \I__10586\ : LocalMux
    port map (
            O => \N__46433\,
            I => \N__46339\
        );

    \I__10585\ : LocalMux
    port map (
            O => \N__46430\,
            I => \N__46339\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46425\,
            I => \N__46336\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__46418\,
            I => \N__46329\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__46415\,
            I => \N__46329\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__46412\,
            I => \N__46329\
        );

    \I__10580\ : InMux
    port map (
            O => \N__46411\,
            I => \N__46324\
        );

    \I__10579\ : InMux
    port map (
            O => \N__46410\,
            I => \N__46324\
        );

    \I__10578\ : InMux
    port map (
            O => \N__46409\,
            I => \N__46319\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46408\,
            I => \N__46319\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46407\,
            I => \N__46312\
        );

    \I__10575\ : InMux
    port map (
            O => \N__46406\,
            I => \N__46312\
        );

    \I__10574\ : InMux
    port map (
            O => \N__46403\,
            I => \N__46303\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46402\,
            I => \N__46292\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__46397\,
            I => \N__46287\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46392\,
            I => \N__46278\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__46387\,
            I => \N__46278\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__46384\,
            I => \N__46278\
        );

    \I__10568\ : LocalMux
    port map (
            O => \N__46381\,
            I => \N__46278\
        );

    \I__10567\ : LocalMux
    port map (
            O => \N__46378\,
            I => \N__46275\
        );

    \I__10566\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46272\
        );

    \I__10565\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46269\
        );

    \I__10564\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46262\
        );

    \I__10563\ : InMux
    port map (
            O => \N__46374\,
            I => \N__46262\
        );

    \I__10562\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46262\
        );

    \I__10561\ : InMux
    port map (
            O => \N__46372\,
            I => \N__46259\
        );

    \I__10560\ : InMux
    port map (
            O => \N__46371\,
            I => \N__46249\
        );

    \I__10559\ : InMux
    port map (
            O => \N__46370\,
            I => \N__46249\
        );

    \I__10558\ : InMux
    port map (
            O => \N__46369\,
            I => \N__46249\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__46360\,
            I => \N__46244\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__46357\,
            I => \N__46244\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__46354\,
            I => \N__46241\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46351\,
            I => \N__46238\
        );

    \I__10553\ : Span4Mux_v
    port map (
            O => \N__46346\,
            I => \N__46225\
        );

    \I__10552\ : Span4Mux_v
    port map (
            O => \N__46339\,
            I => \N__46225\
        );

    \I__10551\ : Span4Mux_v
    port map (
            O => \N__46336\,
            I => \N__46225\
        );

    \I__10550\ : Span4Mux_v
    port map (
            O => \N__46329\,
            I => \N__46225\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__46324\,
            I => \N__46225\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__46319\,
            I => \N__46225\
        );

    \I__10547\ : InMux
    port map (
            O => \N__46318\,
            I => \N__46221\
        );

    \I__10546\ : InMux
    port map (
            O => \N__46317\,
            I => \N__46218\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__46312\,
            I => \N__46215\
        );

    \I__10544\ : InMux
    port map (
            O => \N__46311\,
            I => \N__46210\
        );

    \I__10543\ : InMux
    port map (
            O => \N__46310\,
            I => \N__46210\
        );

    \I__10542\ : InMux
    port map (
            O => \N__46309\,
            I => \N__46203\
        );

    \I__10541\ : InMux
    port map (
            O => \N__46308\,
            I => \N__46203\
        );

    \I__10540\ : InMux
    port map (
            O => \N__46307\,
            I => \N__46203\
        );

    \I__10539\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46200\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__46303\,
            I => \N__46197\
        );

    \I__10537\ : InMux
    port map (
            O => \N__46302\,
            I => \N__46186\
        );

    \I__10536\ : InMux
    port map (
            O => \N__46301\,
            I => \N__46186\
        );

    \I__10535\ : InMux
    port map (
            O => \N__46300\,
            I => \N__46186\
        );

    \I__10534\ : InMux
    port map (
            O => \N__46299\,
            I => \N__46186\
        );

    \I__10533\ : InMux
    port map (
            O => \N__46298\,
            I => \N__46186\
        );

    \I__10532\ : InMux
    port map (
            O => \N__46297\,
            I => \N__46183\
        );

    \I__10531\ : InMux
    port map (
            O => \N__46296\,
            I => \N__46178\
        );

    \I__10530\ : InMux
    port map (
            O => \N__46295\,
            I => \N__46178\
        );

    \I__10529\ : LocalMux
    port map (
            O => \N__46292\,
            I => \N__46175\
        );

    \I__10528\ : InMux
    port map (
            O => \N__46291\,
            I => \N__46172\
        );

    \I__10527\ : InMux
    port map (
            O => \N__46290\,
            I => \N__46169\
        );

    \I__10526\ : Span4Mux_v
    port map (
            O => \N__46287\,
            I => \N__46160\
        );

    \I__10525\ : Span4Mux_v
    port map (
            O => \N__46278\,
            I => \N__46160\
        );

    \I__10524\ : Span4Mux_h
    port map (
            O => \N__46275\,
            I => \N__46160\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__46272\,
            I => \N__46160\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__46269\,
            I => \N__46152\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__46262\,
            I => \N__46152\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__46259\,
            I => \N__46152\
        );

    \I__10519\ : InMux
    port map (
            O => \N__46258\,
            I => \N__46149\
        );

    \I__10518\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46146\
        );

    \I__10517\ : InMux
    port map (
            O => \N__46256\,
            I => \N__46143\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__46249\,
            I => \N__46132\
        );

    \I__10515\ : Span4Mux_v
    port map (
            O => \N__46244\,
            I => \N__46132\
        );

    \I__10514\ : Span4Mux_v
    port map (
            O => \N__46241\,
            I => \N__46132\
        );

    \I__10513\ : Span4Mux_v
    port map (
            O => \N__46238\,
            I => \N__46132\
        );

    \I__10512\ : Span4Mux_h
    port map (
            O => \N__46225\,
            I => \N__46132\
        );

    \I__10511\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46129\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__46221\,
            I => \N__46122\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__46218\,
            I => \N__46122\
        );

    \I__10508\ : Span4Mux_v
    port map (
            O => \N__46215\,
            I => \N__46122\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__46210\,
            I => \N__46111\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__46203\,
            I => \N__46111\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__46200\,
            I => \N__46111\
        );

    \I__10504\ : Span4Mux_v
    port map (
            O => \N__46197\,
            I => \N__46111\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__46186\,
            I => \N__46111\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__46183\,
            I => \N__46098\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__46178\,
            I => \N__46098\
        );

    \I__10500\ : Span4Mux_v
    port map (
            O => \N__46175\,
            I => \N__46098\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__46172\,
            I => \N__46098\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__46169\,
            I => \N__46098\
        );

    \I__10497\ : Span4Mux_v
    port map (
            O => \N__46160\,
            I => \N__46098\
        );

    \I__10496\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46095\
        );

    \I__10495\ : Span12Mux_h
    port map (
            O => \N__46152\,
            I => \N__46092\
        );

    \I__10494\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46089\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__46146\,
            I => \N__46084\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__46143\,
            I => \N__46084\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__46132\,
            I => \N__46081\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__46129\,
            I => \N__46072\
        );

    \I__10489\ : Span4Mux_v
    port map (
            O => \N__46122\,
            I => \N__46072\
        );

    \I__10488\ : Span4Mux_v
    port map (
            O => \N__46111\,
            I => \N__46072\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__46098\,
            I => \N__46072\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__46095\,
            I => comm_cmd_1
        );

    \I__10485\ : Odrv12
    port map (
            O => \N__46092\,
            I => comm_cmd_1
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__46089\,
            I => comm_cmd_1
        );

    \I__10483\ : Odrv4
    port map (
            O => \N__46084\,
            I => comm_cmd_1
        );

    \I__10482\ : Odrv4
    port map (
            O => \N__46081\,
            I => comm_cmd_1
        );

    \I__10481\ : Odrv4
    port map (
            O => \N__46072\,
            I => comm_cmd_1
        );

    \I__10480\ : SRMux
    port map (
            O => \N__46059\,
            I => \N__46056\
        );

    \I__10479\ : LocalMux
    port map (
            O => \N__46056\,
            I => \N__46053\
        );

    \I__10478\ : Span4Mux_v
    port map (
            O => \N__46053\,
            I => \N__46050\
        );

    \I__10477\ : Odrv4
    port map (
            O => \N__46050\,
            I => n16824
        );

    \I__10476\ : InMux
    port map (
            O => \N__46047\,
            I => \N__46044\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__46044\,
            I => \N__46041\
        );

    \I__10474\ : Odrv4
    port map (
            O => \N__46041\,
            I => comm_length_1
        );

    \I__10473\ : InMux
    port map (
            O => \N__46038\,
            I => \N__46033\
        );

    \I__10472\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46030\
        );

    \I__10471\ : InMux
    port map (
            O => \N__46036\,
            I => \N__46027\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__46033\,
            I => \N__46024\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__46030\,
            I => \N__46021\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__46018\
        );

    \I__10467\ : Span4Mux_h
    port map (
            O => \N__46024\,
            I => \N__46015\
        );

    \I__10466\ : Span12Mux_v
    port map (
            O => \N__46021\,
            I => \N__46010\
        );

    \I__10465\ : Span12Mux_h
    port map (
            O => \N__46018\,
            I => \N__46010\
        );

    \I__10464\ : Odrv4
    port map (
            O => \N__46015\,
            I => n5_adj_1524
        );

    \I__10463\ : Odrv12
    port map (
            O => \N__46010\,
            I => n5_adj_1524
        );

    \I__10462\ : InMux
    port map (
            O => \N__46005\,
            I => \N__46002\
        );

    \I__10461\ : LocalMux
    port map (
            O => \N__46002\,
            I => \N__45999\
        );

    \I__10460\ : Span4Mux_h
    port map (
            O => \N__45999\,
            I => \N__45996\
        );

    \I__10459\ : Span4Mux_h
    port map (
            O => \N__45996\,
            I => \N__45993\
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__45993\,
            I => n30_adj_1605
        );

    \I__10457\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45987\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__45987\,
            I => \N__45984\
        );

    \I__10455\ : Span4Mux_v
    port map (
            O => \N__45984\,
            I => \N__45981\
        );

    \I__10454\ : Sp12to4
    port map (
            O => \N__45981\,
            I => \N__45978\
        );

    \I__10453\ : Odrv12
    port map (
            O => \N__45978\,
            I => n30_adj_1608
        );

    \I__10452\ : CascadeMux
    port map (
            O => \N__45975\,
            I => \N__45972\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45969\
        );

    \I__10450\ : LocalMux
    port map (
            O => \N__45969\,
            I => \N__45966\
        );

    \I__10449\ : Odrv4
    port map (
            O => \N__45966\,
            I => comm_buf_2_4
        );

    \I__10448\ : InMux
    port map (
            O => \N__45963\,
            I => \N__45960\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__45960\,
            I => \N__45957\
        );

    \I__10446\ : Span4Mux_v
    port map (
            O => \N__45957\,
            I => \N__45954\
        );

    \I__10445\ : Span4Mux_h
    port map (
            O => \N__45954\,
            I => \N__45951\
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__45951\,
            I => n30_adj_1611
        );

    \I__10443\ : InMux
    port map (
            O => \N__45948\,
            I => \N__45945\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45945\,
            I => \N__45942\
        );

    \I__10441\ : Odrv4
    port map (
            O => \N__45942\,
            I => comm_buf_2_3
        );

    \I__10440\ : InMux
    port map (
            O => \N__45939\,
            I => \N__45936\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__45936\,
            I => \N__45933\
        );

    \I__10438\ : Span12Mux_v
    port map (
            O => \N__45933\,
            I => \N__45930\
        );

    \I__10437\ : Odrv12
    port map (
            O => \N__45930\,
            I => n30_adj_1614
        );

    \I__10436\ : InMux
    port map (
            O => \N__45927\,
            I => \N__45924\
        );

    \I__10435\ : LocalMux
    port map (
            O => \N__45924\,
            I => \N__45921\
        );

    \I__10434\ : Odrv12
    port map (
            O => \N__45921\,
            I => comm_buf_2_2
        );

    \I__10433\ : InMux
    port map (
            O => \N__45918\,
            I => \N__45915\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45915\,
            I => \N__45912\
        );

    \I__10431\ : Span4Mux_h
    port map (
            O => \N__45912\,
            I => \N__45909\
        );

    \I__10430\ : Odrv4
    port map (
            O => \N__45909\,
            I => n30_adj_1618
        );

    \I__10429\ : CEMux
    port map (
            O => \N__45906\,
            I => \N__45903\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45903\,
            I => \N__45899\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45896\
        );

    \I__10426\ : Odrv4
    port map (
            O => \N__45899\,
            I => n12314
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__45896\,
            I => n12314
        );

    \I__10424\ : SRMux
    port map (
            O => \N__45891\,
            I => \N__45888\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45885\
        );

    \I__10422\ : Span4Mux_h
    port map (
            O => \N__45885\,
            I => \N__45882\
        );

    \I__10421\ : Odrv4
    port map (
            O => \N__45882\,
            I => n14972
        );

    \I__10420\ : CascadeMux
    port map (
            O => \N__45879\,
            I => \N__45875\
        );

    \I__10419\ : CascadeMux
    port map (
            O => \N__45878\,
            I => \N__45871\
        );

    \I__10418\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45865\
        );

    \I__10417\ : CascadeMux
    port map (
            O => \N__45874\,
            I => \N__45861\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45858\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45855\
        );

    \I__10414\ : CascadeMux
    port map (
            O => \N__45869\,
            I => \N__45852\
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__45868\,
            I => \N__45849\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__45865\,
            I => \N__45845\
        );

    \I__10411\ : CascadeMux
    port map (
            O => \N__45864\,
            I => \N__45842\
        );

    \I__10410\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45839\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__45858\,
            I => \N__45836\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__45855\,
            I => \N__45833\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45852\,
            I => \N__45830\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45849\,
            I => \N__45824\
        );

    \I__10405\ : InMux
    port map (
            O => \N__45848\,
            I => \N__45824\
        );

    \I__10404\ : Span4Mux_h
    port map (
            O => \N__45845\,
            I => \N__45821\
        );

    \I__10403\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45818\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__45839\,
            I => \N__45809\
        );

    \I__10401\ : Span4Mux_v
    port map (
            O => \N__45836\,
            I => \N__45809\
        );

    \I__10400\ : Span4Mux_h
    port map (
            O => \N__45833\,
            I => \N__45809\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__45830\,
            I => \N__45809\
        );

    \I__10398\ : InMux
    port map (
            O => \N__45829\,
            I => \N__45806\
        );

    \I__10397\ : LocalMux
    port map (
            O => \N__45824\,
            I => \N__45803\
        );

    \I__10396\ : Span4Mux_v
    port map (
            O => \N__45821\,
            I => \N__45800\
        );

    \I__10395\ : LocalMux
    port map (
            O => \N__45818\,
            I => \N__45797\
        );

    \I__10394\ : Span4Mux_h
    port map (
            O => \N__45809\,
            I => \N__45794\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__45806\,
            I => \N__45791\
        );

    \I__10392\ : Span4Mux_h
    port map (
            O => \N__45803\,
            I => \N__45788\
        );

    \I__10391\ : Sp12to4
    port map (
            O => \N__45800\,
            I => \N__45785\
        );

    \I__10390\ : Span4Mux_h
    port map (
            O => \N__45797\,
            I => \N__45782\
        );

    \I__10389\ : Span4Mux_h
    port map (
            O => \N__45794\,
            I => \N__45775\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__45791\,
            I => \N__45775\
        );

    \I__10387\ : Span4Mux_h
    port map (
            O => \N__45788\,
            I => \N__45775\
        );

    \I__10386\ : Odrv12
    port map (
            O => \N__45785\,
            I => comm_buf_0_2
        );

    \I__10385\ : Odrv4
    port map (
            O => \N__45782\,
            I => comm_buf_0_2
        );

    \I__10384\ : Odrv4
    port map (
            O => \N__45775\,
            I => comm_buf_0_2
        );

    \I__10383\ : InMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__10382\ : LocalMux
    port map (
            O => \N__45765\,
            I => \N__45762\
        );

    \I__10381\ : Span4Mux_v
    port map (
            O => \N__45762\,
            I => \N__45759\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__45759\,
            I => \N__45756\
        );

    \I__10379\ : Odrv4
    port map (
            O => \N__45756\,
            I => buf_data_iac_19
        );

    \I__10378\ : InMux
    port map (
            O => \N__45753\,
            I => \N__45750\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45747\
        );

    \I__10376\ : Span4Mux_h
    port map (
            O => \N__45747\,
            I => \N__45744\
        );

    \I__10375\ : Span4Mux_h
    port map (
            O => \N__45744\,
            I => \N__45741\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45741\,
            I => n21543
        );

    \I__10373\ : IoInMux
    port map (
            O => \N__45738\,
            I => \N__45735\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45735\,
            I => \N__45732\
        );

    \I__10371\ : IoSpan4Mux
    port map (
            O => \N__45732\,
            I => \N__45729\
        );

    \I__10370\ : Span4Mux_s3_v
    port map (
            O => \N__45729\,
            I => \N__45725\
        );

    \I__10369\ : InMux
    port map (
            O => \N__45728\,
            I => \N__45722\
        );

    \I__10368\ : Sp12to4
    port map (
            O => \N__45725\,
            I => \N__45719\
        );

    \I__10367\ : LocalMux
    port map (
            O => \N__45722\,
            I => \N__45715\
        );

    \I__10366\ : Span12Mux_s11_v
    port map (
            O => \N__45719\,
            I => \N__45712\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45718\,
            I => \N__45709\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__45715\,
            I => \N__45706\
        );

    \I__10363\ : Odrv12
    port map (
            O => \N__45712\,
            I => \SELIRNG0\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__45709\,
            I => \SELIRNG0\
        );

    \I__10361\ : Odrv4
    port map (
            O => \N__45706\,
            I => \SELIRNG0\
        );

    \I__10360\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45696\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__10358\ : Span4Mux_h
    port map (
            O => \N__45693\,
            I => \N__45690\
        );

    \I__10357\ : Odrv4
    port map (
            O => \N__45690\,
            I => n23_adj_1685
        );

    \I__10356\ : InMux
    port map (
            O => \N__45687\,
            I => \N__45684\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__45684\,
            I => n21273
        );

    \I__10354\ : InMux
    port map (
            O => \N__45681\,
            I => \N__45678\
        );

    \I__10353\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45674\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45671\
        );

    \I__10351\ : Span4Mux_h
    port map (
            O => \N__45674\,
            I => \N__45666\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45671\,
            I => \N__45663\
        );

    \I__10349\ : InMux
    port map (
            O => \N__45670\,
            I => \N__45658\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45669\,
            I => \N__45658\
        );

    \I__10347\ : Odrv4
    port map (
            O => \N__45666\,
            I => comm_buf_1_0
        );

    \I__10346\ : Odrv4
    port map (
            O => \N__45663\,
            I => comm_buf_1_0
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__45658\,
            I => comm_buf_1_0
        );

    \I__10344\ : CascadeMux
    port map (
            O => \N__45651\,
            I => \n22533_cascade_\
        );

    \I__10343\ : InMux
    port map (
            O => \N__45648\,
            I => \N__45642\
        );

    \I__10342\ : CascadeMux
    port map (
            O => \N__45647\,
            I => \N__45639\
        );

    \I__10341\ : CascadeMux
    port map (
            O => \N__45646\,
            I => \N__45636\
        );

    \I__10340\ : CascadeMux
    port map (
            O => \N__45645\,
            I => \N__45631\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__45642\,
            I => \N__45628\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45625\
        );

    \I__10337\ : InMux
    port map (
            O => \N__45636\,
            I => \N__45622\
        );

    \I__10336\ : CascadeMux
    port map (
            O => \N__45635\,
            I => \N__45617\
        );

    \I__10335\ : InMux
    port map (
            O => \N__45634\,
            I => \N__45613\
        );

    \I__10334\ : InMux
    port map (
            O => \N__45631\,
            I => \N__45610\
        );

    \I__10333\ : Span4Mux_h
    port map (
            O => \N__45628\,
            I => \N__45605\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__45625\,
            I => \N__45605\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__45622\,
            I => \N__45602\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45599\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45620\,
            I => \N__45596\
        );

    \I__10328\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45593\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45616\,
            I => \N__45590\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45613\,
            I => \N__45585\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45585\
        );

    \I__10324\ : Span4Mux_v
    port map (
            O => \N__45605\,
            I => \N__45582\
        );

    \I__10323\ : Span4Mux_v
    port map (
            O => \N__45602\,
            I => \N__45579\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__45599\,
            I => \N__45576\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__45596\,
            I => \N__45573\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45593\,
            I => \N__45568\
        );

    \I__10319\ : LocalMux
    port map (
            O => \N__45590\,
            I => \N__45568\
        );

    \I__10318\ : Span4Mux_v
    port map (
            O => \N__45585\,
            I => \N__45563\
        );

    \I__10317\ : Span4Mux_h
    port map (
            O => \N__45582\,
            I => \N__45563\
        );

    \I__10316\ : Span4Mux_h
    port map (
            O => \N__45579\,
            I => \N__45554\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__45576\,
            I => \N__45554\
        );

    \I__10314\ : Span4Mux_v
    port map (
            O => \N__45573\,
            I => \N__45554\
        );

    \I__10313\ : Span4Mux_v
    port map (
            O => \N__45568\,
            I => \N__45554\
        );

    \I__10312\ : Odrv4
    port map (
            O => \N__45563\,
            I => comm_buf_0_0
        );

    \I__10311\ : Odrv4
    port map (
            O => \N__45554\,
            I => comm_buf_0_0
        );

    \I__10310\ : InMux
    port map (
            O => \N__45549\,
            I => \N__45546\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__45546\,
            I => n22536
        );

    \I__10308\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45540\
        );

    \I__10307\ : LocalMux
    port map (
            O => \N__45540\,
            I => n24_adj_1639
        );

    \I__10306\ : CascadeMux
    port map (
            O => \N__45537\,
            I => \n21497_cascade_\
        );

    \I__10305\ : CascadeMux
    port map (
            O => \N__45534\,
            I => \n34_adj_1649_cascade_\
        );

    \I__10304\ : InMux
    port map (
            O => \N__45531\,
            I => \N__45528\
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__45528\,
            I => n30_adj_1531
        );

    \I__10302\ : InMux
    port map (
            O => \N__45525\,
            I => \N__45522\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__45522\,
            I => comm_buf_2_0
        );

    \I__10300\ : InMux
    port map (
            O => \N__45519\,
            I => \N__45516\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__45516\,
            I => \N__45513\
        );

    \I__10298\ : Span12Mux_h
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__10297\ : Odrv12
    port map (
            O => \N__45510\,
            I => n30_adj_1599
        );

    \I__10296\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45504\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__45504\,
            I => comm_buf_2_7
        );

    \I__10294\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45498\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__45498\,
            I => \N__45495\
        );

    \I__10292\ : Span4Mux_h
    port map (
            O => \N__45495\,
            I => \N__45492\
        );

    \I__10291\ : Span4Mux_h
    port map (
            O => \N__45492\,
            I => \N__45489\
        );

    \I__10290\ : Span4Mux_h
    port map (
            O => \N__45489\,
            I => \N__45486\
        );

    \I__10289\ : Span4Mux_v
    port map (
            O => \N__45486\,
            I => \N__45483\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__45483\,
            I => n30_adj_1602
        );

    \I__10287\ : CascadeMux
    port map (
            O => \N__45480\,
            I => \N__45476\
        );

    \I__10286\ : InMux
    port map (
            O => \N__45479\,
            I => \N__45472\
        );

    \I__10285\ : InMux
    port map (
            O => \N__45476\,
            I => \N__45469\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45466\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__45472\,
            I => \N__45462\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__45469\,
            I => \N__45459\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__45466\,
            I => \N__45456\
        );

    \I__10280\ : InMux
    port map (
            O => \N__45465\,
            I => \N__45453\
        );

    \I__10279\ : Span4Mux_h
    port map (
            O => \N__45462\,
            I => \N__45450\
        );

    \I__10278\ : Span4Mux_h
    port map (
            O => \N__45459\,
            I => \N__45445\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__45456\,
            I => \N__45445\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__45453\,
            I => \N__45442\
        );

    \I__10275\ : Span4Mux_v
    port map (
            O => \N__45450\,
            I => \N__45439\
        );

    \I__10274\ : Span4Mux_h
    port map (
            O => \N__45445\,
            I => \N__45434\
        );

    \I__10273\ : Span4Mux_h
    port map (
            O => \N__45442\,
            I => \N__45434\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__45439\,
            I => \N__45431\
        );

    \I__10271\ : Span4Mux_v
    port map (
            O => \N__45434\,
            I => \N__45428\
        );

    \I__10270\ : Odrv4
    port map (
            O => \N__45431\,
            I => comm_buf_1_2
        );

    \I__10269\ : Odrv4
    port map (
            O => \N__45428\,
            I => comm_buf_1_2
        );

    \I__10268\ : CascadeMux
    port map (
            O => \N__45423\,
            I => \n1_cascade_\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45420\,
            I => \N__45417\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__45417\,
            I => n2_adj_1584
        );

    \I__10265\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45411\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__45411\,
            I => \N__45408\
        );

    \I__10263\ : Odrv12
    port map (
            O => \N__45408\,
            I => comm_buf_4_2
        );

    \I__10262\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45402\
        );

    \I__10261\ : LocalMux
    port map (
            O => \N__45402\,
            I => n21528
        );

    \I__10260\ : CascadeMux
    port map (
            O => \N__45399\,
            I => \n4_adj_1585_cascade_\
        );

    \I__10259\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45393\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__45393\,
            I => n22491
        );

    \I__10257\ : CascadeMux
    port map (
            O => \N__45390\,
            I => \N__45385\
        );

    \I__10256\ : InMux
    port map (
            O => \N__45389\,
            I => \N__45382\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45388\,
            I => \N__45377\
        );

    \I__10254\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45377\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__45382\,
            I => \N__45374\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__45377\,
            I => \N__45371\
        );

    \I__10251\ : Span4Mux_v
    port map (
            O => \N__45374\,
            I => \N__45366\
        );

    \I__10250\ : Span4Mux_h
    port map (
            O => \N__45371\,
            I => \N__45366\
        );

    \I__10249\ : Odrv4
    port map (
            O => \N__45366\,
            I => n21143
        );

    \I__10248\ : CascadeMux
    port map (
            O => \N__45363\,
            I => \n19193_cascade_\
        );

    \I__10247\ : CascadeMux
    port map (
            O => \N__45360\,
            I => \n19188_cascade_\
        );

    \I__10246\ : CascadeMux
    port map (
            O => \N__45357\,
            I => \N__45353\
        );

    \I__10245\ : CascadeMux
    port map (
            O => \N__45356\,
            I => \N__45349\
        );

    \I__10244\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45345\
        );

    \I__10243\ : InMux
    port map (
            O => \N__45352\,
            I => \N__45342\
        );

    \I__10242\ : InMux
    port map (
            O => \N__45349\,
            I => \N__45339\
        );

    \I__10241\ : InMux
    port map (
            O => \N__45348\,
            I => \N__45336\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__45345\,
            I => \N__45327\
        );

    \I__10239\ : LocalMux
    port map (
            O => \N__45342\,
            I => \N__45327\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__45339\,
            I => \N__45327\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__45336\,
            I => \N__45323\
        );

    \I__10236\ : InMux
    port map (
            O => \N__45335\,
            I => \N__45320\
        );

    \I__10235\ : InMux
    port map (
            O => \N__45334\,
            I => \N__45317\
        );

    \I__10234\ : Span4Mux_v
    port map (
            O => \N__45327\,
            I => \N__45314\
        );

    \I__10233\ : InMux
    port map (
            O => \N__45326\,
            I => \N__45311\
        );

    \I__10232\ : Span4Mux_h
    port map (
            O => \N__45323\,
            I => \N__45306\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__45320\,
            I => \N__45306\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__45317\,
            I => \N__45303\
        );

    \I__10229\ : Span4Mux_h
    port map (
            O => \N__45314\,
            I => \N__45293\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__45311\,
            I => \N__45293\
        );

    \I__10227\ : Span4Mux_h
    port map (
            O => \N__45306\,
            I => \N__45293\
        );

    \I__10226\ : Span4Mux_h
    port map (
            O => \N__45303\,
            I => \N__45293\
        );

    \I__10225\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45290\
        );

    \I__10224\ : Odrv4
    port map (
            O => \N__45293\,
            I => comm_buf_0_3
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__45290\,
            I => comm_buf_0_3
        );

    \I__10222\ : CascadeMux
    port map (
            O => \N__45285\,
            I => \n22557_cascade_\
        );

    \I__10221\ : InMux
    port map (
            O => \N__45282\,
            I => \N__45275\
        );

    \I__10220\ : InMux
    port map (
            O => \N__45281\,
            I => \N__45275\
        );

    \I__10219\ : InMux
    port map (
            O => \N__45280\,
            I => \N__45272\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__45275\,
            I => \N__45269\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__45272\,
            I => \N__45266\
        );

    \I__10216\ : Span4Mux_h
    port map (
            O => \N__45269\,
            I => \N__45263\
        );

    \I__10215\ : Span4Mux_h
    port map (
            O => \N__45266\,
            I => \N__45260\
        );

    \I__10214\ : Span4Mux_h
    port map (
            O => \N__45263\,
            I => \N__45257\
        );

    \I__10213\ : Odrv4
    port map (
            O => \N__45260\,
            I => comm_buf_1_3
        );

    \I__10212\ : Odrv4
    port map (
            O => \N__45257\,
            I => comm_buf_1_3
        );

    \I__10211\ : InMux
    port map (
            O => \N__45252\,
            I => \N__45249\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__45249\,
            I => \N__45246\
        );

    \I__10209\ : Odrv12
    port map (
            O => \N__45246\,
            I => comm_buf_4_3
        );

    \I__10208\ : CascadeMux
    port map (
            O => \N__45243\,
            I => \n4_adj_1583_cascade_\
        );

    \I__10207\ : InMux
    port map (
            O => \N__45240\,
            I => \N__45237\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__45237\,
            I => n22560
        );

    \I__10205\ : CascadeMux
    port map (
            O => \N__45234\,
            I => \n21288_cascade_\
        );

    \I__10204\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45228\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__45228\,
            I => \N__45225\
        );

    \I__10202\ : Span4Mux_h
    port map (
            O => \N__45225\,
            I => \N__45222\
        );

    \I__10201\ : Odrv4
    port map (
            O => \N__45222\,
            I => n21479
        );

    \I__10200\ : CascadeMux
    port map (
            O => \N__45219\,
            I => \n21477_cascade_\
        );

    \I__10199\ : CascadeMux
    port map (
            O => \N__45216\,
            I => \n44_cascade_\
        );

    \I__10198\ : CEMux
    port map (
            O => \N__45213\,
            I => \N__45206\
        );

    \I__10197\ : CEMux
    port map (
            O => \N__45212\,
            I => \N__45203\
        );

    \I__10196\ : CEMux
    port map (
            O => \N__45211\,
            I => \N__45200\
        );

    \I__10195\ : CEMux
    port map (
            O => \N__45210\,
            I => \N__45196\
        );

    \I__10194\ : CEMux
    port map (
            O => \N__45209\,
            I => \N__45191\
        );

    \I__10193\ : LocalMux
    port map (
            O => \N__45206\,
            I => \N__45186\
        );

    \I__10192\ : LocalMux
    port map (
            O => \N__45203\,
            I => \N__45186\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__45200\,
            I => \N__45183\
        );

    \I__10190\ : CEMux
    port map (
            O => \N__45199\,
            I => \N__45180\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__45196\,
            I => \N__45177\
        );

    \I__10188\ : CEMux
    port map (
            O => \N__45195\,
            I => \N__45174\
        );

    \I__10187\ : CEMux
    port map (
            O => \N__45194\,
            I => \N__45171\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__45191\,
            I => \N__45167\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__45186\,
            I => \N__45164\
        );

    \I__10184\ : Span4Mux_v
    port map (
            O => \N__45183\,
            I => \N__45157\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__45180\,
            I => \N__45157\
        );

    \I__10182\ : Span4Mux_v
    port map (
            O => \N__45177\,
            I => \N__45157\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__45174\,
            I => \N__45154\
        );

    \I__10180\ : LocalMux
    port map (
            O => \N__45171\,
            I => \N__45151\
        );

    \I__10179\ : InMux
    port map (
            O => \N__45170\,
            I => \N__45148\
        );

    \I__10178\ : Span4Mux_h
    port map (
            O => \N__45167\,
            I => \N__45145\
        );

    \I__10177\ : Span4Mux_h
    port map (
            O => \N__45164\,
            I => \N__45140\
        );

    \I__10176\ : Span4Mux_v
    port map (
            O => \N__45157\,
            I => \N__45140\
        );

    \I__10175\ : Span4Mux_h
    port map (
            O => \N__45154\,
            I => \N__45133\
        );

    \I__10174\ : Span4Mux_v
    port map (
            O => \N__45151\,
            I => \N__45133\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__45148\,
            I => \N__45133\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__45145\,
            I => n12260
        );

    \I__10171\ : Odrv4
    port map (
            O => \N__45140\,
            I => n12260
        );

    \I__10170\ : Odrv4
    port map (
            O => \N__45133\,
            I => n12260
        );

    \I__10169\ : InMux
    port map (
            O => \N__45126\,
            I => \N__45123\
        );

    \I__10168\ : LocalMux
    port map (
            O => \N__45123\,
            I => \N__45120\
        );

    \I__10167\ : Span4Mux_h
    port map (
            O => \N__45120\,
            I => \N__45117\
        );

    \I__10166\ : Span4Mux_v
    port map (
            O => \N__45117\,
            I => \N__45114\
        );

    \I__10165\ : Span4Mux_v
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__10164\ : Odrv4
    port map (
            O => \N__45111\,
            I => buf_data_vac_10
        );

    \I__10163\ : InMux
    port map (
            O => \N__45108\,
            I => \N__45105\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__10161\ : Span4Mux_h
    port map (
            O => \N__45102\,
            I => \N__45099\
        );

    \I__10160\ : Span4Mux_v
    port map (
            O => \N__45099\,
            I => \N__45096\
        );

    \I__10159\ : Span4Mux_v
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__10158\ : Odrv4
    port map (
            O => \N__45093\,
            I => buf_data_vac_9
        );

    \I__10157\ : SRMux
    port map (
            O => \N__45090\,
            I => \N__45087\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__45087\,
            I => \N__45084\
        );

    \I__10155\ : Span4Mux_h
    port map (
            O => \N__45084\,
            I => \N__45081\
        );

    \I__10154\ : Odrv4
    port map (
            O => \N__45081\,
            I => n14986
        );

    \I__10153\ : CascadeMux
    port map (
            O => \N__45078\,
            I => \n21268_cascade_\
        );

    \I__10152\ : InMux
    port map (
            O => \N__45075\,
            I => \N__45072\
        );

    \I__10151\ : LocalMux
    port map (
            O => \N__45072\,
            I => n22094
        );

    \I__10150\ : CascadeMux
    port map (
            O => \N__45069\,
            I => \N__45066\
        );

    \I__10149\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45063\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__45063\,
            I => n21266
        );

    \I__10147\ : CEMux
    port map (
            O => \N__45060\,
            I => \N__45056\
        );

    \I__10146\ : InMux
    port map (
            O => \N__45059\,
            I => \N__45053\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__45056\,
            I => \N__45050\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__45053\,
            I => \N__45047\
        );

    \I__10143\ : Odrv12
    port map (
            O => \N__45050\,
            I => n12407
        );

    \I__10142\ : Odrv4
    port map (
            O => \N__45047\,
            I => n12407
        );

    \I__10141\ : CascadeMux
    port map (
            O => \N__45042\,
            I => \n21085_cascade_\
        );

    \I__10140\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45036\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__45036\,
            I => n19188
        );

    \I__10138\ : InMux
    port map (
            O => \N__45033\,
            I => \N__45029\
        );

    \I__10137\ : InMux
    port map (
            O => \N__45032\,
            I => \N__45026\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__45029\,
            I => \N__45020\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__45026\,
            I => \N__45020\
        );

    \I__10134\ : InMux
    port map (
            O => \N__45025\,
            I => \N__45017\
        );

    \I__10133\ : Span4Mux_v
    port map (
            O => \N__45020\,
            I => \N__45011\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__45017\,
            I => \N__45011\
        );

    \I__10131\ : InMux
    port map (
            O => \N__45016\,
            I => \N__45008\
        );

    \I__10130\ : Span4Mux_h
    port map (
            O => \N__45011\,
            I => \N__45005\
        );

    \I__10129\ : LocalMux
    port map (
            O => \N__45008\,
            I => \comm_spi.n23092\
        );

    \I__10128\ : Odrv4
    port map (
            O => \N__45005\,
            I => \comm_spi.n23092\
        );

    \I__10127\ : InMux
    port map (
            O => \N__45000\,
            I => \N__44997\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__44997\,
            I => \N__44994\
        );

    \I__10125\ : Span4Mux_v
    port map (
            O => \N__44994\,
            I => \N__44989\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44993\,
            I => \N__44986\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44992\,
            I => \N__44983\
        );

    \I__10122\ : Odrv4
    port map (
            O => \N__44989\,
            I => clk_cnt_1
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44986\,
            I => clk_cnt_1
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__44983\,
            I => clk_cnt_1
        );

    \I__10119\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44973\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44973\,
            I => \N__44970\
        );

    \I__10117\ : Span4Mux_v
    port map (
            O => \N__44970\,
            I => \N__44964\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44959\
        );

    \I__10115\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44959\
        );

    \I__10114\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44956\
        );

    \I__10113\ : Odrv4
    port map (
            O => \N__44964\,
            I => clk_cnt_0
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__44959\,
            I => clk_cnt_0
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__44956\,
            I => clk_cnt_0
        );

    \I__10110\ : SRMux
    port map (
            O => \N__44949\,
            I => \N__44946\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44946\,
            I => \N__44943\
        );

    \I__10108\ : Odrv4
    port map (
            O => \N__44943\,
            I => n17773
        );

    \I__10107\ : InMux
    port map (
            O => \N__44940\,
            I => \N__44937\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44934\
        );

    \I__10105\ : Span4Mux_h
    port map (
            O => \N__44934\,
            I => \N__44931\
        );

    \I__10104\ : Span4Mux_v
    port map (
            O => \N__44931\,
            I => \N__44928\
        );

    \I__10103\ : Sp12to4
    port map (
            O => \N__44928\,
            I => \N__44925\
        );

    \I__10102\ : Odrv12
    port map (
            O => \N__44925\,
            I => buf_data_vac_8
        );

    \I__10101\ : InMux
    port map (
            O => \N__44922\,
            I => \N__44919\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44919\,
            I => \N__44916\
        );

    \I__10099\ : Span4Mux_h
    port map (
            O => \N__44916\,
            I => \N__44913\
        );

    \I__10098\ : Span4Mux_v
    port map (
            O => \N__44913\,
            I => \N__44910\
        );

    \I__10097\ : Odrv4
    port map (
            O => \N__44910\,
            I => buf_data_vac_15
        );

    \I__10096\ : InMux
    port map (
            O => \N__44907\,
            I => \N__44904\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__44904\,
            I => comm_buf_4_7
        );

    \I__10094\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44898\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44898\,
            I => \N__44895\
        );

    \I__10092\ : Span12Mux_h
    port map (
            O => \N__44895\,
            I => \N__44892\
        );

    \I__10091\ : Odrv12
    port map (
            O => \N__44892\,
            I => buf_data_vac_14
        );

    \I__10090\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44886\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44886\,
            I => \N__44883\
        );

    \I__10088\ : Span4Mux_h
    port map (
            O => \N__44883\,
            I => \N__44880\
        );

    \I__10087\ : Span4Mux_v
    port map (
            O => \N__44880\,
            I => \N__44877\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__44877\,
            I => buf_data_vac_13
        );

    \I__10085\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44871\
        );

    \I__10084\ : LocalMux
    port map (
            O => \N__44871\,
            I => \N__44868\
        );

    \I__10083\ : Span4Mux_h
    port map (
            O => \N__44868\,
            I => \N__44865\
        );

    \I__10082\ : Span4Mux_v
    port map (
            O => \N__44865\,
            I => \N__44862\
        );

    \I__10081\ : Span4Mux_v
    port map (
            O => \N__44862\,
            I => \N__44859\
        );

    \I__10080\ : Odrv4
    port map (
            O => \N__44859\,
            I => buf_data_vac_12
        );

    \I__10079\ : InMux
    port map (
            O => \N__44856\,
            I => \N__44853\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__44853\,
            I => \N__44850\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__44850\,
            I => comm_buf_4_4
        );

    \I__10076\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44844\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44844\,
            I => \N__44841\
        );

    \I__10074\ : Span4Mux_v
    port map (
            O => \N__44841\,
            I => \N__44838\
        );

    \I__10073\ : Span4Mux_v
    port map (
            O => \N__44838\,
            I => \N__44835\
        );

    \I__10072\ : Span4Mux_h
    port map (
            O => \N__44835\,
            I => \N__44832\
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__44832\,
            I => buf_data_vac_11
        );

    \I__10070\ : InMux
    port map (
            O => \N__44829\,
            I => \N__44826\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__44826\,
            I => \N__44823\
        );

    \I__10068\ : Span4Mux_v
    port map (
            O => \N__44823\,
            I => \N__44819\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44822\,
            I => \N__44816\
        );

    \I__10066\ : Span4Mux_v
    port map (
            O => \N__44819\,
            I => \N__44810\
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__44816\,
            I => \N__44810\
        );

    \I__10064\ : InMux
    port map (
            O => \N__44815\,
            I => \N__44807\
        );

    \I__10063\ : Span4Mux_v
    port map (
            O => \N__44810\,
            I => \N__44804\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__44807\,
            I => wdtick_flag
        );

    \I__10061\ : Odrv4
    port map (
            O => \N__44804\,
            I => wdtick_flag
        );

    \I__10060\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44796\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44793\
        );

    \I__10058\ : Span4Mux_v
    port map (
            O => \N__44793\,
            I => \N__44788\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44792\,
            I => \N__44785\
        );

    \I__10056\ : InMux
    port map (
            O => \N__44791\,
            I => \N__44782\
        );

    \I__10055\ : Odrv4
    port map (
            O => \N__44788\,
            I => buf_control_0
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__44785\,
            I => buf_control_0
        );

    \I__10053\ : LocalMux
    port map (
            O => \N__44782\,
            I => buf_control_0
        );

    \I__10052\ : IoInMux
    port map (
            O => \N__44775\,
            I => \N__44772\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44772\,
            I => \N__44769\
        );

    \I__10050\ : Span4Mux_s1_v
    port map (
            O => \N__44769\,
            I => \N__44766\
        );

    \I__10049\ : Span4Mux_h
    port map (
            O => \N__44766\,
            I => \N__44763\
        );

    \I__10048\ : Span4Mux_v
    port map (
            O => \N__44763\,
            I => \N__44760\
        );

    \I__10047\ : Span4Mux_v
    port map (
            O => \N__44760\,
            I => \N__44757\
        );

    \I__10046\ : Odrv4
    port map (
            O => \N__44757\,
            I => \CONT_SD\
        );

    \I__10045\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44749\
        );

    \I__10044\ : CascadeMux
    port map (
            O => \N__44753\,
            I => \N__44745\
        );

    \I__10043\ : InMux
    port map (
            O => \N__44752\,
            I => \N__44741\
        );

    \I__10042\ : LocalMux
    port map (
            O => \N__44749\,
            I => \N__44738\
        );

    \I__10041\ : InMux
    port map (
            O => \N__44748\,
            I => \N__44735\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44745\,
            I => \N__44730\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44744\,
            I => \N__44730\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44741\,
            I => \N__44727\
        );

    \I__10037\ : Span4Mux_v
    port map (
            O => \N__44738\,
            I => \N__44719\
        );

    \I__10036\ : LocalMux
    port map (
            O => \N__44735\,
            I => \N__44719\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44719\
        );

    \I__10034\ : Span4Mux_v
    port map (
            O => \N__44727\,
            I => \N__44716\
        );

    \I__10033\ : InMux
    port map (
            O => \N__44726\,
            I => \N__44713\
        );

    \I__10032\ : Span4Mux_h
    port map (
            O => \N__44719\,
            I => \N__44710\
        );

    \I__10031\ : Sp12to4
    port map (
            O => \N__44716\,
            I => \N__44703\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__44713\,
            I => \N__44703\
        );

    \I__10029\ : Span4Mux_h
    port map (
            O => \N__44710\,
            I => \N__44699\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44709\,
            I => \N__44696\
        );

    \I__10027\ : InMux
    port map (
            O => \N__44708\,
            I => \N__44693\
        );

    \I__10026\ : Span12Mux_v
    port map (
            O => \N__44703\,
            I => \N__44690\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44702\,
            I => \N__44687\
        );

    \I__10024\ : Span4Mux_v
    port map (
            O => \N__44699\,
            I => \N__44684\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__44696\,
            I => \N__44679\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__44693\,
            I => \N__44679\
        );

    \I__10021\ : Odrv12
    port map (
            O => \N__44690\,
            I => dds_state_0
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__44687\,
            I => dds_state_0
        );

    \I__10019\ : Odrv4
    port map (
            O => \N__44684\,
            I => dds_state_0
        );

    \I__10018\ : Odrv12
    port map (
            O => \N__44679\,
            I => dds_state_0
        );

    \I__10017\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44664\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44669\,
            I => \N__44661\
        );

    \I__10015\ : InMux
    port map (
            O => \N__44668\,
            I => \N__44658\
        );

    \I__10014\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44654\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44664\,
            I => \N__44633\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44661\,
            I => \N__44633\
        );

    \I__10011\ : LocalMux
    port map (
            O => \N__44658\,
            I => \N__44630\
        );

    \I__10010\ : InMux
    port map (
            O => \N__44657\,
            I => \N__44623\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__44654\,
            I => \N__44620\
        );

    \I__10008\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44617\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44602\
        );

    \I__10006\ : InMux
    port map (
            O => \N__44651\,
            I => \N__44602\
        );

    \I__10005\ : InMux
    port map (
            O => \N__44650\,
            I => \N__44602\
        );

    \I__10004\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44602\
        );

    \I__10003\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44602\
        );

    \I__10002\ : InMux
    port map (
            O => \N__44647\,
            I => \N__44602\
        );

    \I__10001\ : InMux
    port map (
            O => \N__44646\,
            I => \N__44602\
        );

    \I__10000\ : InMux
    port map (
            O => \N__44645\,
            I => \N__44585\
        );

    \I__9999\ : InMux
    port map (
            O => \N__44644\,
            I => \N__44585\
        );

    \I__9998\ : InMux
    port map (
            O => \N__44643\,
            I => \N__44585\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44642\,
            I => \N__44585\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44585\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44640\,
            I => \N__44585\
        );

    \I__9994\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44585\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44638\,
            I => \N__44585\
        );

    \I__9992\ : Span4Mux_h
    port map (
            O => \N__44633\,
            I => \N__44582\
        );

    \I__9991\ : Span4Mux_v
    port map (
            O => \N__44630\,
            I => \N__44579\
        );

    \I__9990\ : InMux
    port map (
            O => \N__44629\,
            I => \N__44570\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44628\,
            I => \N__44570\
        );

    \I__9988\ : InMux
    port map (
            O => \N__44627\,
            I => \N__44570\
        );

    \I__9987\ : InMux
    port map (
            O => \N__44626\,
            I => \N__44570\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__44623\,
            I => \N__44565\
        );

    \I__9985\ : Span12Mux_v
    port map (
            O => \N__44620\,
            I => \N__44565\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44617\,
            I => dds_state_2
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__44602\,
            I => dds_state_2
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__44585\,
            I => dds_state_2
        );

    \I__9981\ : Odrv4
    port map (
            O => \N__44582\,
            I => dds_state_2
        );

    \I__9980\ : Odrv4
    port map (
            O => \N__44579\,
            I => dds_state_2
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__44570\,
            I => dds_state_2
        );

    \I__9978\ : Odrv12
    port map (
            O => \N__44565\,
            I => dds_state_2
        );

    \I__9977\ : CEMux
    port map (
            O => \N__44550\,
            I => \N__44547\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__44547\,
            I => \N__44544\
        );

    \I__9975\ : Span4Mux_v
    port map (
            O => \N__44544\,
            I => \N__44540\
        );

    \I__9974\ : CEMux
    port map (
            O => \N__44543\,
            I => \N__44537\
        );

    \I__9973\ : Span4Mux_h
    port map (
            O => \N__44540\,
            I => \N__44534\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__44537\,
            I => \N__44531\
        );

    \I__9971\ : Span4Mux_h
    port map (
            O => \N__44534\,
            I => \N__44528\
        );

    \I__9970\ : Span4Mux_v
    port map (
            O => \N__44531\,
            I => \N__44525\
        );

    \I__9969\ : Span4Mux_v
    port map (
            O => \N__44528\,
            I => \N__44520\
        );

    \I__9968\ : Span4Mux_h
    port map (
            O => \N__44525\,
            I => \N__44520\
        );

    \I__9967\ : Odrv4
    port map (
            O => \N__44520\,
            I => \SIG_DDS.n9\
        );

    \I__9966\ : CEMux
    port map (
            O => \N__44517\,
            I => \N__44512\
        );

    \I__9965\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44509\
        );

    \I__9964\ : InMux
    port map (
            O => \N__44515\,
            I => \N__44505\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__44512\,
            I => \N__44500\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__44509\,
            I => \N__44488\
        );

    \I__9961\ : InMux
    port map (
            O => \N__44508\,
            I => \N__44485\
        );

    \I__9960\ : LocalMux
    port map (
            O => \N__44505\,
            I => \N__44482\
        );

    \I__9959\ : InMux
    port map (
            O => \N__44504\,
            I => \N__44479\
        );

    \I__9958\ : SRMux
    port map (
            O => \N__44503\,
            I => \N__44476\
        );

    \I__9957\ : Span4Mux_v
    port map (
            O => \N__44500\,
            I => \N__44473\
        );

    \I__9956\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44456\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44498\,
            I => \N__44456\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44497\,
            I => \N__44456\
        );

    \I__9953\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44456\
        );

    \I__9952\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44456\
        );

    \I__9951\ : InMux
    port map (
            O => \N__44494\,
            I => \N__44456\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44456\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44456\
        );

    \I__9948\ : CascadeMux
    port map (
            O => \N__44491\,
            I => \N__44446\
        );

    \I__9947\ : Span4Mux_h
    port map (
            O => \N__44488\,
            I => \N__44439\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__44485\,
            I => \N__44439\
        );

    \I__9945\ : Span4Mux_v
    port map (
            O => \N__44482\,
            I => \N__44436\
        );

    \I__9944\ : LocalMux
    port map (
            O => \N__44479\,
            I => \N__44433\
        );

    \I__9943\ : LocalMux
    port map (
            O => \N__44476\,
            I => \N__44430\
        );

    \I__9942\ : Span4Mux_h
    port map (
            O => \N__44473\,
            I => \N__44425\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__44456\,
            I => \N__44425\
        );

    \I__9940\ : InMux
    port map (
            O => \N__44455\,
            I => \N__44410\
        );

    \I__9939\ : InMux
    port map (
            O => \N__44454\,
            I => \N__44410\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44453\,
            I => \N__44410\
        );

    \I__9937\ : InMux
    port map (
            O => \N__44452\,
            I => \N__44410\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44451\,
            I => \N__44410\
        );

    \I__9935\ : InMux
    port map (
            O => \N__44450\,
            I => \N__44410\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44449\,
            I => \N__44410\
        );

    \I__9933\ : InMux
    port map (
            O => \N__44446\,
            I => \N__44401\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44445\,
            I => \N__44401\
        );

    \I__9931\ : InMux
    port map (
            O => \N__44444\,
            I => \N__44401\
        );

    \I__9930\ : Span4Mux_v
    port map (
            O => \N__44439\,
            I => \N__44394\
        );

    \I__9929\ : Span4Mux_h
    port map (
            O => \N__44436\,
            I => \N__44394\
        );

    \I__9928\ : Span4Mux_h
    port map (
            O => \N__44433\,
            I => \N__44394\
        );

    \I__9927\ : Span4Mux_h
    port map (
            O => \N__44430\,
            I => \N__44389\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__44425\,
            I => \N__44389\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44410\,
            I => \N__44385\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44380\
        );

    \I__9923\ : InMux
    port map (
            O => \N__44408\,
            I => \N__44380\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__44401\,
            I => \N__44377\
        );

    \I__9921\ : Span4Mux_h
    port map (
            O => \N__44394\,
            I => \N__44373\
        );

    \I__9920\ : Span4Mux_h
    port map (
            O => \N__44389\,
            I => \N__44370\
        );

    \I__9919\ : InMux
    port map (
            O => \N__44388\,
            I => \N__44367\
        );

    \I__9918\ : Span4Mux_h
    port map (
            O => \N__44385\,
            I => \N__44360\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__44380\,
            I => \N__44360\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__44377\,
            I => \N__44360\
        );

    \I__9915\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44357\
        );

    \I__9914\ : Span4Mux_h
    port map (
            O => \N__44373\,
            I => \N__44354\
        );

    \I__9913\ : Odrv4
    port map (
            O => \N__44370\,
            I => dds_state_1
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__44367\,
            I => dds_state_1
        );

    \I__9911\ : Odrv4
    port map (
            O => \N__44360\,
            I => dds_state_1
        );

    \I__9910\ : LocalMux
    port map (
            O => \N__44357\,
            I => dds_state_1
        );

    \I__9909\ : Odrv4
    port map (
            O => \N__44354\,
            I => dds_state_1
        );

    \I__9908\ : InMux
    port map (
            O => \N__44343\,
            I => \N__44340\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__44340\,
            I => \comm_spi.n14813\
        );

    \I__9906\ : InMux
    port map (
            O => \N__44337\,
            I => \N__44334\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__44334\,
            I => \comm_spi.n14812\
        );

    \I__9904\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44327\
        );

    \I__9903\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44324\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__44327\,
            I => \N__44320\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__44324\,
            I => \N__44317\
        );

    \I__9900\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44314\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__44320\,
            I => \N__44304\
        );

    \I__9898\ : Span4Mux_h
    port map (
            O => \N__44317\,
            I => \N__44304\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44304\
        );

    \I__9896\ : InMux
    port map (
            O => \N__44313\,
            I => \N__44301\
        );

    \I__9895\ : InMux
    port map (
            O => \N__44312\,
            I => \N__44298\
        );

    \I__9894\ : InMux
    port map (
            O => \N__44311\,
            I => \N__44295\
        );

    \I__9893\ : Sp12to4
    port map (
            O => \N__44304\,
            I => \N__44288\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__44301\,
            I => \N__44288\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__44298\,
            I => \N__44288\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__44295\,
            I => \comm_spi.n14811\
        );

    \I__9889\ : Odrv12
    port map (
            O => \N__44288\,
            I => \comm_spi.n14811\
        );

    \I__9888\ : IoInMux
    port map (
            O => \N__44283\,
            I => \N__44280\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__44280\,
            I => \N__44277\
        );

    \I__9886\ : IoSpan4Mux
    port map (
            O => \N__44277\,
            I => \N__44274\
        );

    \I__9885\ : IoSpan4Mux
    port map (
            O => \N__44274\,
            I => \N__44271\
        );

    \I__9884\ : Span4Mux_s3_h
    port map (
            O => \N__44271\,
            I => \N__44268\
        );

    \I__9883\ : Span4Mux_h
    port map (
            O => \N__44268\,
            I => \N__44265\
        );

    \I__9882\ : Odrv4
    port map (
            O => \N__44265\,
            I => \ICE_SPI_MISO\
        );

    \I__9881\ : InMux
    port map (
            O => \N__44262\,
            I => \N__44259\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__44259\,
            I => \ADC_VDC.n11895\
        );

    \I__9879\ : InMux
    port map (
            O => \N__44256\,
            I => \N__44253\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__44253\,
            I => \comm_spi.n23086\
        );

    \I__9877\ : CascadeMux
    port map (
            O => \N__44250\,
            I => \comm_spi.n23086_cascade_\
        );

    \I__9876\ : InMux
    port map (
            O => \N__44247\,
            I => \N__44244\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__44244\,
            I => \comm_spi.n14804\
        );

    \I__9874\ : InMux
    port map (
            O => \N__44241\,
            I => \N__44238\
        );

    \I__9873\ : LocalMux
    port map (
            O => \N__44238\,
            I => n80
        );

    \I__9872\ : CascadeMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__9871\ : InMux
    port map (
            O => \N__44232\,
            I => \N__44229\
        );

    \I__9870\ : LocalMux
    port map (
            O => \N__44229\,
            I => \N__44226\
        );

    \I__9869\ : Span4Mux_h
    port map (
            O => \N__44226\,
            I => \N__44223\
        );

    \I__9868\ : Span4Mux_h
    port map (
            O => \N__44223\,
            I => \N__44220\
        );

    \I__9867\ : Odrv4
    port map (
            O => \N__44220\,
            I => n5
        );

    \I__9866\ : InMux
    port map (
            O => \N__44217\,
            I => \N__44214\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__44214\,
            I => \N__44210\
        );

    \I__9864\ : InMux
    port map (
            O => \N__44213\,
            I => \N__44207\
        );

    \I__9863\ : Span12Mux_v
    port map (
            O => \N__44210\,
            I => \N__44204\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__44207\,
            I => data_idxvec_1
        );

    \I__9861\ : Odrv12
    port map (
            O => \N__44204\,
            I => data_idxvec_1
        );

    \I__9860\ : InMux
    port map (
            O => \N__44199\,
            I => \N__44196\
        );

    \I__9859\ : LocalMux
    port map (
            O => \N__44196\,
            I => \N__44191\
        );

    \I__9858\ : InMux
    port map (
            O => \N__44195\,
            I => \N__44188\
        );

    \I__9857\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44185\
        );

    \I__9856\ : Span4Mux_h
    port map (
            O => \N__44191\,
            I => \N__44182\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__44188\,
            I => data_cntvec_1
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__44185\,
            I => data_cntvec_1
        );

    \I__9853\ : Odrv4
    port map (
            O => \N__44182\,
            I => data_cntvec_1
        );

    \I__9852\ : CascadeMux
    port map (
            O => \N__44175\,
            I => \n26_adj_1653_cascade_\
        );

    \I__9851\ : InMux
    port map (
            O => \N__44172\,
            I => \N__44169\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__9849\ : Span4Mux_v
    port map (
            O => \N__44166\,
            I => \N__44161\
        );

    \I__9848\ : InMux
    port map (
            O => \N__44165\,
            I => \N__44156\
        );

    \I__9847\ : InMux
    port map (
            O => \N__44164\,
            I => \N__44156\
        );

    \I__9846\ : Odrv4
    port map (
            O => \N__44161\,
            I => \acadc_skipCount_1\
        );

    \I__9845\ : LocalMux
    port map (
            O => \N__44156\,
            I => \acadc_skipCount_1\
        );

    \I__9844\ : CascadeMux
    port map (
            O => \N__44151\,
            I => \n22497_cascade_\
        );

    \I__9843\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44145\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__44145\,
            I => \N__44142\
        );

    \I__9841\ : Span4Mux_h
    port map (
            O => \N__44142\,
            I => \N__44137\
        );

    \I__9840\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44132\
        );

    \I__9839\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44132\
        );

    \I__9838\ : Odrv4
    port map (
            O => \N__44137\,
            I => req_data_cnt_1
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__44132\,
            I => req_data_cnt_1
        );

    \I__9836\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44124\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__44124\,
            I => n22434
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__44121\,
            I => \n22500_cascade_\
        );

    \I__9833\ : CascadeMux
    port map (
            O => \N__44118\,
            I => \n30_adj_1654_cascade_\
        );

    \I__9832\ : CascadeMux
    port map (
            O => \N__44115\,
            I => \N__44111\
        );

    \I__9831\ : InMux
    port map (
            O => \N__44114\,
            I => \N__44108\
        );

    \I__9830\ : InMux
    port map (
            O => \N__44111\,
            I => \N__44105\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__44108\,
            I => \N__44102\
        );

    \I__9828\ : LocalMux
    port map (
            O => \N__44105\,
            I => \N__44099\
        );

    \I__9827\ : Span4Mux_h
    port map (
            O => \N__44102\,
            I => \N__44096\
        );

    \I__9826\ : Span4Mux_v
    port map (
            O => \N__44099\,
            I => \N__44093\
        );

    \I__9825\ : Span4Mux_v
    port map (
            O => \N__44096\,
            I => \N__44090\
        );

    \I__9824\ : Span4Mux_h
    port map (
            O => \N__44093\,
            I => \N__44087\
        );

    \I__9823\ : Odrv4
    port map (
            O => \N__44090\,
            I => n28
        );

    \I__9822\ : Odrv4
    port map (
            O => \N__44087\,
            I => n28
        );

    \I__9821\ : CascadeMux
    port map (
            O => \N__44082\,
            I => \N__44079\
        );

    \I__9820\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44075\
        );

    \I__9819\ : CascadeMux
    port map (
            O => \N__44078\,
            I => \N__44072\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__44075\,
            I => \N__44068\
        );

    \I__9817\ : InMux
    port map (
            O => \N__44072\,
            I => \N__44065\
        );

    \I__9816\ : InMux
    port map (
            O => \N__44071\,
            I => \N__44062\
        );

    \I__9815\ : Span4Mux_h
    port map (
            O => \N__44068\,
            I => \N__44054\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__44065\,
            I => \N__44054\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__44062\,
            I => \N__44051\
        );

    \I__9812\ : InMux
    port map (
            O => \N__44061\,
            I => \N__44048\
        );

    \I__9811\ : InMux
    port map (
            O => \N__44060\,
            I => \N__44043\
        );

    \I__9810\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44043\
        );

    \I__9809\ : Span4Mux_v
    port map (
            O => \N__44054\,
            I => \N__44040\
        );

    \I__9808\ : Span4Mux_h
    port map (
            O => \N__44051\,
            I => \N__44037\
        );

    \I__9807\ : LocalMux
    port map (
            O => \N__44048\,
            I => \N__44032\
        );

    \I__9806\ : LocalMux
    port map (
            O => \N__44043\,
            I => \N__44032\
        );

    \I__9805\ : Span4Mux_h
    port map (
            O => \N__44040\,
            I => \N__44029\
        );

    \I__9804\ : Span4Mux_v
    port map (
            O => \N__44037\,
            I => \N__44026\
        );

    \I__9803\ : Span12Mux_v
    port map (
            O => \N__44032\,
            I => \N__44023\
        );

    \I__9802\ : Odrv4
    port map (
            O => \N__44029\,
            I => comm_buf_1_7
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__44026\,
            I => comm_buf_1_7
        );

    \I__9800\ : Odrv12
    port map (
            O => \N__44023\,
            I => comm_buf_1_7
        );

    \I__9799\ : SRMux
    port map (
            O => \N__44016\,
            I => \N__44010\
        );

    \I__9798\ : SRMux
    port map (
            O => \N__44015\,
            I => \N__44006\
        );

    \I__9797\ : SRMux
    port map (
            O => \N__44014\,
            I => \N__44003\
        );

    \I__9796\ : SRMux
    port map (
            O => \N__44013\,
            I => \N__43998\
        );

    \I__9795\ : LocalMux
    port map (
            O => \N__44010\,
            I => \N__43995\
        );

    \I__9794\ : SRMux
    port map (
            O => \N__44009\,
            I => \N__43992\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__44006\,
            I => \N__43989\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__44003\,
            I => \N__43986\
        );

    \I__9791\ : SRMux
    port map (
            O => \N__44002\,
            I => \N__43983\
        );

    \I__9790\ : SRMux
    port map (
            O => \N__44001\,
            I => \N__43980\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43998\,
            I => \N__43973\
        );

    \I__9788\ : Span4Mux_h
    port map (
            O => \N__43995\,
            I => \N__43973\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43992\,
            I => \N__43973\
        );

    \I__9786\ : Span4Mux_h
    port map (
            O => \N__43989\,
            I => \N__43966\
        );

    \I__9785\ : Span4Mux_v
    port map (
            O => \N__43986\,
            I => \N__43966\
        );

    \I__9784\ : LocalMux
    port map (
            O => \N__43983\,
            I => \N__43966\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43980\,
            I => \N__43963\
        );

    \I__9782\ : Span4Mux_v
    port map (
            O => \N__43973\,
            I => \N__43957\
        );

    \I__9781\ : Span4Mux_h
    port map (
            O => \N__43966\,
            I => \N__43957\
        );

    \I__9780\ : Span4Mux_h
    port map (
            O => \N__43963\,
            I => \N__43954\
        );

    \I__9779\ : SRMux
    port map (
            O => \N__43962\,
            I => \N__43951\
        );

    \I__9778\ : Odrv4
    port map (
            O => \N__43957\,
            I => n14965
        );

    \I__9777\ : Odrv4
    port map (
            O => \N__43954\,
            I => n14965
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43951\,
            I => n14965
        );

    \I__9775\ : CascadeMux
    port map (
            O => \N__43944\,
            I => \N__43940\
        );

    \I__9774\ : CascadeMux
    port map (
            O => \N__43943\,
            I => \N__43937\
        );

    \I__9773\ : InMux
    port map (
            O => \N__43940\,
            I => \N__43933\
        );

    \I__9772\ : InMux
    port map (
            O => \N__43937\,
            I => \N__43930\
        );

    \I__9771\ : CascadeMux
    port map (
            O => \N__43936\,
            I => \N__43927\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__43933\,
            I => \N__43921\
        );

    \I__9769\ : LocalMux
    port map (
            O => \N__43930\,
            I => \N__43921\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43927\,
            I => \N__43916\
        );

    \I__9767\ : InMux
    port map (
            O => \N__43926\,
            I => \N__43916\
        );

    \I__9766\ : Odrv4
    port map (
            O => \N__43921\,
            I => trig_dds0
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__43916\,
            I => trig_dds0
        );

    \I__9764\ : CEMux
    port map (
            O => \N__43911\,
            I => \N__43907\
        );

    \I__9763\ : CEMux
    port map (
            O => \N__43910\,
            I => \N__43904\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43907\,
            I => \N__43900\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__43904\,
            I => \N__43897\
        );

    \I__9760\ : CEMux
    port map (
            O => \N__43903\,
            I => \N__43894\
        );

    \I__9759\ : Span4Mux_v
    port map (
            O => \N__43900\,
            I => \N__43891\
        );

    \I__9758\ : Span4Mux_h
    port map (
            O => \N__43897\,
            I => \N__43888\
        );

    \I__9757\ : LocalMux
    port map (
            O => \N__43894\,
            I => \N__43885\
        );

    \I__9756\ : Span4Mux_h
    port map (
            O => \N__43891\,
            I => \N__43882\
        );

    \I__9755\ : Span4Mux_h
    port map (
            O => \N__43888\,
            I => \N__43879\
        );

    \I__9754\ : Span12Mux_h
    port map (
            O => \N__43885\,
            I => \N__43876\
        );

    \I__9753\ : Odrv4
    port map (
            O => \N__43882\,
            I => \SIG_DDS.n12895\
        );

    \I__9752\ : Odrv4
    port map (
            O => \N__43879\,
            I => \SIG_DDS.n12895\
        );

    \I__9751\ : Odrv12
    port map (
            O => \N__43876\,
            I => \SIG_DDS.n12895\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43869\,
            I => \N__43866\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43862\
        );

    \I__9748\ : CascadeMux
    port map (
            O => \N__43865\,
            I => \N__43859\
        );

    \I__9747\ : Span4Mux_v
    port map (
            O => \N__43862\,
            I => \N__43856\
        );

    \I__9746\ : InMux
    port map (
            O => \N__43859\,
            I => \N__43853\
        );

    \I__9745\ : Span4Mux_h
    port map (
            O => \N__43856\,
            I => \N__43850\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__43853\,
            I => data_idxvec_0
        );

    \I__9743\ : Odrv4
    port map (
            O => \N__43850\,
            I => data_idxvec_0
        );

    \I__9742\ : InMux
    port map (
            O => \N__43845\,
            I => \N__43841\
        );

    \I__9741\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43837\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__43841\,
            I => \N__43834\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43840\,
            I => \N__43831\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__43837\,
            I => \N__43828\
        );

    \I__9737\ : Span4Mux_h
    port map (
            O => \N__43834\,
            I => \N__43825\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43831\,
            I => data_cntvec_0
        );

    \I__9735\ : Odrv12
    port map (
            O => \N__43828\,
            I => data_cntvec_0
        );

    \I__9734\ : Odrv4
    port map (
            O => \N__43825\,
            I => data_cntvec_0
        );

    \I__9733\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43815\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__43815\,
            I => \N__43812\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__43812\,
            I => \N__43809\
        );

    \I__9730\ : Span4Mux_h
    port map (
            O => \N__43809\,
            I => \N__43806\
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__43806\,
            I => buf_data_iac_8
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__43803\,
            I => \n26_cascade_\
        );

    \I__9727\ : CascadeMux
    port map (
            O => \N__43800\,
            I => \n21261_cascade_\
        );

    \I__9726\ : CascadeMux
    port map (
            O => \N__43797\,
            I => \n22563_cascade_\
        );

    \I__9725\ : InMux
    port map (
            O => \N__43794\,
            I => \N__43791\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__43791\,
            I => \N__43788\
        );

    \I__9723\ : Odrv4
    port map (
            O => \N__43788\,
            I => n21257
        );

    \I__9722\ : CascadeMux
    port map (
            O => \N__43785\,
            I => \n22566_cascade_\
        );

    \I__9721\ : InMux
    port map (
            O => \N__43782\,
            I => \N__43779\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43779\,
            I => \N__43776\
        );

    \I__9719\ : Span4Mux_v
    port map (
            O => \N__43776\,
            I => \N__43773\
        );

    \I__9718\ : Sp12to4
    port map (
            O => \N__43773\,
            I => \N__43770\
        );

    \I__9717\ : Span12Mux_h
    port map (
            O => \N__43770\,
            I => \N__43766\
        );

    \I__9716\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43763\
        );

    \I__9715\ : Odrv12
    port map (
            O => \N__43766\,
            I => buf_adcdata_vdc_8
        );

    \I__9714\ : LocalMux
    port map (
            O => \N__43763\,
            I => buf_adcdata_vdc_8
        );

    \I__9713\ : InMux
    port map (
            O => \N__43758\,
            I => \N__43754\
        );

    \I__9712\ : CascadeMux
    port map (
            O => \N__43757\,
            I => \N__43751\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43754\,
            I => \N__43748\
        );

    \I__9710\ : InMux
    port map (
            O => \N__43751\,
            I => \N__43745\
        );

    \I__9709\ : Span4Mux_v
    port map (
            O => \N__43748\,
            I => \N__43742\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43745\,
            I => \N__43738\
        );

    \I__9707\ : Span4Mux_h
    port map (
            O => \N__43742\,
            I => \N__43735\
        );

    \I__9706\ : CascadeMux
    port map (
            O => \N__43741\,
            I => \N__43732\
        );

    \I__9705\ : Span4Mux_v
    port map (
            O => \N__43738\,
            I => \N__43729\
        );

    \I__9704\ : Span4Mux_h
    port map (
            O => \N__43735\,
            I => \N__43726\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43732\,
            I => \N__43723\
        );

    \I__9702\ : Span4Mux_h
    port map (
            O => \N__43729\,
            I => \N__43720\
        );

    \I__9701\ : Span4Mux_h
    port map (
            O => \N__43726\,
            I => \N__43717\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__43723\,
            I => buf_adcdata_vac_8
        );

    \I__9699\ : Odrv4
    port map (
            O => \N__43720\,
            I => buf_adcdata_vac_8
        );

    \I__9698\ : Odrv4
    port map (
            O => \N__43717\,
            I => buf_adcdata_vac_8
        );

    \I__9697\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43707\
        );

    \I__9696\ : LocalMux
    port map (
            O => \N__43707\,
            I => \N__43704\
        );

    \I__9695\ : Span4Mux_h
    port map (
            O => \N__43704\,
            I => \N__43701\
        );

    \I__9694\ : Span4Mux_v
    port map (
            O => \N__43701\,
            I => \N__43698\
        );

    \I__9693\ : Span4Mux_h
    port map (
            O => \N__43698\,
            I => \N__43694\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43697\,
            I => \N__43691\
        );

    \I__9691\ : Odrv4
    port map (
            O => \N__43694\,
            I => \buf_readRTD_0\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__43691\,
            I => \buf_readRTD_0\
        );

    \I__9689\ : CascadeMux
    port map (
            O => \N__43686\,
            I => \n19_cascade_\
        );

    \I__9688\ : InMux
    port map (
            O => \N__43683\,
            I => \N__43680\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__43680\,
            I => n21258
        );

    \I__9686\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43673\
        );

    \I__9685\ : InMux
    port map (
            O => \N__43676\,
            I => \N__43669\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__43673\,
            I => \N__43666\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43663\
        );

    \I__9682\ : LocalMux
    port map (
            O => \N__43669\,
            I => \acadc_skipCount_0\
        );

    \I__9681\ : Odrv12
    port map (
            O => \N__43666\,
            I => \acadc_skipCount_0\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__43663\,
            I => \acadc_skipCount_0\
        );

    \I__9679\ : InMux
    port map (
            O => \N__43656\,
            I => \N__43653\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__43653\,
            I => \N__43650\
        );

    \I__9677\ : Span4Mux_h
    port map (
            O => \N__43650\,
            I => \N__43645\
        );

    \I__9676\ : CascadeMux
    port map (
            O => \N__43649\,
            I => \N__43642\
        );

    \I__9675\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43639\
        );

    \I__9674\ : Span4Mux_h
    port map (
            O => \N__43645\,
            I => \N__43636\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43642\,
            I => \N__43633\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__43639\,
            I => req_data_cnt_0
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__43636\,
            I => req_data_cnt_0
        );

    \I__9670\ : LocalMux
    port map (
            O => \N__43633\,
            I => req_data_cnt_0
        );

    \I__9669\ : InMux
    port map (
            O => \N__43626\,
            I => \N__43623\
        );

    \I__9668\ : LocalMux
    port map (
            O => \N__43623\,
            I => n21260
        );

    \I__9667\ : InMux
    port map (
            O => \N__43620\,
            I => \N__43617\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__43617\,
            I => \N__43614\
        );

    \I__9665\ : Span4Mux_h
    port map (
            O => \N__43614\,
            I => \N__43610\
        );

    \I__9664\ : InMux
    port map (
            O => \N__43613\,
            I => \N__43607\
        );

    \I__9663\ : Span4Mux_v
    port map (
            O => \N__43610\,
            I => \N__43602\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__43607\,
            I => \N__43602\
        );

    \I__9661\ : Span4Mux_h
    port map (
            O => \N__43602\,
            I => \N__43598\
        );

    \I__9660\ : InMux
    port map (
            O => \N__43601\,
            I => \N__43595\
        );

    \I__9659\ : Span4Mux_h
    port map (
            O => \N__43598\,
            I => \N__43592\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__43595\,
            I => buf_adcdata_iac_9
        );

    \I__9657\ : Odrv4
    port map (
            O => \N__43592\,
            I => buf_adcdata_iac_9
        );

    \I__9656\ : CascadeMux
    port map (
            O => \N__43587\,
            I => \N__43584\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43581\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__43581\,
            I => \N__43578\
        );

    \I__9653\ : Odrv12
    port map (
            O => \N__43578\,
            I => n16_adj_1651
        );

    \I__9652\ : InMux
    port map (
            O => \N__43575\,
            I => \N__43572\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__43572\,
            I => \N__43569\
        );

    \I__9650\ : Span4Mux_v
    port map (
            O => \N__43569\,
            I => \N__43566\
        );

    \I__9649\ : Span4Mux_h
    port map (
            O => \N__43566\,
            I => \N__43563\
        );

    \I__9648\ : Odrv4
    port map (
            O => \N__43563\,
            I => n22431
        );

    \I__9647\ : CascadeMux
    port map (
            O => \N__43560\,
            I => \N__43556\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43553\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43550\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__43553\,
            I => \N__43547\
        );

    \I__9643\ : LocalMux
    port map (
            O => \N__43550\,
            I => comm_buf_6_7
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__43547\,
            I => comm_buf_6_7
        );

    \I__9641\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43539\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__43539\,
            I => \N__43535\
        );

    \I__9639\ : InMux
    port map (
            O => \N__43538\,
            I => \N__43531\
        );

    \I__9638\ : Span4Mux_h
    port map (
            O => \N__43535\,
            I => \N__43528\
        );

    \I__9637\ : InMux
    port map (
            O => \N__43534\,
            I => \N__43525\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__43531\,
            I => \acadc_skipCount_6\
        );

    \I__9635\ : Odrv4
    port map (
            O => \N__43528\,
            I => \acadc_skipCount_6\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__43525\,
            I => \acadc_skipCount_6\
        );

    \I__9633\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43514\
        );

    \I__9632\ : InMux
    port map (
            O => \N__43517\,
            I => \N__43510\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__43514\,
            I => \N__43507\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43504\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__43510\,
            I => req_data_cnt_6
        );

    \I__9628\ : Odrv12
    port map (
            O => \N__43507\,
            I => req_data_cnt_6
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43504\,
            I => req_data_cnt_6
        );

    \I__9626\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43494\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__43494\,
            I => \N__43491\
        );

    \I__9624\ : Odrv12
    port map (
            O => \N__43491\,
            I => n19_adj_1625
        );

    \I__9623\ : CascadeMux
    port map (
            O => \N__43488\,
            I => \N__43485\
        );

    \I__9622\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43482\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__43482\,
            I => \N__43479\
        );

    \I__9620\ : Span4Mux_v
    port map (
            O => \N__43479\,
            I => \N__43476\
        );

    \I__9619\ : Span4Mux_h
    port map (
            O => \N__43476\,
            I => \N__43473\
        );

    \I__9618\ : Sp12to4
    port map (
            O => \N__43473\,
            I => \N__43469\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43466\
        );

    \I__9616\ : Odrv12
    port map (
            O => \N__43469\,
            I => \buf_readRTD_6\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__43466\,
            I => \buf_readRTD_6\
        );

    \I__9614\ : InMux
    port map (
            O => \N__43461\,
            I => \N__43458\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__43458\,
            I => \N__43454\
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__43457\,
            I => \N__43451\
        );

    \I__9611\ : Span4Mux_h
    port map (
            O => \N__43454\,
            I => \N__43448\
        );

    \I__9610\ : InMux
    port map (
            O => \N__43451\,
            I => \N__43445\
        );

    \I__9609\ : Span4Mux_h
    port map (
            O => \N__43448\,
            I => \N__43442\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__43445\,
            I => data_idxvec_6
        );

    \I__9607\ : Odrv4
    port map (
            O => \N__43442\,
            I => data_idxvec_6
        );

    \I__9606\ : InMux
    port map (
            O => \N__43437\,
            I => \N__43433\
        );

    \I__9605\ : InMux
    port map (
            O => \N__43436\,
            I => \N__43429\
        );

    \I__9604\ : LocalMux
    port map (
            O => \N__43433\,
            I => \N__43426\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43432\,
            I => \N__43423\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__43429\,
            I => \N__43416\
        );

    \I__9601\ : Span4Mux_h
    port map (
            O => \N__43426\,
            I => \N__43416\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__43423\,
            I => \N__43416\
        );

    \I__9599\ : Odrv4
    port map (
            O => \N__43416\,
            I => data_cntvec_6
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__43413\,
            I => \n26_adj_1626_cascade_\
        );

    \I__9597\ : InMux
    port map (
            O => \N__43410\,
            I => \N__43407\
        );

    \I__9596\ : LocalMux
    port map (
            O => \N__43407\,
            I => n22515
        );

    \I__9595\ : InMux
    port map (
            O => \N__43404\,
            I => \N__43401\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__43401\,
            I => \N__43398\
        );

    \I__9593\ : Span4Mux_h
    port map (
            O => \N__43398\,
            I => \N__43395\
        );

    \I__9592\ : Odrv4
    port map (
            O => \N__43395\,
            I => n16_adj_1624
        );

    \I__9591\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43389\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__43389\,
            I => \N__43385\
        );

    \I__9589\ : CascadeMux
    port map (
            O => \N__43388\,
            I => \N__43382\
        );

    \I__9588\ : Span4Mux_v
    port map (
            O => \N__43385\,
            I => \N__43379\
        );

    \I__9587\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43375\
        );

    \I__9586\ : Sp12to4
    port map (
            O => \N__43379\,
            I => \N__43372\
        );

    \I__9585\ : InMux
    port map (
            O => \N__43378\,
            I => \N__43369\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__43375\,
            I => \N__43364\
        );

    \I__9583\ : Span12Mux_s10_h
    port map (
            O => \N__43372\,
            I => \N__43364\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__43369\,
            I => buf_adcdata_iac_14
        );

    \I__9581\ : Odrv12
    port map (
            O => \N__43364\,
            I => buf_adcdata_iac_14
        );

    \I__9580\ : InMux
    port map (
            O => \N__43359\,
            I => \N__43356\
        );

    \I__9579\ : LocalMux
    port map (
            O => \N__43356\,
            I => n22527
        );

    \I__9578\ : CascadeMux
    port map (
            O => \N__43353\,
            I => \n22530_cascade_\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43347\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__43347\,
            I => n22518
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__43344\,
            I => \n30_adj_1627_cascade_\
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__43341\,
            I => \n30_adj_1695_cascade_\
        );

    \I__9573\ : CEMux
    port map (
            O => \N__43338\,
            I => \N__43333\
        );

    \I__9572\ : CEMux
    port map (
            O => \N__43337\,
            I => \N__43330\
        );

    \I__9571\ : CEMux
    port map (
            O => \N__43336\,
            I => \N__43327\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__43333\,
            I => \N__43321\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__43330\,
            I => \N__43318\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__43327\,
            I => \N__43315\
        );

    \I__9567\ : CEMux
    port map (
            O => \N__43326\,
            I => \N__43312\
        );

    \I__9566\ : CEMux
    port map (
            O => \N__43325\,
            I => \N__43309\
        );

    \I__9565\ : CEMux
    port map (
            O => \N__43324\,
            I => \N__43306\
        );

    \I__9564\ : Span4Mux_h
    port map (
            O => \N__43321\,
            I => \N__43302\
        );

    \I__9563\ : Span4Mux_v
    port map (
            O => \N__43318\,
            I => \N__43295\
        );

    \I__9562\ : Span4Mux_h
    port map (
            O => \N__43315\,
            I => \N__43295\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43312\,
            I => \N__43295\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__43309\,
            I => \N__43292\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__43306\,
            I => \N__43289\
        );

    \I__9558\ : InMux
    port map (
            O => \N__43305\,
            I => \N__43286\
        );

    \I__9557\ : Odrv4
    port map (
            O => \N__43302\,
            I => n12184
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__43295\,
            I => n12184
        );

    \I__9555\ : Odrv12
    port map (
            O => \N__43292\,
            I => n12184
        );

    \I__9554\ : Odrv4
    port map (
            O => \N__43289\,
            I => n12184
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__43286\,
            I => n12184
        );

    \I__9552\ : SRMux
    port map (
            O => \N__43275\,
            I => \N__43271\
        );

    \I__9551\ : SRMux
    port map (
            O => \N__43274\,
            I => \N__43268\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__43271\,
            I => \N__43265\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__43268\,
            I => \N__43260\
        );

    \I__9548\ : Span4Mux_h
    port map (
            O => \N__43265\,
            I => \N__43257\
        );

    \I__9547\ : SRMux
    port map (
            O => \N__43264\,
            I => \N__43254\
        );

    \I__9546\ : SRMux
    port map (
            O => \N__43263\,
            I => \N__43251\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__43260\,
            I => \N__43242\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__43257\,
            I => \N__43242\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__43254\,
            I => \N__43242\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__43251\,
            I => \N__43239\
        );

    \I__9541\ : SRMux
    port map (
            O => \N__43250\,
            I => \N__43236\
        );

    \I__9540\ : SRMux
    port map (
            O => \N__43249\,
            I => \N__43233\
        );

    \I__9539\ : Span4Mux_v
    port map (
            O => \N__43242\,
            I => \N__43230\
        );

    \I__9538\ : Sp12to4
    port map (
            O => \N__43239\,
            I => \N__43225\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__43236\,
            I => \N__43225\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__43233\,
            I => \N__43222\
        );

    \I__9535\ : Odrv4
    port map (
            O => \N__43230\,
            I => n14958
        );

    \I__9534\ : Odrv12
    port map (
            O => \N__43225\,
            I => n14958
        );

    \I__9533\ : Odrv12
    port map (
            O => \N__43222\,
            I => n14958
        );

    \I__9532\ : InMux
    port map (
            O => \N__43215\,
            I => \N__43212\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__43212\,
            I => \N__43209\
        );

    \I__9530\ : Odrv12
    port map (
            O => \N__43209\,
            I => n22539
        );

    \I__9529\ : InMux
    port map (
            O => \N__43206\,
            I => \N__43203\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__43203\,
            I => \N__43200\
        );

    \I__9527\ : Span4Mux_v
    port map (
            O => \N__43200\,
            I => \N__43195\
        );

    \I__9526\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43191\
        );

    \I__9525\ : InMux
    port map (
            O => \N__43198\,
            I => \N__43188\
        );

    \I__9524\ : Span4Mux_h
    port map (
            O => \N__43195\,
            I => \N__43185\
        );

    \I__9523\ : InMux
    port map (
            O => \N__43194\,
            I => \N__43182\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__43191\,
            I => \N__43179\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__43188\,
            I => \N__43176\
        );

    \I__9520\ : Span4Mux_h
    port map (
            O => \N__43185\,
            I => \N__43173\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__43182\,
            I => \N__43170\
        );

    \I__9518\ : Span4Mux_v
    port map (
            O => \N__43179\,
            I => \N__43165\
        );

    \I__9517\ : Span4Mux_v
    port map (
            O => \N__43176\,
            I => \N__43165\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__43173\,
            I => \N__43162\
        );

    \I__9515\ : Span4Mux_v
    port map (
            O => \N__43170\,
            I => \N__43157\
        );

    \I__9514\ : Span4Mux_h
    port map (
            O => \N__43165\,
            I => \N__43157\
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__43162\,
            I => n14_adj_1541
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__43157\,
            I => n14_adj_1541
        );

    \I__9511\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43149\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__43149\,
            I => \N__43146\
        );

    \I__9509\ : Span4Mux_h
    port map (
            O => \N__43146\,
            I => \N__43143\
        );

    \I__9508\ : Span4Mux_v
    port map (
            O => \N__43143\,
            I => \N__43140\
        );

    \I__9507\ : Odrv4
    port map (
            O => \N__43140\,
            I => buf_data_iac_0
        );

    \I__9506\ : InMux
    port map (
            O => \N__43137\,
            I => \N__43134\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__43134\,
            I => \N__43131\
        );

    \I__9504\ : Span12Mux_v
    port map (
            O => \N__43131\,
            I => \N__43128\
        );

    \I__9503\ : Odrv12
    port map (
            O => \N__43128\,
            I => n22_adj_1532
        );

    \I__9502\ : CascadeMux
    port map (
            O => \N__43125\,
            I => \N__43122\
        );

    \I__9501\ : InMux
    port map (
            O => \N__43122\,
            I => \N__43119\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__43119\,
            I => \N__43116\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__43116\,
            I => n21586
        );

    \I__9498\ : CascadeMux
    port map (
            O => \N__43113\,
            I => \n21474_cascade_\
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__43110\,
            I => \n12_adj_1596_cascade_\
        );

    \I__9496\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43103\
        );

    \I__9495\ : CascadeMux
    port map (
            O => \N__43106\,
            I => \N__43100\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__43103\,
            I => \N__43097\
        );

    \I__9493\ : InMux
    port map (
            O => \N__43100\,
            I => \N__43094\
        );

    \I__9492\ : Span12Mux_v
    port map (
            O => \N__43097\,
            I => \N__43091\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__43094\,
            I => data_idxvec_9
        );

    \I__9490\ : Odrv12
    port map (
            O => \N__43091\,
            I => data_idxvec_9
        );

    \I__9489\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43082\
        );

    \I__9488\ : InMux
    port map (
            O => \N__43085\,
            I => \N__43079\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__43082\,
            I => \N__43075\
        );

    \I__9486\ : LocalMux
    port map (
            O => \N__43079\,
            I => \N__43072\
        );

    \I__9485\ : InMux
    port map (
            O => \N__43078\,
            I => \N__43069\
        );

    \I__9484\ : Span4Mux_v
    port map (
            O => \N__43075\,
            I => \N__43064\
        );

    \I__9483\ : Span4Mux_h
    port map (
            O => \N__43072\,
            I => \N__43064\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__43069\,
            I => data_cntvec_9
        );

    \I__9481\ : Odrv4
    port map (
            O => \N__43064\,
            I => data_cntvec_9
        );

    \I__9480\ : InMux
    port map (
            O => \N__43059\,
            I => \N__43056\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__43056\,
            I => \N__43053\
        );

    \I__9478\ : Odrv12
    port map (
            O => \N__43053\,
            I => buf_data_iac_17
        );

    \I__9477\ : CascadeMux
    port map (
            O => \N__43050\,
            I => \n26_adj_1694_cascade_\
        );

    \I__9476\ : InMux
    port map (
            O => \N__43047\,
            I => \N__43044\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__43044\,
            I => \N__43038\
        );

    \I__9474\ : InMux
    port map (
            O => \N__43043\,
            I => \N__43035\
        );

    \I__9473\ : InMux
    port map (
            O => \N__43042\,
            I => \N__43032\
        );

    \I__9472\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43029\
        );

    \I__9471\ : Span4Mux_h
    port map (
            O => \N__43038\,
            I => \N__43025\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__43035\,
            I => \N__43018\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__43032\,
            I => \N__43018\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__43029\,
            I => \N__43018\
        );

    \I__9467\ : InMux
    port map (
            O => \N__43028\,
            I => \N__43015\
        );

    \I__9466\ : Span4Mux_h
    port map (
            O => \N__43025\,
            I => \N__43012\
        );

    \I__9465\ : Span4Mux_v
    port map (
            O => \N__43018\,
            I => \N__43009\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__43015\,
            I => eis_stop
        );

    \I__9463\ : Odrv4
    port map (
            O => \N__43012\,
            I => eis_stop
        );

    \I__9462\ : Odrv4
    port map (
            O => \N__43009\,
            I => eis_stop
        );

    \I__9461\ : InMux
    port map (
            O => \N__43002\,
            I => \N__42999\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__42999\,
            I => \N__42996\
        );

    \I__9459\ : Span4Mux_h
    port map (
            O => \N__42996\,
            I => \N__42991\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42995\,
            I => \N__42986\
        );

    \I__9457\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42986\
        );

    \I__9456\ : Odrv4
    port map (
            O => \N__42991\,
            I => req_data_cnt_9
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__42986\,
            I => req_data_cnt_9
        );

    \I__9454\ : InMux
    port map (
            O => \N__42981\,
            I => \N__42978\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__42978\,
            I => \N__42974\
        );

    \I__9452\ : InMux
    port map (
            O => \N__42977\,
            I => \N__42970\
        );

    \I__9451\ : Span12Mux_v
    port map (
            O => \N__42974\,
            I => \N__42967\
        );

    \I__9450\ : InMux
    port map (
            O => \N__42973\,
            I => \N__42964\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__42970\,
            I => \acadc_skipCount_9\
        );

    \I__9448\ : Odrv12
    port map (
            O => \N__42967\,
            I => \acadc_skipCount_9\
        );

    \I__9447\ : LocalMux
    port map (
            O => \N__42964\,
            I => \acadc_skipCount_9\
        );

    \I__9446\ : IoInMux
    port map (
            O => \N__42957\,
            I => \N__42954\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42954\,
            I => \N__42950\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42947\
        );

    \I__9443\ : Span12Mux_s0_v
    port map (
            O => \N__42950\,
            I => \N__42944\
        );

    \I__9442\ : LocalMux
    port map (
            O => \N__42947\,
            I => \N__42941\
        );

    \I__9441\ : Span12Mux_v
    port map (
            O => \N__42944\,
            I => \N__42938\
        );

    \I__9440\ : Span4Mux_v
    port map (
            O => \N__42941\,
            I => \N__42934\
        );

    \I__9439\ : Span12Mux_h
    port map (
            O => \N__42938\,
            I => \N__42931\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42928\
        );

    \I__9437\ : Span4Mux_h
    port map (
            O => \N__42934\,
            I => \N__42925\
        );

    \I__9436\ : Odrv12
    port map (
            O => \N__42931\,
            I => \DDS_RNG_0\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__42928\,
            I => \DDS_RNG_0\
        );

    \I__9434\ : Odrv4
    port map (
            O => \N__42925\,
            I => \DDS_RNG_0\
        );

    \I__9433\ : CascadeMux
    port map (
            O => \N__42918\,
            I => \n22617_cascade_\
        );

    \I__9432\ : CascadeMux
    port map (
            O => \N__42915\,
            I => \n22620_cascade_\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__9430\ : LocalMux
    port map (
            O => \N__42909\,
            I => n21360
        );

    \I__9429\ : InMux
    port map (
            O => \N__42906\,
            I => \N__42903\
        );

    \I__9428\ : LocalMux
    port map (
            O => \N__42903\,
            I => \N__42900\
        );

    \I__9427\ : Span4Mux_v
    port map (
            O => \N__42900\,
            I => \N__42897\
        );

    \I__9426\ : Sp12to4
    port map (
            O => \N__42897\,
            I => \N__42894\
        );

    \I__9425\ : Odrv12
    port map (
            O => \N__42894\,
            I => n22410
        );

    \I__9424\ : CascadeMux
    port map (
            O => \N__42891\,
            I => \n21361_cascade_\
        );

    \I__9423\ : SRMux
    port map (
            O => \N__42888\,
            I => \N__42884\
        );

    \I__9422\ : SRMux
    port map (
            O => \N__42887\,
            I => \N__42881\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__42884\,
            I => \N__42877\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42881\,
            I => \N__42874\
        );

    \I__9419\ : SRMux
    port map (
            O => \N__42880\,
            I => \N__42871\
        );

    \I__9418\ : Span4Mux_v
    port map (
            O => \N__42877\,
            I => \N__42866\
        );

    \I__9417\ : Span4Mux_v
    port map (
            O => \N__42874\,
            I => \N__42866\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__42871\,
            I => \N__42863\
        );

    \I__9415\ : Span4Mux_v
    port map (
            O => \N__42866\,
            I => \N__42860\
        );

    \I__9414\ : Span4Mux_v
    port map (
            O => \N__42863\,
            I => \N__42857\
        );

    \I__9413\ : Odrv4
    port map (
            O => \N__42860\,
            I => \comm_spi.data_tx_7__N_814\
        );

    \I__9412\ : Odrv4
    port map (
            O => \N__42857\,
            I => \comm_spi.data_tx_7__N_814\
        );

    \I__9411\ : CascadeMux
    port map (
            O => \N__42852\,
            I => \N__42848\
        );

    \I__9410\ : InMux
    port map (
            O => \N__42851\,
            I => \N__42840\
        );

    \I__9409\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42840\
        );

    \I__9408\ : InMux
    port map (
            O => \N__42847\,
            I => \N__42840\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42840\,
            I => comm_tx_buf_7
        );

    \I__9406\ : SRMux
    port map (
            O => \N__42837\,
            I => \N__42833\
        );

    \I__9405\ : SRMux
    port map (
            O => \N__42836\,
            I => \N__42830\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__42833\,
            I => \N__42826\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__42830\,
            I => \N__42823\
        );

    \I__9402\ : SRMux
    port map (
            O => \N__42829\,
            I => \N__42820\
        );

    \I__9401\ : Span4Mux_v
    port map (
            O => \N__42826\,
            I => \N__42815\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__42823\,
            I => \N__42815\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__42820\,
            I => \N__42812\
        );

    \I__9398\ : Span4Mux_v
    port map (
            O => \N__42815\,
            I => \N__42809\
        );

    \I__9397\ : Span4Mux_v
    port map (
            O => \N__42812\,
            I => \N__42806\
        );

    \I__9396\ : Odrv4
    port map (
            O => \N__42809\,
            I => \comm_spi.data_tx_7__N_806\
        );

    \I__9395\ : Odrv4
    port map (
            O => \N__42806\,
            I => \comm_spi.data_tx_7__N_806\
        );

    \I__9394\ : InMux
    port map (
            O => \N__42801\,
            I => \N__42798\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__42798\,
            I => \N__42792\
        );

    \I__9392\ : CascadeMux
    port map (
            O => \N__42797\,
            I => \N__42788\
        );

    \I__9391\ : CascadeMux
    port map (
            O => \N__42796\,
            I => \N__42785\
        );

    \I__9390\ : CascadeMux
    port map (
            O => \N__42795\,
            I => \N__42782\
        );

    \I__9389\ : Span4Mux_v
    port map (
            O => \N__42792\,
            I => \N__42775\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42772\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42757\
        );

    \I__9386\ : InMux
    port map (
            O => \N__42785\,
            I => \N__42757\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42782\,
            I => \N__42757\
        );

    \I__9384\ : InMux
    port map (
            O => \N__42781\,
            I => \N__42757\
        );

    \I__9383\ : InMux
    port map (
            O => \N__42780\,
            I => \N__42757\
        );

    \I__9382\ : InMux
    port map (
            O => \N__42779\,
            I => \N__42757\
        );

    \I__9381\ : InMux
    port map (
            O => \N__42778\,
            I => \N__42757\
        );

    \I__9380\ : Odrv4
    port map (
            O => \N__42775\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__42772\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__42757\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__9377\ : InMux
    port map (
            O => \N__42750\,
            I => \N__42747\
        );

    \I__9376\ : LocalMux
    port map (
            O => \N__42747\,
            I => \N__42737\
        );

    \I__9375\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42722\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42745\,
            I => \N__42722\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42744\,
            I => \N__42722\
        );

    \I__9372\ : InMux
    port map (
            O => \N__42743\,
            I => \N__42722\
        );

    \I__9371\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42722\
        );

    \I__9370\ : InMux
    port map (
            O => \N__42741\,
            I => \N__42722\
        );

    \I__9369\ : InMux
    port map (
            O => \N__42740\,
            I => \N__42722\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__42737\,
            I => \comm_spi.n17254\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__42722\,
            I => \comm_spi.n17254\
        );

    \I__9366\ : CascadeMux
    port map (
            O => \N__42717\,
            I => \n22551_cascade_\
        );

    \I__9365\ : CascadeMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__9364\ : InMux
    port map (
            O => \N__42711\,
            I => \N__42704\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42701\
        );

    \I__9362\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42698\
        );

    \I__9361\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42695\
        );

    \I__9360\ : CascadeMux
    port map (
            O => \N__42707\,
            I => \N__42692\
        );

    \I__9359\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42689\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__42701\,
            I => \N__42686\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__42698\,
            I => \N__42683\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__42695\,
            I => \N__42680\
        );

    \I__9355\ : InMux
    port map (
            O => \N__42692\,
            I => \N__42677\
        );

    \I__9354\ : Span4Mux_h
    port map (
            O => \N__42689\,
            I => \N__42672\
        );

    \I__9353\ : Span4Mux_h
    port map (
            O => \N__42686\,
            I => \N__42672\
        );

    \I__9352\ : Span4Mux_v
    port map (
            O => \N__42683\,
            I => \N__42669\
        );

    \I__9351\ : Span4Mux_h
    port map (
            O => \N__42680\,
            I => \N__42666\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__42677\,
            I => \N__42663\
        );

    \I__9349\ : Span4Mux_h
    port map (
            O => \N__42672\,
            I => \N__42660\
        );

    \I__9348\ : Span4Mux_h
    port map (
            O => \N__42669\,
            I => \N__42655\
        );

    \I__9347\ : Span4Mux_v
    port map (
            O => \N__42666\,
            I => \N__42655\
        );

    \I__9346\ : Odrv4
    port map (
            O => \N__42663\,
            I => comm_buf_1_4
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__42660\,
            I => comm_buf_1_4
        );

    \I__9344\ : Odrv4
    port map (
            O => \N__42655\,
            I => comm_buf_1_4
        );

    \I__9343\ : CascadeMux
    port map (
            O => \N__42648\,
            I => \n4_adj_1582_cascade_\
        );

    \I__9342\ : CascadeMux
    port map (
            O => \N__42645\,
            I => \n21285_cascade_\
        );

    \I__9341\ : InMux
    port map (
            O => \N__42642\,
            I => \N__42639\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__42639\,
            I => n22554
        );

    \I__9339\ : CEMux
    port map (
            O => \N__42636\,
            I => \N__42632\
        );

    \I__9338\ : CEMux
    port map (
            O => \N__42635\,
            I => \N__42627\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__42632\,
            I => \N__42624\
        );

    \I__9336\ : CEMux
    port map (
            O => \N__42631\,
            I => \N__42621\
        );

    \I__9335\ : CEMux
    port map (
            O => \N__42630\,
            I => \N__42618\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__42627\,
            I => \N__42615\
        );

    \I__9333\ : Span4Mux_v
    port map (
            O => \N__42624\,
            I => \N__42612\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__42621\,
            I => \N__42609\
        );

    \I__9331\ : LocalMux
    port map (
            O => \N__42618\,
            I => \N__42606\
        );

    \I__9330\ : Span4Mux_h
    port map (
            O => \N__42615\,
            I => \N__42601\
        );

    \I__9329\ : Span4Mux_h
    port map (
            O => \N__42612\,
            I => \N__42601\
        );

    \I__9328\ : Span4Mux_h
    port map (
            O => \N__42609\,
            I => \N__42598\
        );

    \I__9327\ : Span4Mux_h
    port map (
            O => \N__42606\,
            I => \N__42595\
        );

    \I__9326\ : Odrv4
    port map (
            O => \N__42601\,
            I => n11910
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__42598\,
            I => n11910
        );

    \I__9324\ : Odrv4
    port map (
            O => \N__42595\,
            I => n11910
        );

    \I__9323\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42585\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__42585\,
            I => \N__42582\
        );

    \I__9321\ : Span4Mux_v
    port map (
            O => \N__42582\,
            I => \N__42579\
        );

    \I__9320\ : Span4Mux_v
    port map (
            O => \N__42579\,
            I => \N__42576\
        );

    \I__9319\ : Span4Mux_h
    port map (
            O => \N__42576\,
            I => \N__42573\
        );

    \I__9318\ : Odrv4
    port map (
            O => \N__42573\,
            I => buf_data_iac_10
        );

    \I__9317\ : InMux
    port map (
            O => \N__42570\,
            I => \N__42567\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__42567\,
            I => \N__42564\
        );

    \I__9315\ : Span4Mux_v
    port map (
            O => \N__42564\,
            I => \N__42561\
        );

    \I__9314\ : Span4Mux_h
    port map (
            O => \N__42561\,
            I => \N__42558\
        );

    \I__9313\ : Odrv4
    port map (
            O => \N__42558\,
            I => n21385
        );

    \I__9312\ : InMux
    port map (
            O => \N__42555\,
            I => \N__42551\
        );

    \I__9311\ : CascadeMux
    port map (
            O => \N__42554\,
            I => \N__42547\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__42551\,
            I => \N__42544\
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__42550\,
            I => \N__42539\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42547\,
            I => \N__42536\
        );

    \I__9307\ : Span4Mux_h
    port map (
            O => \N__42544\,
            I => \N__42532\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42527\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42542\,
            I => \N__42527\
        );

    \I__9304\ : InMux
    port map (
            O => \N__42539\,
            I => \N__42524\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__42536\,
            I => \N__42521\
        );

    \I__9302\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42518\
        );

    \I__9301\ : Sp12to4
    port map (
            O => \N__42532\,
            I => \N__42512\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__42527\,
            I => \N__42512\
        );

    \I__9299\ : LocalMux
    port map (
            O => \N__42524\,
            I => \N__42509\
        );

    \I__9298\ : Span4Mux_v
    port map (
            O => \N__42521\,
            I => \N__42504\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__42518\,
            I => \N__42504\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42517\,
            I => \N__42501\
        );

    \I__9295\ : Span12Mux_v
    port map (
            O => \N__42512\,
            I => \N__42498\
        );

    \I__9294\ : Span4Mux_v
    port map (
            O => \N__42509\,
            I => \N__42495\
        );

    \I__9293\ : Span4Mux_h
    port map (
            O => \N__42504\,
            I => \N__42490\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__42501\,
            I => \N__42490\
        );

    \I__9291\ : Odrv12
    port map (
            O => \N__42498\,
            I => comm_buf_0_7
        );

    \I__9290\ : Odrv4
    port map (
            O => \N__42495\,
            I => comm_buf_0_7
        );

    \I__9289\ : Odrv4
    port map (
            O => \N__42490\,
            I => comm_buf_0_7
        );

    \I__9288\ : InMux
    port map (
            O => \N__42483\,
            I => \N__42480\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__42480\,
            I => \N__42477\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__42477\,
            I => n21276
        );

    \I__9285\ : CascadeMux
    port map (
            O => \N__42474\,
            I => \n22542_cascade_\
        );

    \I__9284\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42468\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__42468\,
            I => \N__42465\
        );

    \I__9282\ : Odrv4
    port map (
            O => \N__42465\,
            I => n4_adj_1580
        );

    \I__9281\ : IoInMux
    port map (
            O => \N__42462\,
            I => \N__42459\
        );

    \I__9280\ : LocalMux
    port map (
            O => \N__42459\,
            I => \N__42456\
        );

    \I__9279\ : IoSpan4Mux
    port map (
            O => \N__42456\,
            I => \N__42453\
        );

    \I__9278\ : Span4Mux_s0_h
    port map (
            O => \N__42453\,
            I => \N__42450\
        );

    \I__9277\ : Sp12to4
    port map (
            O => \N__42450\,
            I => \N__42447\
        );

    \I__9276\ : Span12Mux_h
    port map (
            O => \N__42447\,
            I => \N__42443\
        );

    \I__9275\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42440\
        );

    \I__9274\ : Odrv12
    port map (
            O => \N__42443\,
            I => \VDC_SCLK\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__42440\,
            I => \VDC_SCLK\
        );

    \I__9272\ : IoInMux
    port map (
            O => \N__42435\,
            I => \N__42431\
        );

    \I__9271\ : ClkMux
    port map (
            O => \N__42434\,
            I => \N__42426\
        );

    \I__9270\ : LocalMux
    port map (
            O => \N__42431\,
            I => \N__42421\
        );

    \I__9269\ : ClkMux
    port map (
            O => \N__42430\,
            I => \N__42418\
        );

    \I__9268\ : ClkMux
    port map (
            O => \N__42429\,
            I => \N__42415\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__42426\,
            I => \N__42406\
        );

    \I__9266\ : ClkMux
    port map (
            O => \N__42425\,
            I => \N__42403\
        );

    \I__9265\ : ClkMux
    port map (
            O => \N__42424\,
            I => \N__42400\
        );

    \I__9264\ : Span4Mux_s1_h
    port map (
            O => \N__42421\,
            I => \N__42395\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__42418\,
            I => \N__42391\
        );

    \I__9262\ : LocalMux
    port map (
            O => \N__42415\,
            I => \N__42388\
        );

    \I__9261\ : ClkMux
    port map (
            O => \N__42414\,
            I => \N__42385\
        );

    \I__9260\ : ClkMux
    port map (
            O => \N__42413\,
            I => \N__42380\
        );

    \I__9259\ : ClkMux
    port map (
            O => \N__42412\,
            I => \N__42377\
        );

    \I__9258\ : ClkMux
    port map (
            O => \N__42411\,
            I => \N__42374\
        );

    \I__9257\ : ClkMux
    port map (
            O => \N__42410\,
            I => \N__42369\
        );

    \I__9256\ : ClkMux
    port map (
            O => \N__42409\,
            I => \N__42366\
        );

    \I__9255\ : Span4Mux_h
    port map (
            O => \N__42406\,
            I => \N__42357\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__42403\,
            I => \N__42357\
        );

    \I__9253\ : LocalMux
    port map (
            O => \N__42400\,
            I => \N__42354\
        );

    \I__9252\ : ClkMux
    port map (
            O => \N__42399\,
            I => \N__42351\
        );

    \I__9251\ : ClkMux
    port map (
            O => \N__42398\,
            I => \N__42348\
        );

    \I__9250\ : Span4Mux_h
    port map (
            O => \N__42395\,
            I => \N__42345\
        );

    \I__9249\ : ClkMux
    port map (
            O => \N__42394\,
            I => \N__42342\
        );

    \I__9248\ : Span4Mux_v
    port map (
            O => \N__42391\,
            I => \N__42335\
        );

    \I__9247\ : Span4Mux_v
    port map (
            O => \N__42388\,
            I => \N__42335\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__42385\,
            I => \N__42335\
        );

    \I__9245\ : ClkMux
    port map (
            O => \N__42384\,
            I => \N__42331\
        );

    \I__9244\ : ClkMux
    port map (
            O => \N__42383\,
            I => \N__42328\
        );

    \I__9243\ : LocalMux
    port map (
            O => \N__42380\,
            I => \N__42325\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__42377\,
            I => \N__42320\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42374\,
            I => \N__42320\
        );

    \I__9240\ : ClkMux
    port map (
            O => \N__42373\,
            I => \N__42317\
        );

    \I__9239\ : ClkMux
    port map (
            O => \N__42372\,
            I => \N__42314\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__42369\,
            I => \N__42309\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__42366\,
            I => \N__42309\
        );

    \I__9236\ : ClkMux
    port map (
            O => \N__42365\,
            I => \N__42306\
        );

    \I__9235\ : ClkMux
    port map (
            O => \N__42364\,
            I => \N__42302\
        );

    \I__9234\ : ClkMux
    port map (
            O => \N__42363\,
            I => \N__42298\
        );

    \I__9233\ : ClkMux
    port map (
            O => \N__42362\,
            I => \N__42295\
        );

    \I__9232\ : Span4Mux_v
    port map (
            O => \N__42357\,
            I => \N__42286\
        );

    \I__9231\ : Span4Mux_h
    port map (
            O => \N__42354\,
            I => \N__42286\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__42351\,
            I => \N__42286\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__42348\,
            I => \N__42286\
        );

    \I__9228\ : Span4Mux_h
    port map (
            O => \N__42345\,
            I => \N__42279\
        );

    \I__9227\ : LocalMux
    port map (
            O => \N__42342\,
            I => \N__42279\
        );

    \I__9226\ : Span4Mux_h
    port map (
            O => \N__42335\,
            I => \N__42279\
        );

    \I__9225\ : ClkMux
    port map (
            O => \N__42334\,
            I => \N__42276\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__42331\,
            I => \N__42269\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__42328\,
            I => \N__42269\
        );

    \I__9222\ : Span4Mux_v
    port map (
            O => \N__42325\,
            I => \N__42269\
        );

    \I__9221\ : Span4Mux_v
    port map (
            O => \N__42320\,
            I => \N__42264\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__42317\,
            I => \N__42264\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__42314\,
            I => \N__42261\
        );

    \I__9218\ : Span4Mux_v
    port map (
            O => \N__42309\,
            I => \N__42256\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__42306\,
            I => \N__42256\
        );

    \I__9216\ : ClkMux
    port map (
            O => \N__42305\,
            I => \N__42253\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__42302\,
            I => \N__42250\
        );

    \I__9214\ : ClkMux
    port map (
            O => \N__42301\,
            I => \N__42247\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__42298\,
            I => \N__42244\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__42295\,
            I => \N__42235\
        );

    \I__9211\ : Span4Mux_v
    port map (
            O => \N__42286\,
            I => \N__42235\
        );

    \I__9210\ : Span4Mux_h
    port map (
            O => \N__42279\,
            I => \N__42235\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__42276\,
            I => \N__42235\
        );

    \I__9208\ : Span4Mux_v
    port map (
            O => \N__42269\,
            I => \N__42230\
        );

    \I__9207\ : Span4Mux_h
    port map (
            O => \N__42264\,
            I => \N__42230\
        );

    \I__9206\ : Span4Mux_v
    port map (
            O => \N__42261\,
            I => \N__42227\
        );

    \I__9205\ : Span4Mux_h
    port map (
            O => \N__42256\,
            I => \N__42222\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__42253\,
            I => \N__42222\
        );

    \I__9203\ : Span4Mux_h
    port map (
            O => \N__42250\,
            I => \N__42218\
        );

    \I__9202\ : LocalMux
    port map (
            O => \N__42247\,
            I => \N__42215\
        );

    \I__9201\ : Span4Mux_v
    port map (
            O => \N__42244\,
            I => \N__42212\
        );

    \I__9200\ : Span4Mux_h
    port map (
            O => \N__42235\,
            I => \N__42209\
        );

    \I__9199\ : Span4Mux_h
    port map (
            O => \N__42230\,
            I => \N__42204\
        );

    \I__9198\ : Span4Mux_v
    port map (
            O => \N__42227\,
            I => \N__42204\
        );

    \I__9197\ : Span4Mux_h
    port map (
            O => \N__42222\,
            I => \N__42201\
        );

    \I__9196\ : ClkMux
    port map (
            O => \N__42221\,
            I => \N__42198\
        );

    \I__9195\ : Odrv4
    port map (
            O => \N__42218\,
            I => \VDC_CLK\
        );

    \I__9194\ : Odrv12
    port map (
            O => \N__42215\,
            I => \VDC_CLK\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__42212\,
            I => \VDC_CLK\
        );

    \I__9192\ : Odrv4
    port map (
            O => \N__42209\,
            I => \VDC_CLK\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__42204\,
            I => \VDC_CLK\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__42201\,
            I => \VDC_CLK\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__42198\,
            I => \VDC_CLK\
        );

    \I__9188\ : InMux
    port map (
            O => \N__42183\,
            I => \N__42180\
        );

    \I__9187\ : LocalMux
    port map (
            O => \N__42180\,
            I => \N__42177\
        );

    \I__9186\ : Span4Mux_h
    port map (
            O => \N__42177\,
            I => \N__42174\
        );

    \I__9185\ : Span4Mux_h
    port map (
            O => \N__42174\,
            I => \N__42171\
        );

    \I__9184\ : Odrv4
    port map (
            O => \N__42171\,
            I => buf_data_iac_20
        );

    \I__9183\ : InMux
    port map (
            O => \N__42168\,
            I => \N__42165\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__42165\,
            I => \N__42162\
        );

    \I__9181\ : Span4Mux_h
    port map (
            O => \N__42162\,
            I => \N__42159\
        );

    \I__9180\ : Span4Mux_v
    port map (
            O => \N__42159\,
            I => \N__42156\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__42156\,
            I => n21557
        );

    \I__9178\ : SRMux
    port map (
            O => \N__42153\,
            I => \N__42148\
        );

    \I__9177\ : SRMux
    port map (
            O => \N__42152\,
            I => \N__42144\
        );

    \I__9176\ : SRMux
    port map (
            O => \N__42151\,
            I => \N__42140\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__42148\,
            I => \N__42137\
        );

    \I__9174\ : SRMux
    port map (
            O => \N__42147\,
            I => \N__42134\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__42144\,
            I => \N__42131\
        );

    \I__9172\ : SRMux
    port map (
            O => \N__42143\,
            I => \N__42128\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__42140\,
            I => \N__42125\
        );

    \I__9170\ : Span4Mux_v
    port map (
            O => \N__42137\,
            I => \N__42120\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__42134\,
            I => \N__42120\
        );

    \I__9168\ : Span4Mux_h
    port map (
            O => \N__42131\,
            I => \N__42115\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__42128\,
            I => \N__42115\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__42125\,
            I => \N__42112\
        );

    \I__9165\ : Span4Mux_h
    port map (
            O => \N__42120\,
            I => \N__42109\
        );

    \I__9164\ : Odrv4
    port map (
            O => \N__42115\,
            I => flagcntwd
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__42112\,
            I => flagcntwd
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__42109\,
            I => flagcntwd
        );

    \I__9161\ : CascadeMux
    port map (
            O => \N__42102\,
            I => \n21187_cascade_\
        );

    \I__9160\ : CEMux
    port map (
            O => \N__42099\,
            I => \N__42096\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__42096\,
            I => n11605
        );

    \I__9158\ : SRMux
    port map (
            O => \N__42093\,
            I => \N__42090\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__42090\,
            I => \N__42087\
        );

    \I__9156\ : Span4Mux_h
    port map (
            O => \N__42087\,
            I => \N__42084\
        );

    \I__9155\ : Span4Mux_h
    port map (
            O => \N__42084\,
            I => \N__42080\
        );

    \I__9154\ : SRMux
    port map (
            O => \N__42083\,
            I => \N__42077\
        );

    \I__9153\ : Odrv4
    port map (
            O => \N__42080\,
            I => n20578
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__42077\,
            I => n20578
        );

    \I__9151\ : CascadeMux
    port map (
            O => \N__42072\,
            I => \n11576_cascade_\
        );

    \I__9150\ : CEMux
    port map (
            O => \N__42069\,
            I => \N__42066\
        );

    \I__9149\ : LocalMux
    port map (
            O => \N__42066\,
            I => \N__42063\
        );

    \I__9148\ : Span4Mux_h
    port map (
            O => \N__42063\,
            I => \N__42060\
        );

    \I__9147\ : Span4Mux_h
    port map (
            O => \N__42060\,
            I => \N__42057\
        );

    \I__9146\ : Odrv4
    port map (
            O => \N__42057\,
            I => n12148
        );

    \I__9145\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42051\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__42051\,
            I => \N__42047\
        );

    \I__9143\ : InMux
    port map (
            O => \N__42050\,
            I => \N__42043\
        );

    \I__9142\ : Span4Mux_v
    port map (
            O => \N__42047\,
            I => \N__42040\
        );

    \I__9141\ : CascadeMux
    port map (
            O => \N__42046\,
            I => \N__42037\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__42043\,
            I => \N__42032\
        );

    \I__9139\ : Span4Mux_h
    port map (
            O => \N__42040\,
            I => \N__42032\
        );

    \I__9138\ : InMux
    port map (
            O => \N__42037\,
            I => \N__42029\
        );

    \I__9137\ : Span4Mux_h
    port map (
            O => \N__42032\,
            I => \N__42026\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__42029\,
            I => buf_adcdata_iac_15
        );

    \I__9135\ : Odrv4
    port map (
            O => \N__42026\,
            I => buf_adcdata_iac_15
        );

    \I__9134\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42018\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__42018\,
            I => \N__42015\
        );

    \I__9132\ : Span4Mux_h
    port map (
            O => \N__42015\,
            I => \N__42012\
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__42012\,
            I => n16_adj_1620
        );

    \I__9130\ : CascadeMux
    port map (
            O => \N__42009\,
            I => \N__42005\
        );

    \I__9129\ : InMux
    port map (
            O => \N__42008\,
            I => \N__42002\
        );

    \I__9128\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41998\
        );

    \I__9127\ : LocalMux
    port map (
            O => \N__42002\,
            I => \N__41995\
        );

    \I__9126\ : InMux
    port map (
            O => \N__42001\,
            I => \N__41992\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41998\,
            I => \N__41985\
        );

    \I__9124\ : Span4Mux_h
    port map (
            O => \N__41995\,
            I => \N__41982\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__41992\,
            I => \N__41979\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41991\,
            I => \N__41974\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41974\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41969\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41969\
        );

    \I__9118\ : Span4Mux_h
    port map (
            O => \N__41985\,
            I => \N__41966\
        );

    \I__9117\ : Sp12to4
    port map (
            O => \N__41982\,
            I => \N__41963\
        );

    \I__9116\ : Sp12to4
    port map (
            O => \N__41979\,
            I => \N__41960\
        );

    \I__9115\ : LocalMux
    port map (
            O => \N__41974\,
            I => n12144
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41969\,
            I => n12144
        );

    \I__9113\ : Odrv4
    port map (
            O => \N__41966\,
            I => n12144
        );

    \I__9112\ : Odrv12
    port map (
            O => \N__41963\,
            I => n12144
        );

    \I__9111\ : Odrv12
    port map (
            O => \N__41960\,
            I => n12144
        );

    \I__9110\ : IoInMux
    port map (
            O => \N__41949\,
            I => \N__41946\
        );

    \I__9109\ : LocalMux
    port map (
            O => \N__41946\,
            I => \N__41943\
        );

    \I__9108\ : Span12Mux_s0_v
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__9107\ : Span12Mux_h
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__9106\ : Odrv12
    port map (
            O => \N__41937\,
            I => \DDS_CS\
        );

    \I__9105\ : CEMux
    port map (
            O => \N__41934\,
            I => \N__41931\
        );

    \I__9104\ : LocalMux
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__9103\ : Span4Mux_h
    port map (
            O => \N__41928\,
            I => \N__41925\
        );

    \I__9102\ : Odrv4
    port map (
            O => \N__41925\,
            I => \SIG_DDS.n9_adj_1434\
        );

    \I__9101\ : CascadeMux
    port map (
            O => \N__41922\,
            I => \N__41919\
        );

    \I__9100\ : InMux
    port map (
            O => \N__41919\,
            I => \N__41916\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__41916\,
            I => \N__41912\
        );

    \I__9098\ : InMux
    port map (
            O => \N__41915\,
            I => \N__41909\
        );

    \I__9097\ : Odrv4
    port map (
            O => \N__41912\,
            I => n8_adj_1556
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__41909\,
            I => n8_adj_1556
        );

    \I__9095\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41901\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41901\,
            I => \N__41897\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41900\,
            I => \N__41894\
        );

    \I__9092\ : Span4Mux_v
    port map (
            O => \N__41897\,
            I => \N__41891\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__41894\,
            I => n7_adj_1555
        );

    \I__9090\ : Odrv4
    port map (
            O => \N__41891\,
            I => n7_adj_1555
        );

    \I__9089\ : CascadeMux
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__9088\ : CascadeBuf
    port map (
            O => \N__41883\,
            I => \N__41880\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__41880\,
            I => \N__41877\
        );

    \I__9086\ : CascadeBuf
    port map (
            O => \N__41877\,
            I => \N__41874\
        );

    \I__9085\ : CascadeMux
    port map (
            O => \N__41874\,
            I => \N__41871\
        );

    \I__9084\ : CascadeBuf
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__9083\ : CascadeMux
    port map (
            O => \N__41868\,
            I => \N__41865\
        );

    \I__9082\ : CascadeBuf
    port map (
            O => \N__41865\,
            I => \N__41862\
        );

    \I__9081\ : CascadeMux
    port map (
            O => \N__41862\,
            I => \N__41859\
        );

    \I__9080\ : CascadeBuf
    port map (
            O => \N__41859\,
            I => \N__41856\
        );

    \I__9079\ : CascadeMux
    port map (
            O => \N__41856\,
            I => \N__41853\
        );

    \I__9078\ : CascadeBuf
    port map (
            O => \N__41853\,
            I => \N__41850\
        );

    \I__9077\ : CascadeMux
    port map (
            O => \N__41850\,
            I => \N__41847\
        );

    \I__9076\ : CascadeBuf
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__9075\ : CascadeMux
    port map (
            O => \N__41844\,
            I => \N__41840\
        );

    \I__9074\ : CascadeMux
    port map (
            O => \N__41843\,
            I => \N__41837\
        );

    \I__9073\ : CascadeBuf
    port map (
            O => \N__41840\,
            I => \N__41834\
        );

    \I__9072\ : CascadeBuf
    port map (
            O => \N__41837\,
            I => \N__41831\
        );

    \I__9071\ : CascadeMux
    port map (
            O => \N__41834\,
            I => \N__41828\
        );

    \I__9070\ : CascadeMux
    port map (
            O => \N__41831\,
            I => \N__41825\
        );

    \I__9069\ : CascadeBuf
    port map (
            O => \N__41828\,
            I => \N__41822\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41819\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__41822\,
            I => \N__41816\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__41819\,
            I => \N__41813\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41816\,
            I => \N__41810\
        );

    \I__9064\ : Span12Mux_h
    port map (
            O => \N__41813\,
            I => \N__41807\
        );

    \I__9063\ : LocalMux
    port map (
            O => \N__41810\,
            I => \N__41804\
        );

    \I__9062\ : Odrv12
    port map (
            O => \N__41807\,
            I => \data_index_9_N_212_9\
        );

    \I__9061\ : Odrv12
    port map (
            O => \N__41804\,
            I => \data_index_9_N_212_9\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41795\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41792\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41795\,
            I => \comm_spi.n14818\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__41792\,
            I => \comm_spi.n14818\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41784\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41784\,
            I => \N__41780\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41783\,
            I => \N__41777\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__41780\,
            I => \N__41772\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41777\,
            I => \N__41772\
        );

    \I__9051\ : Odrv4
    port map (
            O => \N__41772\,
            I => \comm_spi.n14819\
        );

    \I__9050\ : InMux
    port map (
            O => \N__41769\,
            I => \N__41766\
        );

    \I__9049\ : LocalMux
    port map (
            O => \N__41766\,
            I => \N__41763\
        );

    \I__9048\ : Span4Mux_h
    port map (
            O => \N__41763\,
            I => \N__41760\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__41760\,
            I => \N__41757\
        );

    \I__9046\ : Odrv4
    port map (
            O => \N__41757\,
            I => buf_data_iac_21
        );

    \I__9045\ : InMux
    port map (
            O => \N__41754\,
            I => \N__41751\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__41751\,
            I => \N__41748\
        );

    \I__9043\ : Span4Mux_h
    port map (
            O => \N__41748\,
            I => \N__41745\
        );

    \I__9042\ : Span4Mux_v
    port map (
            O => \N__41745\,
            I => \N__41742\
        );

    \I__9041\ : Odrv4
    port map (
            O => \N__41742\,
            I => n21672
        );

    \I__9040\ : CascadeMux
    port map (
            O => \N__41739\,
            I => \ADC_VDC.n22124_cascade_\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__41736\,
            I => \N__41733\
        );

    \I__9038\ : InMux
    port map (
            O => \N__41733\,
            I => \N__41730\
        );

    \I__9037\ : LocalMux
    port map (
            O => \N__41730\,
            I => \N__41727\
        );

    \I__9036\ : Span4Mux_h
    port map (
            O => \N__41727\,
            I => \N__41724\
        );

    \I__9035\ : Span4Mux_h
    port map (
            O => \N__41724\,
            I => \N__41719\
        );

    \I__9034\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41714\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41714\
        );

    \I__9032\ : Odrv4
    port map (
            O => \N__41719\,
            I => buf_dds1_0
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41714\,
            I => buf_dds1_0
        );

    \I__9030\ : CascadeMux
    port map (
            O => \N__41709\,
            I => \n16_cascade_\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41706\,
            I => \N__41702\
        );

    \I__9028\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41698\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__41702\,
            I => \N__41695\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__41701\,
            I => \N__41692\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41698\,
            I => \N__41689\
        );

    \I__9024\ : Span4Mux_v
    port map (
            O => \N__41695\,
            I => \N__41686\
        );

    \I__9023\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41683\
        );

    \I__9022\ : Span4Mux_v
    port map (
            O => \N__41689\,
            I => \N__41680\
        );

    \I__9021\ : Sp12to4
    port map (
            O => \N__41686\,
            I => \N__41677\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__41683\,
            I => buf_adcdata_iac_8
        );

    \I__9019\ : Odrv4
    port map (
            O => \N__41680\,
            I => buf_adcdata_iac_8
        );

    \I__9018\ : Odrv12
    port map (
            O => \N__41677\,
            I => buf_adcdata_iac_8
        );

    \I__9017\ : CascadeMux
    port map (
            O => \N__41670\,
            I => \N__41659\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41669\,
            I => \N__41654\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41668\,
            I => \N__41651\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41648\
        );

    \I__9013\ : InMux
    port map (
            O => \N__41666\,
            I => \N__41645\
        );

    \I__9012\ : InMux
    port map (
            O => \N__41665\,
            I => \N__41641\
        );

    \I__9011\ : InMux
    port map (
            O => \N__41664\,
            I => \N__41638\
        );

    \I__9010\ : InMux
    port map (
            O => \N__41663\,
            I => \N__41634\
        );

    \I__9009\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41631\
        );

    \I__9008\ : InMux
    port map (
            O => \N__41659\,
            I => \N__41628\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41658\,
            I => \N__41625\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41622\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__41654\,
            I => \N__41619\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__41651\,
            I => \N__41616\
        );

    \I__9003\ : LocalMux
    port map (
            O => \N__41648\,
            I => \N__41610\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__41645\,
            I => \N__41607\
        );

    \I__9001\ : InMux
    port map (
            O => \N__41644\,
            I => \N__41604\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41641\,
            I => \N__41599\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41638\,
            I => \N__41599\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41637\,
            I => \N__41596\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__41634\,
            I => \N__41591\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__41631\,
            I => \N__41591\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__41628\,
            I => \N__41584\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__41625\,
            I => \N__41584\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__41622\,
            I => \N__41584\
        );

    \I__8992\ : Span4Mux_v
    port map (
            O => \N__41619\,
            I => \N__41579\
        );

    \I__8991\ : Span4Mux_h
    port map (
            O => \N__41616\,
            I => \N__41579\
        );

    \I__8990\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41574\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41574\
        );

    \I__8988\ : InMux
    port map (
            O => \N__41613\,
            I => \N__41571\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__41610\,
            I => \N__41568\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__41607\,
            I => \N__41565\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__41604\,
            I => \N__41560\
        );

    \I__8984\ : Span4Mux_h
    port map (
            O => \N__41599\,
            I => \N__41560\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__41596\,
            I => \N__41551\
        );

    \I__8982\ : Span4Mux_h
    port map (
            O => \N__41591\,
            I => \N__41551\
        );

    \I__8981\ : Span4Mux_v
    port map (
            O => \N__41584\,
            I => \N__41551\
        );

    \I__8980\ : Span4Mux_v
    port map (
            O => \N__41579\,
            I => \N__41551\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__41574\,
            I => n12596
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__41571\,
            I => n12596
        );

    \I__8977\ : Odrv4
    port map (
            O => \N__41568\,
            I => n12596
        );

    \I__8976\ : Odrv4
    port map (
            O => \N__41565\,
            I => n12596
        );

    \I__8975\ : Odrv4
    port map (
            O => \N__41560\,
            I => n12596
        );

    \I__8974\ : Odrv4
    port map (
            O => \N__41551\,
            I => n12596
        );

    \I__8973\ : InMux
    port map (
            O => \N__41538\,
            I => \N__41535\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__41535\,
            I => \N__41532\
        );

    \I__8971\ : Span4Mux_v
    port map (
            O => \N__41532\,
            I => \N__41527\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41531\,
            I => \N__41522\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41530\,
            I => \N__41522\
        );

    \I__8968\ : Odrv4
    port map (
            O => \N__41527\,
            I => buf_dds0_0
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__41522\,
            I => buf_dds0_0
        );

    \I__8966\ : IoInMux
    port map (
            O => \N__41517\,
            I => \N__41514\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__41514\,
            I => \N__41511\
        );

    \I__8964\ : Span4Mux_s2_h
    port map (
            O => \N__41511\,
            I => \N__41508\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__41508\,
            I => \N__41505\
        );

    \I__8962\ : Sp12to4
    port map (
            O => \N__41505\,
            I => \N__41502\
        );

    \I__8961\ : Span12Mux_v
    port map (
            O => \N__41502\,
            I => \N__41498\
        );

    \I__8960\ : CascadeMux
    port map (
            O => \N__41501\,
            I => \N__41494\
        );

    \I__8959\ : Span12Mux_h
    port map (
            O => \N__41498\,
            I => \N__41491\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41497\,
            I => \N__41488\
        );

    \I__8957\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41485\
        );

    \I__8956\ : Odrv12
    port map (
            O => \N__41491\,
            I => \VDC_RNG0\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__41488\,
            I => \VDC_RNG0\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__41485\,
            I => \VDC_RNG0\
        );

    \I__8953\ : CascadeMux
    port map (
            O => \N__41478\,
            I => \N__41475\
        );

    \I__8952\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41472\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__41472\,
            I => \N__41469\
        );

    \I__8950\ : Span4Mux_v
    port map (
            O => \N__41469\,
            I => \N__41466\
        );

    \I__8949\ : Odrv4
    port map (
            O => \N__41466\,
            I => n23_adj_1675
        );

    \I__8948\ : InMux
    port map (
            O => \N__41463\,
            I => \N__41460\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__41460\,
            I => \N__41457\
        );

    \I__8946\ : Span4Mux_v
    port map (
            O => \N__41457\,
            I => \N__41452\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41456\,
            I => \N__41449\
        );

    \I__8944\ : InMux
    port map (
            O => \N__41455\,
            I => \N__41446\
        );

    \I__8943\ : Odrv4
    port map (
            O => \N__41452\,
            I => buf_dds0_6
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__41449\,
            I => buf_dds0_6
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__41446\,
            I => buf_dds0_6
        );

    \I__8940\ : InMux
    port map (
            O => \N__41439\,
            I => \N__41435\
        );

    \I__8939\ : InMux
    port map (
            O => \N__41438\,
            I => \N__41432\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__41435\,
            I => n17705
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__41432\,
            I => n17705
        );

    \I__8936\ : CascadeMux
    port map (
            O => \N__41427\,
            I => \n9342_cascade_\
        );

    \I__8935\ : CascadeMux
    port map (
            O => \N__41424\,
            I => \N__41421\
        );

    \I__8934\ : InMux
    port map (
            O => \N__41421\,
            I => \N__41418\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41418\,
            I => \N__41414\
        );

    \I__8932\ : InMux
    port map (
            O => \N__41417\,
            I => \N__41411\
        );

    \I__8931\ : Odrv4
    port map (
            O => \N__41414\,
            I => n17703
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__41411\,
            I => n17703
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__41406\,
            I => \N__41403\
        );

    \I__8928\ : CascadeBuf
    port map (
            O => \N__41403\,
            I => \N__41400\
        );

    \I__8927\ : CascadeMux
    port map (
            O => \N__41400\,
            I => \N__41397\
        );

    \I__8926\ : CascadeBuf
    port map (
            O => \N__41397\,
            I => \N__41394\
        );

    \I__8925\ : CascadeMux
    port map (
            O => \N__41394\,
            I => \N__41391\
        );

    \I__8924\ : CascadeBuf
    port map (
            O => \N__41391\,
            I => \N__41388\
        );

    \I__8923\ : CascadeMux
    port map (
            O => \N__41388\,
            I => \N__41385\
        );

    \I__8922\ : CascadeBuf
    port map (
            O => \N__41385\,
            I => \N__41382\
        );

    \I__8921\ : CascadeMux
    port map (
            O => \N__41382\,
            I => \N__41379\
        );

    \I__8920\ : CascadeBuf
    port map (
            O => \N__41379\,
            I => \N__41376\
        );

    \I__8919\ : CascadeMux
    port map (
            O => \N__41376\,
            I => \N__41373\
        );

    \I__8918\ : CascadeBuf
    port map (
            O => \N__41373\,
            I => \N__41370\
        );

    \I__8917\ : CascadeMux
    port map (
            O => \N__41370\,
            I => \N__41366\
        );

    \I__8916\ : CascadeMux
    port map (
            O => \N__41369\,
            I => \N__41363\
        );

    \I__8915\ : CascadeBuf
    port map (
            O => \N__41366\,
            I => \N__41360\
        );

    \I__8914\ : CascadeBuf
    port map (
            O => \N__41363\,
            I => \N__41357\
        );

    \I__8913\ : CascadeMux
    port map (
            O => \N__41360\,
            I => \N__41354\
        );

    \I__8912\ : CascadeMux
    port map (
            O => \N__41357\,
            I => \N__41351\
        );

    \I__8911\ : CascadeBuf
    port map (
            O => \N__41354\,
            I => \N__41348\
        );

    \I__8910\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41345\
        );

    \I__8909\ : CascadeMux
    port map (
            O => \N__41348\,
            I => \N__41342\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__41345\,
            I => \N__41339\
        );

    \I__8907\ : CascadeBuf
    port map (
            O => \N__41342\,
            I => \N__41336\
        );

    \I__8906\ : Span4Mux_h
    port map (
            O => \N__41339\,
            I => \N__41333\
        );

    \I__8905\ : CascadeMux
    port map (
            O => \N__41336\,
            I => \N__41330\
        );

    \I__8904\ : Span4Mux_v
    port map (
            O => \N__41333\,
            I => \N__41327\
        );

    \I__8903\ : InMux
    port map (
            O => \N__41330\,
            I => \N__41324\
        );

    \I__8902\ : Span4Mux_v
    port map (
            O => \N__41327\,
            I => \N__41321\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__41324\,
            I => \N__41318\
        );

    \I__8900\ : Span4Mux_h
    port map (
            O => \N__41321\,
            I => \N__41315\
        );

    \I__8899\ : Span4Mux_h
    port map (
            O => \N__41318\,
            I => \N__41312\
        );

    \I__8898\ : Span4Mux_h
    port map (
            O => \N__41315\,
            I => \N__41307\
        );

    \I__8897\ : Span4Mux_h
    port map (
            O => \N__41312\,
            I => \N__41307\
        );

    \I__8896\ : Odrv4
    port map (
            O => \N__41307\,
            I => \data_index_9_N_212_5\
        );

    \I__8895\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41300\
        );

    \I__8894\ : InMux
    port map (
            O => \N__41303\,
            I => \N__41297\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41300\,
            I => \N__41293\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__41297\,
            I => \N__41290\
        );

    \I__8891\ : CascadeMux
    port map (
            O => \N__41296\,
            I => \N__41287\
        );

    \I__8890\ : Span4Mux_h
    port map (
            O => \N__41293\,
            I => \N__41284\
        );

    \I__8889\ : Span12Mux_s11_v
    port map (
            O => \N__41290\,
            I => \N__41281\
        );

    \I__8888\ : InMux
    port map (
            O => \N__41287\,
            I => \N__41278\
        );

    \I__8887\ : Span4Mux_h
    port map (
            O => \N__41284\,
            I => \N__41275\
        );

    \I__8886\ : Span12Mux_h
    port map (
            O => \N__41281\,
            I => \N__41272\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__41278\,
            I => buf_adcdata_iac_11
        );

    \I__8884\ : Odrv4
    port map (
            O => \N__41275\,
            I => buf_adcdata_iac_11
        );

    \I__8883\ : Odrv12
    port map (
            O => \N__41272\,
            I => buf_adcdata_iac_11
        );

    \I__8882\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41262\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__41262\,
            I => \N__41259\
        );

    \I__8880\ : Odrv12
    port map (
            O => \N__41259\,
            I => n16_adj_1640
        );

    \I__8879\ : CascadeMux
    port map (
            O => \N__41256\,
            I => \n22623_cascade_\
        );

    \I__8878\ : CascadeMux
    port map (
            O => \N__41253\,
            I => \n22626_cascade_\
        );

    \I__8877\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41247\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__41247\,
            I => n30_adj_1643
        );

    \I__8875\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41241\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__41241\,
            I => \N__41238\
        );

    \I__8873\ : Span4Mux_h
    port map (
            O => \N__41238\,
            I => \N__41234\
        );

    \I__8872\ : InMux
    port map (
            O => \N__41237\,
            I => \N__41231\
        );

    \I__8871\ : Span4Mux_h
    port map (
            O => \N__41234\,
            I => \N__41228\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__41231\,
            I => data_idxvec_3
        );

    \I__8869\ : Odrv4
    port map (
            O => \N__41228\,
            I => data_idxvec_3
        );

    \I__8868\ : InMux
    port map (
            O => \N__41223\,
            I => \N__41220\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__41220\,
            I => \N__41216\
        );

    \I__8866\ : InMux
    port map (
            O => \N__41219\,
            I => \N__41212\
        );

    \I__8865\ : Span4Mux_v
    port map (
            O => \N__41216\,
            I => \N__41209\
        );

    \I__8864\ : InMux
    port map (
            O => \N__41215\,
            I => \N__41206\
        );

    \I__8863\ : LocalMux
    port map (
            O => \N__41212\,
            I => data_cntvec_3
        );

    \I__8862\ : Odrv4
    port map (
            O => \N__41209\,
            I => data_cntvec_3
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__41206\,
            I => data_cntvec_3
        );

    \I__8860\ : CascadeMux
    port map (
            O => \N__41199\,
            I => \n26_adj_1642_cascade_\
        );

    \I__8859\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41193\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__41193\,
            I => \N__41189\
        );

    \I__8857\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41185\
        );

    \I__8856\ : Span4Mux_v
    port map (
            O => \N__41189\,
            I => \N__41182\
        );

    \I__8855\ : InMux
    port map (
            O => \N__41188\,
            I => \N__41179\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__41185\,
            I => req_data_cnt_3
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__41182\,
            I => req_data_cnt_3
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__41179\,
            I => req_data_cnt_3
        );

    \I__8851\ : CascadeMux
    port map (
            O => \N__41172\,
            I => \n22425_cascade_\
        );

    \I__8850\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41166\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__41166\,
            I => \N__41163\
        );

    \I__8848\ : Span4Mux_h
    port map (
            O => \N__41163\,
            I => \N__41158\
        );

    \I__8847\ : InMux
    port map (
            O => \N__41162\,
            I => \N__41153\
        );

    \I__8846\ : InMux
    port map (
            O => \N__41161\,
            I => \N__41153\
        );

    \I__8845\ : Odrv4
    port map (
            O => \N__41158\,
            I => \acadc_skipCount_3\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__41153\,
            I => \acadc_skipCount_3\
        );

    \I__8843\ : InMux
    port map (
            O => \N__41148\,
            I => \N__41145\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__41145\,
            I => n22428
        );

    \I__8841\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41137\
        );

    \I__8840\ : InMux
    port map (
            O => \N__41141\,
            I => \N__41134\
        );

    \I__8839\ : InMux
    port map (
            O => \N__41140\,
            I => \N__41131\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__41137\,
            I => data_index_0
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__41134\,
            I => data_index_0
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__41131\,
            I => data_index_0
        );

    \I__8835\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41116\
        );

    \I__8834\ : InMux
    port map (
            O => \N__41123\,
            I => \N__41113\
        );

    \I__8833\ : InMux
    port map (
            O => \N__41122\,
            I => \N__41108\
        );

    \I__8832\ : InMux
    port map (
            O => \N__41121\,
            I => \N__41108\
        );

    \I__8831\ : InMux
    port map (
            O => \N__41120\,
            I => \N__41103\
        );

    \I__8830\ : InMux
    port map (
            O => \N__41119\,
            I => \N__41103\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__41116\,
            I => \N__41097\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__41113\,
            I => \N__41093\
        );

    \I__8827\ : LocalMux
    port map (
            O => \N__41108\,
            I => \N__41088\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__41103\,
            I => \N__41088\
        );

    \I__8825\ : InMux
    port map (
            O => \N__41102\,
            I => \N__41085\
        );

    \I__8824\ : InMux
    port map (
            O => \N__41101\,
            I => \N__41080\
        );

    \I__8823\ : InMux
    port map (
            O => \N__41100\,
            I => \N__41080\
        );

    \I__8822\ : Span4Mux_v
    port map (
            O => \N__41097\,
            I => \N__41076\
        );

    \I__8821\ : InMux
    port map (
            O => \N__41096\,
            I => \N__41073\
        );

    \I__8820\ : Span4Mux_v
    port map (
            O => \N__41093\,
            I => \N__41064\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__41088\,
            I => \N__41064\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__41085\,
            I => \N__41064\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__41080\,
            I => \N__41064\
        );

    \I__8816\ : InMux
    port map (
            O => \N__41079\,
            I => \N__41061\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__41076\,
            I => n8841
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__41073\,
            I => n8841
        );

    \I__8813\ : Odrv4
    port map (
            O => \N__41064\,
            I => n8841
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__41061\,
            I => n8841
        );

    \I__8811\ : InMux
    port map (
            O => \N__41052\,
            I => \N__41049\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__41049\,
            I => n8_adj_1540
        );

    \I__8809\ : InMux
    port map (
            O => \N__41046\,
            I => \N__41040\
        );

    \I__8808\ : InMux
    port map (
            O => \N__41045\,
            I => \N__41040\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__41040\,
            I => n7_adj_1539
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__41037\,
            I => \n8_adj_1540_cascade_\
        );

    \I__8805\ : CascadeMux
    port map (
            O => \N__41034\,
            I => \N__41031\
        );

    \I__8804\ : CascadeBuf
    port map (
            O => \N__41031\,
            I => \N__41028\
        );

    \I__8803\ : CascadeMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__8802\ : CascadeBuf
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__8801\ : CascadeMux
    port map (
            O => \N__41022\,
            I => \N__41019\
        );

    \I__8800\ : CascadeBuf
    port map (
            O => \N__41019\,
            I => \N__41016\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__41016\,
            I => \N__41013\
        );

    \I__8798\ : CascadeBuf
    port map (
            O => \N__41013\,
            I => \N__41010\
        );

    \I__8797\ : CascadeMux
    port map (
            O => \N__41010\,
            I => \N__41007\
        );

    \I__8796\ : CascadeBuf
    port map (
            O => \N__41007\,
            I => \N__41004\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__41004\,
            I => \N__41001\
        );

    \I__8794\ : CascadeBuf
    port map (
            O => \N__41001\,
            I => \N__40998\
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__40998\,
            I => \N__40995\
        );

    \I__8792\ : CascadeBuf
    port map (
            O => \N__40995\,
            I => \N__40991\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__40994\,
            I => \N__40988\
        );

    \I__8790\ : CascadeMux
    port map (
            O => \N__40991\,
            I => \N__40985\
        );

    \I__8789\ : CascadeBuf
    port map (
            O => \N__40988\,
            I => \N__40982\
        );

    \I__8788\ : CascadeBuf
    port map (
            O => \N__40985\,
            I => \N__40979\
        );

    \I__8787\ : CascadeMux
    port map (
            O => \N__40982\,
            I => \N__40976\
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__40979\,
            I => \N__40973\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40976\,
            I => \N__40970\
        );

    \I__8784\ : CascadeBuf
    port map (
            O => \N__40973\,
            I => \N__40967\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__40970\,
            I => \N__40964\
        );

    \I__8782\ : CascadeMux
    port map (
            O => \N__40967\,
            I => \N__40961\
        );

    \I__8781\ : Span4Mux_h
    port map (
            O => \N__40964\,
            I => \N__40958\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40955\
        );

    \I__8779\ : Span4Mux_v
    port map (
            O => \N__40958\,
            I => \N__40952\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40955\,
            I => \N__40949\
        );

    \I__8777\ : Span4Mux_h
    port map (
            O => \N__40952\,
            I => \N__40946\
        );

    \I__8776\ : Span4Mux_h
    port map (
            O => \N__40949\,
            I => \N__40943\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__40946\,
            I => \N__40940\
        );

    \I__8774\ : Span4Mux_v
    port map (
            O => \N__40943\,
            I => \N__40937\
        );

    \I__8773\ : Odrv4
    port map (
            O => \N__40940\,
            I => \data_index_9_N_212_0\
        );

    \I__8772\ : Odrv4
    port map (
            O => \N__40937\,
            I => \data_index_9_N_212_0\
        );

    \I__8771\ : CascadeMux
    port map (
            O => \N__40932\,
            I => \n30_adj_1688_cascade_\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40926\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40926\,
            I => \N__40922\
        );

    \I__8768\ : CascadeMux
    port map (
            O => \N__40925\,
            I => \N__40919\
        );

    \I__8767\ : Span4Mux_h
    port map (
            O => \N__40922\,
            I => \N__40916\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40919\,
            I => \N__40913\
        );

    \I__8765\ : Span4Mux_h
    port map (
            O => \N__40916\,
            I => \N__40910\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40913\,
            I => data_idxvec_8
        );

    \I__8763\ : Odrv4
    port map (
            O => \N__40910\,
            I => data_idxvec_8
        );

    \I__8762\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40902\,
            I => \N__40898\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40901\,
            I => \N__40894\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__40898\,
            I => \N__40891\
        );

    \I__8758\ : InMux
    port map (
            O => \N__40897\,
            I => \N__40888\
        );

    \I__8757\ : LocalMux
    port map (
            O => \N__40894\,
            I => data_cntvec_8
        );

    \I__8756\ : Odrv4
    port map (
            O => \N__40891\,
            I => data_cntvec_8
        );

    \I__8755\ : LocalMux
    port map (
            O => \N__40888\,
            I => data_cntvec_8
        );

    \I__8754\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40878\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__40878\,
            I => \N__40875\
        );

    \I__8752\ : Span4Mux_h
    port map (
            O => \N__40875\,
            I => \N__40872\
        );

    \I__8751\ : Span4Mux_h
    port map (
            O => \N__40872\,
            I => \N__40869\
        );

    \I__8750\ : Odrv4
    port map (
            O => \N__40869\,
            I => buf_data_iac_16
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__40866\,
            I => \n26_adj_1533_cascade_\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40863\,
            I => \N__40860\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__40860\,
            I => \N__40857\
        );

    \I__8746\ : Odrv12
    port map (
            O => \N__40857\,
            I => n22398
        );

    \I__8745\ : CascadeMux
    port map (
            O => \N__40854\,
            I => \n21246_cascade_\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40848\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__40848\,
            I => \N__40845\
        );

    \I__8742\ : Span4Mux_h
    port map (
            O => \N__40845\,
            I => \N__40842\
        );

    \I__8741\ : Odrv4
    port map (
            O => \N__40842\,
            I => n22392
        );

    \I__8740\ : InMux
    port map (
            O => \N__40839\,
            I => \N__40836\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__40836\,
            I => \N__40833\
        );

    \I__8738\ : Span4Mux_v
    port map (
            O => \N__40833\,
            I => \N__40830\
        );

    \I__8737\ : Span4Mux_h
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__40827\,
            I => n22578
        );

    \I__8735\ : CascadeMux
    port map (
            O => \N__40824\,
            I => \n22581_cascade_\
        );

    \I__8734\ : CascadeMux
    port map (
            O => \N__40821\,
            I => \n22584_cascade_\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40818\,
            I => \N__40815\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40815\,
            I => \N__40812\
        );

    \I__8731\ : Span4Mux_h
    port map (
            O => \N__40812\,
            I => \N__40809\
        );

    \I__8730\ : Span4Mux_h
    port map (
            O => \N__40809\,
            I => \N__40806\
        );

    \I__8729\ : Span4Mux_h
    port map (
            O => \N__40806\,
            I => \N__40802\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40805\,
            I => \N__40799\
        );

    \I__8727\ : Odrv4
    port map (
            O => \N__40802\,
            I => \buf_readRTD_3\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40799\,
            I => \buf_readRTD_3\
        );

    \I__8725\ : CascadeMux
    port map (
            O => \N__40794\,
            I => \N__40791\
        );

    \I__8724\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40788\,
            I => \N__40785\
        );

    \I__8722\ : Span4Mux_v
    port map (
            O => \N__40785\,
            I => \N__40782\
        );

    \I__8721\ : Odrv4
    port map (
            O => \N__40782\,
            I => n19_adj_1641
        );

    \I__8720\ : CascadeMux
    port map (
            O => \N__40779\,
            I => \n21556_cascade_\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40776\,
            I => \N__40773\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__8717\ : Span4Mux_v
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__8716\ : Odrv4
    port map (
            O => \N__40767\,
            I => n21703
        );

    \I__8715\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40761\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__40761\,
            I => n22521
        );

    \I__8713\ : InMux
    port map (
            O => \N__40758\,
            I => \N__40755\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__40755\,
            I => n22464
        );

    \I__8711\ : CascadeMux
    port map (
            O => \N__40752\,
            I => \n22524_cascade_\
        );

    \I__8710\ : CascadeMux
    port map (
            O => \N__40749\,
            I => \n30_adj_1676_cascade_\
        );

    \I__8709\ : InMux
    port map (
            O => \N__40746\,
            I => \N__40743\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__40743\,
            I => \N__40740\
        );

    \I__8707\ : Span4Mux_h
    port map (
            O => \N__40740\,
            I => \N__40737\
        );

    \I__8706\ : Span4Mux_h
    port map (
            O => \N__40737\,
            I => \N__40734\
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__40734\,
            I => n17_adj_1682
        );

    \I__8704\ : CascadeMux
    port map (
            O => \N__40731\,
            I => \N__40728\
        );

    \I__8703\ : InMux
    port map (
            O => \N__40728\,
            I => \N__40725\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40725\,
            I => \N__40722\
        );

    \I__8701\ : Span4Mux_v
    port map (
            O => \N__40722\,
            I => \N__40719\
        );

    \I__8700\ : Odrv4
    port map (
            O => \N__40719\,
            I => n16_adj_1681
        );

    \I__8699\ : InMux
    port map (
            O => \N__40716\,
            I => \N__40713\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40713\,
            I => \N__40710\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__40710\,
            I => \N__40707\
        );

    \I__8696\ : Odrv4
    port map (
            O => \N__40707\,
            I => n22485
        );

    \I__8695\ : InMux
    port map (
            O => \N__40704\,
            I => \N__40700\
        );

    \I__8694\ : CascadeMux
    port map (
            O => \N__40703\,
            I => \N__40697\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__40700\,
            I => \N__40694\
        );

    \I__8692\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40691\
        );

    \I__8691\ : Span12Mux_v
    port map (
            O => \N__40694\,
            I => \N__40688\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__40691\,
            I => data_idxvec_10
        );

    \I__8689\ : Odrv12
    port map (
            O => \N__40688\,
            I => data_idxvec_10
        );

    \I__8688\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40679\
        );

    \I__8687\ : InMux
    port map (
            O => \N__40682\,
            I => \N__40675\
        );

    \I__8686\ : LocalMux
    port map (
            O => \N__40679\,
            I => \N__40672\
        );

    \I__8685\ : InMux
    port map (
            O => \N__40678\,
            I => \N__40669\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__40675\,
            I => \N__40666\
        );

    \I__8683\ : Span4Mux_v
    port map (
            O => \N__40672\,
            I => \N__40663\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40669\,
            I => data_cntvec_10
        );

    \I__8681\ : Odrv4
    port map (
            O => \N__40666\,
            I => data_cntvec_10
        );

    \I__8680\ : Odrv4
    port map (
            O => \N__40663\,
            I => data_cntvec_10
        );

    \I__8679\ : CascadeMux
    port map (
            O => \N__40656\,
            I => \n26_adj_1687_cascade_\
        );

    \I__8678\ : CascadeMux
    port map (
            O => \N__40653\,
            I => \n22455_cascade_\
        );

    \I__8677\ : InMux
    port map (
            O => \N__40650\,
            I => \N__40647\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__40647\,
            I => \N__40644\
        );

    \I__8675\ : Span4Mux_v
    port map (
            O => \N__40644\,
            I => \N__40641\
        );

    \I__8674\ : Span4Mux_h
    port map (
            O => \N__40641\,
            I => \N__40638\
        );

    \I__8673\ : Sp12to4
    port map (
            O => \N__40638\,
            I => \N__40635\
        );

    \I__8672\ : Odrv12
    port map (
            O => \N__40635\,
            I => n24_adj_1686
        );

    \I__8671\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40629\
        );

    \I__8670\ : LocalMux
    port map (
            O => \N__40629\,
            I => n22488
        );

    \I__8669\ : CascadeMux
    port map (
            O => \N__40626\,
            I => \n22458_cascade_\
        );

    \I__8668\ : ClkMux
    port map (
            O => \N__40623\,
            I => \N__40618\
        );

    \I__8667\ : ClkMux
    port map (
            O => \N__40622\,
            I => \N__40604\
        );

    \I__8666\ : ClkMux
    port map (
            O => \N__40621\,
            I => \N__40601\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__40618\,
            I => \N__40598\
        );

    \I__8664\ : ClkMux
    port map (
            O => \N__40617\,
            I => \N__40595\
        );

    \I__8663\ : ClkMux
    port map (
            O => \N__40616\,
            I => \N__40592\
        );

    \I__8662\ : ClkMux
    port map (
            O => \N__40615\,
            I => \N__40589\
        );

    \I__8661\ : ClkMux
    port map (
            O => \N__40614\,
            I => \N__40586\
        );

    \I__8660\ : ClkMux
    port map (
            O => \N__40613\,
            I => \N__40583\
        );

    \I__8659\ : ClkMux
    port map (
            O => \N__40612\,
            I => \N__40579\
        );

    \I__8658\ : ClkMux
    port map (
            O => \N__40611\,
            I => \N__40576\
        );

    \I__8657\ : ClkMux
    port map (
            O => \N__40610\,
            I => \N__40573\
        );

    \I__8656\ : ClkMux
    port map (
            O => \N__40609\,
            I => \N__40570\
        );

    \I__8655\ : ClkMux
    port map (
            O => \N__40608\,
            I => \N__40566\
        );

    \I__8654\ : ClkMux
    port map (
            O => \N__40607\,
            I => \N__40563\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__40604\,
            I => \N__40558\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__40601\,
            I => \N__40558\
        );

    \I__8651\ : Span4Mux_v
    port map (
            O => \N__40598\,
            I => \N__40555\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__40595\,
            I => \N__40550\
        );

    \I__8649\ : LocalMux
    port map (
            O => \N__40592\,
            I => \N__40550\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__40589\,
            I => \N__40547\
        );

    \I__8647\ : LocalMux
    port map (
            O => \N__40586\,
            I => \N__40542\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__40583\,
            I => \N__40542\
        );

    \I__8645\ : ClkMux
    port map (
            O => \N__40582\,
            I => \N__40539\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40579\,
            I => \N__40535\
        );

    \I__8643\ : LocalMux
    port map (
            O => \N__40576\,
            I => \N__40530\
        );

    \I__8642\ : LocalMux
    port map (
            O => \N__40573\,
            I => \N__40530\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__40570\,
            I => \N__40527\
        );

    \I__8640\ : ClkMux
    port map (
            O => \N__40569\,
            I => \N__40524\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__40566\,
            I => \N__40519\
        );

    \I__8638\ : LocalMux
    port map (
            O => \N__40563\,
            I => \N__40519\
        );

    \I__8637\ : Span4Mux_v
    port map (
            O => \N__40558\,
            I => \N__40516\
        );

    \I__8636\ : Span4Mux_v
    port map (
            O => \N__40555\,
            I => \N__40505\
        );

    \I__8635\ : Span4Mux_v
    port map (
            O => \N__40550\,
            I => \N__40505\
        );

    \I__8634\ : Span4Mux_h
    port map (
            O => \N__40547\,
            I => \N__40505\
        );

    \I__8633\ : Span4Mux_v
    port map (
            O => \N__40542\,
            I => \N__40505\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__40539\,
            I => \N__40505\
        );

    \I__8631\ : ClkMux
    port map (
            O => \N__40538\,
            I => \N__40502\
        );

    \I__8630\ : Span4Mux_v
    port map (
            O => \N__40535\,
            I => \N__40497\
        );

    \I__8629\ : Span4Mux_v
    port map (
            O => \N__40530\,
            I => \N__40497\
        );

    \I__8628\ : Span4Mux_v
    port map (
            O => \N__40527\,
            I => \N__40492\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__40524\,
            I => \N__40492\
        );

    \I__8626\ : Span4Mux_v
    port map (
            O => \N__40519\,
            I => \N__40485\
        );

    \I__8625\ : Span4Mux_h
    port map (
            O => \N__40516\,
            I => \N__40485\
        );

    \I__8624\ : Span4Mux_h
    port map (
            O => \N__40505\,
            I => \N__40485\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40502\,
            I => \N__40482\
        );

    \I__8622\ : Span4Mux_h
    port map (
            O => \N__40497\,
            I => \N__40477\
        );

    \I__8621\ : Span4Mux_h
    port map (
            O => \N__40492\,
            I => \N__40477\
        );

    \I__8620\ : Span4Mux_h
    port map (
            O => \N__40485\,
            I => \N__40474\
        );

    \I__8619\ : Span12Mux_h
    port map (
            O => \N__40482\,
            I => \N__40470\
        );

    \I__8618\ : Span4Mux_h
    port map (
            O => \N__40477\,
            I => \N__40467\
        );

    \I__8617\ : Span4Mux_h
    port map (
            O => \N__40474\,
            I => \N__40464\
        );

    \I__8616\ : InMux
    port map (
            O => \N__40473\,
            I => \N__40461\
        );

    \I__8615\ : Odrv12
    port map (
            O => \N__40470\,
            I => \clk_RTD\
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__40467\,
            I => \clk_RTD\
        );

    \I__8613\ : Odrv4
    port map (
            O => \N__40464\,
            I => \clk_RTD\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__40461\,
            I => \clk_RTD\
        );

    \I__8611\ : InMux
    port map (
            O => \N__40452\,
            I => \N__40449\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__40449\,
            I => \N__40444\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40448\,
            I => \N__40441\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40447\,
            I => \N__40438\
        );

    \I__8607\ : Span4Mux_h
    port map (
            O => \N__40444\,
            I => \N__40435\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__40441\,
            I => \N__40430\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40430\
        );

    \I__8604\ : Span4Mux_h
    port map (
            O => \N__40435\,
            I => \N__40427\
        );

    \I__8603\ : Odrv12
    port map (
            O => \N__40430\,
            I => n14_adj_1550
        );

    \I__8602\ : Odrv4
    port map (
            O => \N__40427\,
            I => n14_adj_1550
        );

    \I__8601\ : InMux
    port map (
            O => \N__40422\,
            I => \N__40419\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__40419\,
            I => \N__40416\
        );

    \I__8599\ : Odrv12
    port map (
            O => \N__40416\,
            I => n17_adj_1672
        );

    \I__8598\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40410\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__40410\,
            I => \N__40407\
        );

    \I__8596\ : Span4Mux_h
    port map (
            O => \N__40407\,
            I => \N__40404\
        );

    \I__8595\ : Odrv4
    port map (
            O => \N__40404\,
            I => n22461
        );

    \I__8594\ : CascadeMux
    port map (
            O => \N__40401\,
            I => \N__40398\
        );

    \I__8593\ : InMux
    port map (
            O => \N__40398\,
            I => \N__40395\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__40395\,
            I => \N__40392\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__40392\,
            I => \N__40389\
        );

    \I__8590\ : Span4Mux_v
    port map (
            O => \N__40389\,
            I => \N__40386\
        );

    \I__8589\ : Odrv4
    port map (
            O => \N__40386\,
            I => n16_adj_1671
        );

    \I__8588\ : InMux
    port map (
            O => \N__40383\,
            I => \N__40380\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__40380\,
            I => \N__40376\
        );

    \I__8586\ : CascadeMux
    port map (
            O => \N__40379\,
            I => \N__40373\
        );

    \I__8585\ : Span4Mux_h
    port map (
            O => \N__40376\,
            I => \N__40370\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40367\
        );

    \I__8583\ : Span4Mux_h
    port map (
            O => \N__40370\,
            I => \N__40364\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__40367\,
            I => data_idxvec_12
        );

    \I__8581\ : Odrv4
    port map (
            O => \N__40364\,
            I => data_idxvec_12
        );

    \I__8580\ : InMux
    port map (
            O => \N__40359\,
            I => \N__40355\
        );

    \I__8579\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40352\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__40355\,
            I => wdtick_cnt_22
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__40352\,
            I => wdtick_cnt_22
        );

    \I__8576\ : InMux
    port map (
            O => \N__40347\,
            I => n19953
        );

    \I__8575\ : InMux
    port map (
            O => \N__40344\,
            I => \N__40340\
        );

    \I__8574\ : InMux
    port map (
            O => \N__40343\,
            I => \N__40337\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__40340\,
            I => wdtick_cnt_23
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__40337\,
            I => wdtick_cnt_23
        );

    \I__8571\ : InMux
    port map (
            O => \N__40332\,
            I => n19954
        );

    \I__8570\ : InMux
    port map (
            O => \N__40329\,
            I => \N__40296\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40328\,
            I => \N__40296\
        );

    \I__8568\ : InMux
    port map (
            O => \N__40327\,
            I => \N__40296\
        );

    \I__8567\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40296\
        );

    \I__8566\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40293\
        );

    \I__8565\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40284\
        );

    \I__8564\ : InMux
    port map (
            O => \N__40323\,
            I => \N__40284\
        );

    \I__8563\ : InMux
    port map (
            O => \N__40322\,
            I => \N__40284\
        );

    \I__8562\ : InMux
    port map (
            O => \N__40321\,
            I => \N__40284\
        );

    \I__8561\ : InMux
    port map (
            O => \N__40320\,
            I => \N__40275\
        );

    \I__8560\ : InMux
    port map (
            O => \N__40319\,
            I => \N__40275\
        );

    \I__8559\ : InMux
    port map (
            O => \N__40318\,
            I => \N__40275\
        );

    \I__8558\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40275\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40316\,
            I => \N__40266\
        );

    \I__8556\ : InMux
    port map (
            O => \N__40315\,
            I => \N__40266\
        );

    \I__8555\ : InMux
    port map (
            O => \N__40314\,
            I => \N__40266\
        );

    \I__8554\ : InMux
    port map (
            O => \N__40313\,
            I => \N__40266\
        );

    \I__8553\ : InMux
    port map (
            O => \N__40312\,
            I => \N__40257\
        );

    \I__8552\ : InMux
    port map (
            O => \N__40311\,
            I => \N__40257\
        );

    \I__8551\ : InMux
    port map (
            O => \N__40310\,
            I => \N__40257\
        );

    \I__8550\ : InMux
    port map (
            O => \N__40309\,
            I => \N__40257\
        );

    \I__8549\ : InMux
    port map (
            O => \N__40308\,
            I => \N__40248\
        );

    \I__8548\ : InMux
    port map (
            O => \N__40307\,
            I => \N__40248\
        );

    \I__8547\ : InMux
    port map (
            O => \N__40306\,
            I => \N__40248\
        );

    \I__8546\ : InMux
    port map (
            O => \N__40305\,
            I => \N__40248\
        );

    \I__8545\ : LocalMux
    port map (
            O => \N__40296\,
            I => \N__40243\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__40293\,
            I => \N__40243\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__40284\,
            I => n49
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__40275\,
            I => n49
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__40266\,
            I => n49
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__40257\,
            I => n49
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__40248\,
            I => n49
        );

    \I__8538\ : Odrv4
    port map (
            O => \N__40243\,
            I => n49
        );

    \I__8537\ : InMux
    port map (
            O => \N__40230\,
            I => \bfn_15_8_0_\
        );

    \I__8536\ : InMux
    port map (
            O => \N__40227\,
            I => \N__40223\
        );

    \I__8535\ : InMux
    port map (
            O => \N__40226\,
            I => \N__40220\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__40223\,
            I => \N__40217\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__40220\,
            I => wdtick_cnt_24
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__40217\,
            I => wdtick_cnt_24
        );

    \I__8531\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40208\
        );

    \I__8530\ : InMux
    port map (
            O => \N__40211\,
            I => \N__40205\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__40208\,
            I => \N__40200\
        );

    \I__8528\ : LocalMux
    port map (
            O => \N__40205\,
            I => \N__40200\
        );

    \I__8527\ : Odrv4
    port map (
            O => \N__40200\,
            I => wdtick_cnt_14
        );

    \I__8526\ : InMux
    port map (
            O => \N__40197\,
            I => n19945
        );

    \I__8525\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40190\
        );

    \I__8524\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40187\
        );

    \I__8523\ : LocalMux
    port map (
            O => \N__40190\,
            I => wdtick_cnt_15
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__40187\,
            I => wdtick_cnt_15
        );

    \I__8521\ : InMux
    port map (
            O => \N__40182\,
            I => n19946
        );

    \I__8520\ : InMux
    port map (
            O => \N__40179\,
            I => \N__40175\
        );

    \I__8519\ : InMux
    port map (
            O => \N__40178\,
            I => \N__40172\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__40175\,
            I => wdtick_cnt_16
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__40172\,
            I => wdtick_cnt_16
        );

    \I__8516\ : InMux
    port map (
            O => \N__40167\,
            I => \bfn_15_7_0_\
        );

    \I__8515\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40160\
        );

    \I__8514\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40157\
        );

    \I__8513\ : LocalMux
    port map (
            O => \N__40160\,
            I => wdtick_cnt_17
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__40157\,
            I => wdtick_cnt_17
        );

    \I__8511\ : InMux
    port map (
            O => \N__40152\,
            I => n19948
        );

    \I__8510\ : CascadeMux
    port map (
            O => \N__40149\,
            I => \N__40145\
        );

    \I__8509\ : InMux
    port map (
            O => \N__40148\,
            I => \N__40142\
        );

    \I__8508\ : InMux
    port map (
            O => \N__40145\,
            I => \N__40139\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__40142\,
            I => wdtick_cnt_18
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__40139\,
            I => wdtick_cnt_18
        );

    \I__8505\ : InMux
    port map (
            O => \N__40134\,
            I => n19949
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__40131\,
            I => \N__40127\
        );

    \I__8503\ : InMux
    port map (
            O => \N__40130\,
            I => \N__40124\
        );

    \I__8502\ : InMux
    port map (
            O => \N__40127\,
            I => \N__40121\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__40124\,
            I => wdtick_cnt_19
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__40121\,
            I => wdtick_cnt_19
        );

    \I__8499\ : InMux
    port map (
            O => \N__40116\,
            I => n19950
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__40113\,
            I => \N__40109\
        );

    \I__8497\ : InMux
    port map (
            O => \N__40112\,
            I => \N__40106\
        );

    \I__8496\ : InMux
    port map (
            O => \N__40109\,
            I => \N__40103\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__40106\,
            I => wdtick_cnt_20
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__40103\,
            I => wdtick_cnt_20
        );

    \I__8493\ : InMux
    port map (
            O => \N__40098\,
            I => n19951
        );

    \I__8492\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40091\
        );

    \I__8491\ : InMux
    port map (
            O => \N__40094\,
            I => \N__40088\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__40091\,
            I => wdtick_cnt_21
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__40088\,
            I => wdtick_cnt_21
        );

    \I__8488\ : InMux
    port map (
            O => \N__40083\,
            I => n19952
        );

    \I__8487\ : CascadeMux
    port map (
            O => \N__40080\,
            I => \N__40077\
        );

    \I__8486\ : InMux
    port map (
            O => \N__40077\,
            I => \N__40074\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__40074\,
            I => \N__40070\
        );

    \I__8484\ : InMux
    port map (
            O => \N__40073\,
            I => \N__40067\
        );

    \I__8483\ : Span4Mux_h
    port map (
            O => \N__40070\,
            I => \N__40064\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__40067\,
            I => wdtick_cnt_6
        );

    \I__8481\ : Odrv4
    port map (
            O => \N__40064\,
            I => wdtick_cnt_6
        );

    \I__8480\ : InMux
    port map (
            O => \N__40059\,
            I => n19937
        );

    \I__8479\ : InMux
    port map (
            O => \N__40056\,
            I => \N__40052\
        );

    \I__8478\ : InMux
    port map (
            O => \N__40055\,
            I => \N__40049\
        );

    \I__8477\ : LocalMux
    port map (
            O => \N__40052\,
            I => \N__40046\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__40049\,
            I => wdtick_cnt_7
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__40046\,
            I => wdtick_cnt_7
        );

    \I__8474\ : InMux
    port map (
            O => \N__40041\,
            I => n19938
        );

    \I__8473\ : CascadeMux
    port map (
            O => \N__40038\,
            I => \N__40035\
        );

    \I__8472\ : InMux
    port map (
            O => \N__40035\,
            I => \N__40031\
        );

    \I__8471\ : InMux
    port map (
            O => \N__40034\,
            I => \N__40028\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__40031\,
            I => \N__40025\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__40028\,
            I => wdtick_cnt_8
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__40025\,
            I => wdtick_cnt_8
        );

    \I__8467\ : InMux
    port map (
            O => \N__40020\,
            I => \bfn_15_6_0_\
        );

    \I__8466\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40013\
        );

    \I__8465\ : InMux
    port map (
            O => \N__40016\,
            I => \N__40010\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__40013\,
            I => wdtick_cnt_9
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__40010\,
            I => wdtick_cnt_9
        );

    \I__8462\ : InMux
    port map (
            O => \N__40005\,
            I => n19940
        );

    \I__8461\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39999\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__39999\,
            I => \N__39995\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39998\,
            I => \N__39992\
        );

    \I__8458\ : Span4Mux_h
    port map (
            O => \N__39995\,
            I => \N__39989\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__39992\,
            I => wdtick_cnt_10
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__39989\,
            I => wdtick_cnt_10
        );

    \I__8455\ : InMux
    port map (
            O => \N__39984\,
            I => n19941
        );

    \I__8454\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39977\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39974\
        );

    \I__8452\ : LocalMux
    port map (
            O => \N__39977\,
            I => wdtick_cnt_11
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39974\,
            I => wdtick_cnt_11
        );

    \I__8450\ : InMux
    port map (
            O => \N__39969\,
            I => n19942
        );

    \I__8449\ : InMux
    port map (
            O => \N__39966\,
            I => \N__39963\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39963\,
            I => \N__39959\
        );

    \I__8447\ : InMux
    port map (
            O => \N__39962\,
            I => \N__39956\
        );

    \I__8446\ : Span4Mux_v
    port map (
            O => \N__39959\,
            I => \N__39953\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39956\,
            I => wdtick_cnt_12
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__39953\,
            I => wdtick_cnt_12
        );

    \I__8443\ : InMux
    port map (
            O => \N__39948\,
            I => n19943
        );

    \I__8442\ : InMux
    port map (
            O => \N__39945\,
            I => \N__39941\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39944\,
            I => \N__39938\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__39941\,
            I => wdtick_cnt_13
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__39938\,
            I => wdtick_cnt_13
        );

    \I__8438\ : InMux
    port map (
            O => \N__39933\,
            I => n19944
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__39930\,
            I => \N__39926\
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__39929\,
            I => \N__39923\
        );

    \I__8435\ : InMux
    port map (
            O => \N__39926\,
            I => \N__39918\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39923\,
            I => \N__39918\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__39918\,
            I => n8_adj_1568
        );

    \I__8432\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39909\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39914\,
            I => \N__39909\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39909\,
            I => \N__39906\
        );

    \I__8429\ : Odrv12
    port map (
            O => \N__39906\,
            I => n7_adj_1567
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__39903\,
            I => \N__39900\
        );

    \I__8427\ : CascadeBuf
    port map (
            O => \N__39900\,
            I => \N__39897\
        );

    \I__8426\ : CascadeMux
    port map (
            O => \N__39897\,
            I => \N__39894\
        );

    \I__8425\ : CascadeBuf
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__39891\,
            I => \N__39888\
        );

    \I__8423\ : CascadeBuf
    port map (
            O => \N__39888\,
            I => \N__39885\
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__8421\ : CascadeBuf
    port map (
            O => \N__39882\,
            I => \N__39879\
        );

    \I__8420\ : CascadeMux
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__8419\ : CascadeBuf
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__39873\,
            I => \N__39870\
        );

    \I__8417\ : CascadeBuf
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__8416\ : CascadeMux
    port map (
            O => \N__39867\,
            I => \N__39864\
        );

    \I__8415\ : CascadeBuf
    port map (
            O => \N__39864\,
            I => \N__39860\
        );

    \I__8414\ : CascadeMux
    port map (
            O => \N__39863\,
            I => \N__39857\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__39860\,
            I => \N__39854\
        );

    \I__8412\ : CascadeBuf
    port map (
            O => \N__39857\,
            I => \N__39851\
        );

    \I__8411\ : CascadeBuf
    port map (
            O => \N__39854\,
            I => \N__39848\
        );

    \I__8410\ : CascadeMux
    port map (
            O => \N__39851\,
            I => \N__39845\
        );

    \I__8409\ : CascadeMux
    port map (
            O => \N__39848\,
            I => \N__39842\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39845\,
            I => \N__39839\
        );

    \I__8407\ : CascadeBuf
    port map (
            O => \N__39842\,
            I => \N__39836\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39839\,
            I => \N__39833\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__39836\,
            I => \N__39830\
        );

    \I__8404\ : Span12Mux_h
    port map (
            O => \N__39833\,
            I => \N__39827\
        );

    \I__8403\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39824\
        );

    \I__8402\ : Span12Mux_v
    port map (
            O => \N__39827\,
            I => \N__39821\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__39824\,
            I => \N__39818\
        );

    \I__8400\ : Odrv12
    port map (
            O => \N__39821\,
            I => \data_index_9_N_212_2\
        );

    \I__8399\ : Odrv12
    port map (
            O => \N__39818\,
            I => \data_index_9_N_212_2\
        );

    \I__8398\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39809\
        );

    \I__8397\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39806\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__39809\,
            I => \N__39803\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__39806\,
            I => \comm_spi.n14815\
        );

    \I__8394\ : Odrv4
    port map (
            O => \N__39803\,
            I => \comm_spi.n14815\
        );

    \I__8393\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39794\
        );

    \I__8392\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39791\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__39794\,
            I => \comm_spi.n14816\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__39791\,
            I => \comm_spi.n14816\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39782\
        );

    \I__8388\ : InMux
    port map (
            O => \N__39785\,
            I => \N__39779\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__39782\,
            I => \comm_spi.imosi\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__39779\,
            I => \comm_spi.imosi\
        );

    \I__8385\ : SRMux
    port map (
            O => \N__39774\,
            I => \N__39771\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39771\,
            I => \N__39768\
        );

    \I__8383\ : Span4Mux_v
    port map (
            O => \N__39768\,
            I => \N__39765\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__39765\,
            I => \N__39762\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__39762\,
            I => \comm_spi.DOUT_7__N_787\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39759\,
            I => \N__39755\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39758\,
            I => \N__39752\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39755\,
            I => wdtick_cnt_0
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__39752\,
            I => wdtick_cnt_0
        );

    \I__8376\ : InMux
    port map (
            O => \N__39747\,
            I => \bfn_15_5_0_\
        );

    \I__8375\ : InMux
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__39741\,
            I => \N__39737\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39740\,
            I => \N__39734\
        );

    \I__8372\ : Span4Mux_h
    port map (
            O => \N__39737\,
            I => \N__39731\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__39734\,
            I => wdtick_cnt_1
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__39731\,
            I => wdtick_cnt_1
        );

    \I__8369\ : InMux
    port map (
            O => \N__39726\,
            I => n19932
        );

    \I__8368\ : InMux
    port map (
            O => \N__39723\,
            I => \N__39719\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39722\,
            I => \N__39716\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__39719\,
            I => wdtick_cnt_2
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__39716\,
            I => wdtick_cnt_2
        );

    \I__8364\ : InMux
    port map (
            O => \N__39711\,
            I => n19933
        );

    \I__8363\ : InMux
    port map (
            O => \N__39708\,
            I => \N__39704\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39707\,
            I => \N__39701\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__39704\,
            I => wdtick_cnt_3
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__39701\,
            I => wdtick_cnt_3
        );

    \I__8359\ : InMux
    port map (
            O => \N__39696\,
            I => n19934
        );

    \I__8358\ : InMux
    port map (
            O => \N__39693\,
            I => \N__39689\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39692\,
            I => \N__39686\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39689\,
            I => wdtick_cnt_4
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39686\,
            I => wdtick_cnt_4
        );

    \I__8354\ : InMux
    port map (
            O => \N__39681\,
            I => n19935
        );

    \I__8353\ : InMux
    port map (
            O => \N__39678\,
            I => \N__39674\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39677\,
            I => \N__39671\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__39674\,
            I => wdtick_cnt_5
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__39671\,
            I => wdtick_cnt_5
        );

    \I__8349\ : InMux
    port map (
            O => \N__39666\,
            I => n19936
        );

    \I__8348\ : InMux
    port map (
            O => \N__39663\,
            I => \N__39659\
        );

    \I__8347\ : InMux
    port map (
            O => \N__39662\,
            I => \N__39656\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__39659\,
            I => \N__39653\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__39656\,
            I => \N__39650\
        );

    \I__8344\ : Span4Mux_v
    port map (
            O => \N__39653\,
            I => \N__39646\
        );

    \I__8343\ : Span4Mux_h
    port map (
            O => \N__39650\,
            I => \N__39643\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39636\
        );

    \I__8341\ : Span4Mux_h
    port map (
            O => \N__39646\,
            I => \N__39631\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__39643\,
            I => \N__39631\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39628\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39641\,
            I => \N__39625\
        );

    \I__8337\ : InMux
    port map (
            O => \N__39640\,
            I => \N__39622\
        );

    \I__8336\ : InMux
    port map (
            O => \N__39639\,
            I => \N__39619\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39616\
        );

    \I__8334\ : Span4Mux_v
    port map (
            O => \N__39631\,
            I => \N__39613\
        );

    \I__8333\ : LocalMux
    port map (
            O => \N__39628\,
            I => n12624
        );

    \I__8332\ : LocalMux
    port map (
            O => \N__39625\,
            I => n12624
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__39622\,
            I => n12624
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__39619\,
            I => n12624
        );

    \I__8329\ : Odrv12
    port map (
            O => \N__39616\,
            I => n12624
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__39613\,
            I => n12624
        );

    \I__8327\ : CascadeMux
    port map (
            O => \N__39600\,
            I => \N__39597\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39592\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39596\,
            I => \N__39589\
        );

    \I__8324\ : CascadeMux
    port map (
            O => \N__39595\,
            I => \N__39586\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__39592\,
            I => \N__39582\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39589\,
            I => \N__39579\
        );

    \I__8321\ : InMux
    port map (
            O => \N__39586\,
            I => \N__39574\
        );

    \I__8320\ : InMux
    port map (
            O => \N__39585\,
            I => \N__39574\
        );

    \I__8319\ : Span4Mux_v
    port map (
            O => \N__39582\,
            I => \N__39567\
        );

    \I__8318\ : Span4Mux_v
    port map (
            O => \N__39579\,
            I => \N__39567\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39574\,
            I => \N__39567\
        );

    \I__8316\ : Span4Mux_h
    port map (
            O => \N__39567\,
            I => \N__39564\
        );

    \I__8315\ : Span4Mux_v
    port map (
            O => \N__39564\,
            I => \N__39560\
        );

    \I__8314\ : CascadeMux
    port map (
            O => \N__39563\,
            I => \N__39557\
        );

    \I__8313\ : Span4Mux_v
    port map (
            O => \N__39560\,
            I => \N__39554\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39557\,
            I => \N__39551\
        );

    \I__8311\ : Span4Mux_h
    port map (
            O => \N__39554\,
            I => \N__39548\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__39551\,
            I => \buf_cfgRTD_1\
        );

    \I__8309\ : Odrv4
    port map (
            O => \N__39548\,
            I => \buf_cfgRTD_1\
        );

    \I__8308\ : InMux
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__39540\,
            I => \N__39535\
        );

    \I__8306\ : InMux
    port map (
            O => \N__39539\,
            I => \N__39532\
        );

    \I__8305\ : InMux
    port map (
            O => \N__39538\,
            I => \N__39529\
        );

    \I__8304\ : Span4Mux_v
    port map (
            O => \N__39535\,
            I => \N__39525\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__39532\,
            I => \N__39520\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__39529\,
            I => \N__39520\
        );

    \I__8301\ : InMux
    port map (
            O => \N__39528\,
            I => \N__39517\
        );

    \I__8300\ : Span4Mux_h
    port map (
            O => \N__39525\,
            I => \N__39509\
        );

    \I__8299\ : Span4Mux_v
    port map (
            O => \N__39520\,
            I => \N__39509\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39506\
        );

    \I__8297\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39503\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39515\,
            I => \N__39498\
        );

    \I__8295\ : InMux
    port map (
            O => \N__39514\,
            I => \N__39498\
        );

    \I__8294\ : Span4Mux_v
    port map (
            O => \N__39509\,
            I => \N__39495\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__39506\,
            I => \N__39490\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__39503\,
            I => \N__39490\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__39498\,
            I => \N__39487\
        );

    \I__8290\ : Sp12to4
    port map (
            O => \N__39495\,
            I => \N__39484\
        );

    \I__8289\ : Span4Mux_v
    port map (
            O => \N__39490\,
            I => \N__39479\
        );

    \I__8288\ : Span4Mux_h
    port map (
            O => \N__39487\,
            I => \N__39479\
        );

    \I__8287\ : Odrv12
    port map (
            O => \N__39484\,
            I => n12610
        );

    \I__8286\ : Odrv4
    port map (
            O => \N__39479\,
            I => n12610
        );

    \I__8285\ : IoInMux
    port map (
            O => \N__39474\,
            I => \N__39471\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__39471\,
            I => \N__39468\
        );

    \I__8283\ : Span4Mux_s0_v
    port map (
            O => \N__39468\,
            I => \N__39465\
        );

    \I__8282\ : Span4Mux_v
    port map (
            O => \N__39465\,
            I => \N__39462\
        );

    \I__8281\ : Span4Mux_v
    port map (
            O => \N__39462\,
            I => \N__39457\
        );

    \I__8280\ : InMux
    port map (
            O => \N__39461\,
            I => \N__39454\
        );

    \I__8279\ : InMux
    port map (
            O => \N__39460\,
            I => \N__39451\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__39457\,
            I => \IAC_OSR0\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__39454\,
            I => \IAC_OSR0\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__39451\,
            I => \IAC_OSR0\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__39444\,
            I => \N__39441\
        );

    \I__8274\ : CascadeBuf
    port map (
            O => \N__39441\,
            I => \N__39438\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__39438\,
            I => \N__39435\
        );

    \I__8272\ : CascadeBuf
    port map (
            O => \N__39435\,
            I => \N__39432\
        );

    \I__8271\ : CascadeMux
    port map (
            O => \N__39432\,
            I => \N__39429\
        );

    \I__8270\ : CascadeBuf
    port map (
            O => \N__39429\,
            I => \N__39426\
        );

    \I__8269\ : CascadeMux
    port map (
            O => \N__39426\,
            I => \N__39423\
        );

    \I__8268\ : CascadeBuf
    port map (
            O => \N__39423\,
            I => \N__39420\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__39420\,
            I => \N__39417\
        );

    \I__8266\ : CascadeBuf
    port map (
            O => \N__39417\,
            I => \N__39414\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__39414\,
            I => \N__39411\
        );

    \I__8264\ : CascadeBuf
    port map (
            O => \N__39411\,
            I => \N__39408\
        );

    \I__8263\ : CascadeMux
    port map (
            O => \N__39408\,
            I => \N__39405\
        );

    \I__8262\ : CascadeBuf
    port map (
            O => \N__39405\,
            I => \N__39402\
        );

    \I__8261\ : CascadeMux
    port map (
            O => \N__39402\,
            I => \N__39398\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__39401\,
            I => \N__39395\
        );

    \I__8259\ : CascadeBuf
    port map (
            O => \N__39398\,
            I => \N__39392\
        );

    \I__8258\ : CascadeBuf
    port map (
            O => \N__39395\,
            I => \N__39389\
        );

    \I__8257\ : CascadeMux
    port map (
            O => \N__39392\,
            I => \N__39386\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__39389\,
            I => \N__39383\
        );

    \I__8255\ : CascadeBuf
    port map (
            O => \N__39386\,
            I => \N__39380\
        );

    \I__8254\ : InMux
    port map (
            O => \N__39383\,
            I => \N__39377\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__39380\,
            I => \N__39374\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__39377\,
            I => \N__39371\
        );

    \I__8251\ : InMux
    port map (
            O => \N__39374\,
            I => \N__39368\
        );

    \I__8250\ : Span12Mux_h
    port map (
            O => \N__39371\,
            I => \N__39365\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__39368\,
            I => \N__39362\
        );

    \I__8248\ : Odrv12
    port map (
            O => \N__39365\,
            I => \data_index_9_N_212_8\
        );

    \I__8247\ : Odrv12
    port map (
            O => \N__39362\,
            I => \data_index_9_N_212_8\
        );

    \I__8246\ : InMux
    port map (
            O => \N__39357\,
            I => \N__39352\
        );

    \I__8245\ : InMux
    port map (
            O => \N__39356\,
            I => \N__39349\
        );

    \I__8244\ : InMux
    port map (
            O => \N__39355\,
            I => \N__39346\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__39352\,
            I => \N__39341\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39349\,
            I => \N__39341\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__39346\,
            I => data_index_1
        );

    \I__8240\ : Odrv4
    port map (
            O => \N__39341\,
            I => data_index_1
        );

    \I__8239\ : InMux
    port map (
            O => \N__39336\,
            I => \N__39333\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__39333\,
            I => n8_adj_1570
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__39330\,
            I => \n8_adj_1570_cascade_\
        );

    \I__8236\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39323\
        );

    \I__8235\ : InMux
    port map (
            O => \N__39326\,
            I => \N__39320\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__39323\,
            I => \N__39315\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__39320\,
            I => \N__39315\
        );

    \I__8232\ : Odrv12
    port map (
            O => \N__39315\,
            I => n7_adj_1569
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__39312\,
            I => \N__39309\
        );

    \I__8230\ : CascadeBuf
    port map (
            O => \N__39309\,
            I => \N__39306\
        );

    \I__8229\ : CascadeMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8228\ : CascadeBuf
    port map (
            O => \N__39303\,
            I => \N__39300\
        );

    \I__8227\ : CascadeMux
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8226\ : CascadeBuf
    port map (
            O => \N__39297\,
            I => \N__39294\
        );

    \I__8225\ : CascadeMux
    port map (
            O => \N__39294\,
            I => \N__39291\
        );

    \I__8224\ : CascadeBuf
    port map (
            O => \N__39291\,
            I => \N__39288\
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__39288\,
            I => \N__39285\
        );

    \I__8222\ : CascadeBuf
    port map (
            O => \N__39285\,
            I => \N__39282\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__39282\,
            I => \N__39279\
        );

    \I__8220\ : CascadeBuf
    port map (
            O => \N__39279\,
            I => \N__39276\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__39276\,
            I => \N__39273\
        );

    \I__8218\ : CascadeBuf
    port map (
            O => \N__39273\,
            I => \N__39269\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__39272\,
            I => \N__39266\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__39269\,
            I => \N__39263\
        );

    \I__8215\ : CascadeBuf
    port map (
            O => \N__39266\,
            I => \N__39260\
        );

    \I__8214\ : CascadeBuf
    port map (
            O => \N__39263\,
            I => \N__39257\
        );

    \I__8213\ : CascadeMux
    port map (
            O => \N__39260\,
            I => \N__39254\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__39257\,
            I => \N__39251\
        );

    \I__8211\ : InMux
    port map (
            O => \N__39254\,
            I => \N__39248\
        );

    \I__8210\ : CascadeBuf
    port map (
            O => \N__39251\,
            I => \N__39245\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__39248\,
            I => \N__39242\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__39245\,
            I => \N__39239\
        );

    \I__8207\ : Span12Mux_s9_h
    port map (
            O => \N__39242\,
            I => \N__39236\
        );

    \I__8206\ : InMux
    port map (
            O => \N__39239\,
            I => \N__39233\
        );

    \I__8205\ : Span12Mux_v
    port map (
            O => \N__39236\,
            I => \N__39230\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__39233\,
            I => \N__39227\
        );

    \I__8203\ : Odrv12
    port map (
            O => \N__39230\,
            I => \data_index_9_N_212_1\
        );

    \I__8202\ : Odrv12
    port map (
            O => \N__39227\,
            I => \data_index_9_N_212_1\
        );

    \I__8201\ : InMux
    port map (
            O => \N__39222\,
            I => \N__39218\
        );

    \I__8200\ : InMux
    port map (
            O => \N__39221\,
            I => \N__39215\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__39218\,
            I => \N__39209\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__39215\,
            I => \N__39209\
        );

    \I__8197\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39206\
        );

    \I__8196\ : Span4Mux_h
    port map (
            O => \N__39209\,
            I => \N__39203\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__39206\,
            I => data_index_2
        );

    \I__8194\ : Odrv4
    port map (
            O => \N__39203\,
            I => data_index_2
        );

    \I__8193\ : InMux
    port map (
            O => \N__39198\,
            I => \N__39192\
        );

    \I__8192\ : InMux
    port map (
            O => \N__39197\,
            I => \N__39192\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__39192\,
            I => n8_adj_1558
        );

    \I__8190\ : InMux
    port map (
            O => \N__39189\,
            I => \N__39183\
        );

    \I__8189\ : InMux
    port map (
            O => \N__39188\,
            I => \N__39183\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__8187\ : Odrv12
    port map (
            O => \N__39180\,
            I => n7_adj_1557
        );

    \I__8186\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39173\
        );

    \I__8185\ : InMux
    port map (
            O => \N__39176\,
            I => \N__39170\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__39173\,
            I => \N__39166\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__39170\,
            I => \N__39163\
        );

    \I__8182\ : InMux
    port map (
            O => \N__39169\,
            I => \N__39160\
        );

    \I__8181\ : Span4Mux_v
    port map (
            O => \N__39166\,
            I => \N__39155\
        );

    \I__8180\ : Span4Mux_h
    port map (
            O => \N__39163\,
            I => \N__39155\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__39160\,
            I => data_index_8
        );

    \I__8178\ : Odrv4
    port map (
            O => \N__39155\,
            I => data_index_8
        );

    \I__8177\ : CascadeMux
    port map (
            O => \N__39150\,
            I => \N__39147\
        );

    \I__8176\ : InMux
    port map (
            O => \N__39147\,
            I => \N__39144\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__39144\,
            I => \N__39139\
        );

    \I__8174\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39136\
        );

    \I__8173\ : CascadeMux
    port map (
            O => \N__39142\,
            I => \N__39133\
        );

    \I__8172\ : Span4Mux_h
    port map (
            O => \N__39139\,
            I => \N__39130\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__39136\,
            I => \N__39127\
        );

    \I__8170\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39124\
        );

    \I__8169\ : Span4Mux_h
    port map (
            O => \N__39130\,
            I => \N__39121\
        );

    \I__8168\ : Span12Mux_v
    port map (
            O => \N__39127\,
            I => \N__39118\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__39124\,
            I => buf_adcdata_iac_16
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__39121\,
            I => buf_adcdata_iac_16
        );

    \I__8165\ : Odrv12
    port map (
            O => \N__39118\,
            I => buf_adcdata_iac_16
        );

    \I__8164\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39108\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__39108\,
            I => \N__39105\
        );

    \I__8162\ : Span4Mux_v
    port map (
            O => \N__39105\,
            I => \N__39100\
        );

    \I__8161\ : InMux
    port map (
            O => \N__39104\,
            I => \N__39097\
        );

    \I__8160\ : InMux
    port map (
            O => \N__39103\,
            I => \N__39094\
        );

    \I__8159\ : Span4Mux_h
    port map (
            O => \N__39100\,
            I => \N__39091\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__39097\,
            I => buf_dds1_8
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__39094\,
            I => buf_dds1_8
        );

    \I__8156\ : Odrv4
    port map (
            O => \N__39091\,
            I => buf_dds1_8
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__39084\,
            I => \n22389_cascade_\
        );

    \I__8154\ : CascadeMux
    port map (
            O => \N__39081\,
            I => \N__39078\
        );

    \I__8153\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39073\
        );

    \I__8152\ : InMux
    port map (
            O => \N__39077\,
            I => \N__39070\
        );

    \I__8151\ : InMux
    port map (
            O => \N__39076\,
            I => \N__39067\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__39073\,
            I => \N__39062\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__39070\,
            I => \N__39062\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__39067\,
            I => buf_dds0_8
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__39062\,
            I => buf_dds0_8
        );

    \I__8146\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39052\
        );

    \I__8145\ : InMux
    port map (
            O => \N__39056\,
            I => \N__39049\
        );

    \I__8144\ : InMux
    port map (
            O => \N__39055\,
            I => \N__39046\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__39052\,
            I => \N__39041\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__39049\,
            I => \N__39041\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__39046\,
            I => data_index_5
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__39041\,
            I => data_index_5
        );

    \I__8139\ : IoInMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39030\
        );

    \I__8137\ : Span4Mux_s0_v
    port map (
            O => \N__39030\,
            I => \N__39027\
        );

    \I__8136\ : Sp12to4
    port map (
            O => \N__39027\,
            I => \N__39023\
        );

    \I__8135\ : CascadeMux
    port map (
            O => \N__39026\,
            I => \N__39020\
        );

    \I__8134\ : Span12Mux_h
    port map (
            O => \N__39023\,
            I => \N__39017\
        );

    \I__8133\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39014\
        );

    \I__8132\ : Odrv12
    port map (
            O => \N__39017\,
            I => \DDS_SCK\
        );

    \I__8131\ : LocalMux
    port map (
            O => \N__39014\,
            I => \DDS_SCK\
        );

    \I__8130\ : InMux
    port map (
            O => \N__39009\,
            I => \N__39006\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__39006\,
            I => \N__39002\
        );

    \I__8128\ : CascadeMux
    port map (
            O => \N__39005\,
            I => \N__38999\
        );

    \I__8127\ : Span4Mux_v
    port map (
            O => \N__39002\,
            I => \N__38996\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38999\,
            I => \N__38993\
        );

    \I__8125\ : Span4Mux_h
    port map (
            O => \N__38996\,
            I => \N__38988\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38993\,
            I => \N__38988\
        );

    \I__8123\ : Odrv4
    port map (
            O => \N__38988\,
            I => tmp_buf_15
        );

    \I__8122\ : IoInMux
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__38982\,
            I => \N__38979\
        );

    \I__8120\ : Span12Mux_s11_v
    port map (
            O => \N__38979\,
            I => \N__38976\
        );

    \I__8119\ : Span12Mux_h
    port map (
            O => \N__38976\,
            I => \N__38972\
        );

    \I__8118\ : InMux
    port map (
            O => \N__38975\,
            I => \N__38969\
        );

    \I__8117\ : Odrv12
    port map (
            O => \N__38972\,
            I => \DDS_MOSI\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__38969\,
            I => \DDS_MOSI\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38959\
        );

    \I__8114\ : InMux
    port map (
            O => \N__38963\,
            I => \N__38956\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38962\,
            I => \N__38953\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__38959\,
            I => data_index_9
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38956\,
            I => data_index_9
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__38953\,
            I => data_index_9
        );

    \I__8109\ : InMux
    port map (
            O => \N__38946\,
            I => \N__38941\
        );

    \I__8108\ : CascadeMux
    port map (
            O => \N__38945\,
            I => \N__38938\
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__38944\,
            I => \N__38935\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__38941\,
            I => \N__38924\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38938\,
            I => \N__38921\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38918\
        );

    \I__8103\ : CascadeMux
    port map (
            O => \N__38934\,
            I => \N__38915\
        );

    \I__8102\ : CascadeMux
    port map (
            O => \N__38933\,
            I => \N__38912\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__38932\,
            I => \N__38909\
        );

    \I__8100\ : CascadeMux
    port map (
            O => \N__38931\,
            I => \N__38906\
        );

    \I__8099\ : CascadeMux
    port map (
            O => \N__38930\,
            I => \N__38903\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__38929\,
            I => \N__38900\
        );

    \I__8097\ : CascadeMux
    port map (
            O => \N__38928\,
            I => \N__38897\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__38927\,
            I => \N__38894\
        );

    \I__8095\ : Span4Mux_h
    port map (
            O => \N__38924\,
            I => \N__38891\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__38921\,
            I => \N__38886\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38918\,
            I => \N__38886\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38877\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38877\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38909\,
            I => \N__38877\
        );

    \I__8089\ : InMux
    port map (
            O => \N__38906\,
            I => \N__38877\
        );

    \I__8088\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38868\
        );

    \I__8087\ : InMux
    port map (
            O => \N__38900\,
            I => \N__38868\
        );

    \I__8086\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38868\
        );

    \I__8085\ : InMux
    port map (
            O => \N__38894\,
            I => \N__38868\
        );

    \I__8084\ : Odrv4
    port map (
            O => \N__38891\,
            I => n10756
        );

    \I__8083\ : Odrv4
    port map (
            O => \N__38886\,
            I => n10756
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__38877\,
            I => n10756
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__38868\,
            I => n10756
        );

    \I__8080\ : InMux
    port map (
            O => \N__38859\,
            I => n19812
        );

    \I__8079\ : InMux
    port map (
            O => \N__38856\,
            I => \N__38853\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__38853\,
            I => \N__38850\
        );

    \I__8077\ : Span4Mux_v
    port map (
            O => \N__38850\,
            I => \N__38847\
        );

    \I__8076\ : Span4Mux_h
    port map (
            O => \N__38847\,
            I => \N__38844\
        );

    \I__8075\ : Span4Mux_h
    port map (
            O => \N__38844\,
            I => \N__38841\
        );

    \I__8074\ : Span4Mux_v
    port map (
            O => \N__38841\,
            I => \N__38838\
        );

    \I__8073\ : Odrv4
    port map (
            O => \N__38838\,
            I => buf_data_iac_1
        );

    \I__8072\ : InMux
    port map (
            O => \N__38835\,
            I => \N__38832\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__38832\,
            I => n22_adj_1617
        );

    \I__8070\ : CascadeMux
    port map (
            O => \N__38829\,
            I => \N__38825\
        );

    \I__8069\ : CascadeMux
    port map (
            O => \N__38828\,
            I => \N__38821\
        );

    \I__8068\ : InMux
    port map (
            O => \N__38825\,
            I => \N__38814\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38824\,
            I => \N__38814\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38814\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__38814\,
            I => \N__38811\
        );

    \I__8064\ : Span4Mux_h
    port map (
            O => \N__38811\,
            I => \N__38807\
        );

    \I__8063\ : CascadeMux
    port map (
            O => \N__38810\,
            I => \N__38804\
        );

    \I__8062\ : Span4Mux_v
    port map (
            O => \N__38807\,
            I => \N__38801\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38804\,
            I => \N__38798\
        );

    \I__8060\ : Sp12to4
    port map (
            O => \N__38801\,
            I => \N__38795\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__38798\,
            I => trig_dds1
        );

    \I__8058\ : Odrv12
    port map (
            O => \N__38795\,
            I => trig_dds1
        );

    \I__8057\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38785\
        );

    \I__8056\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38780\
        );

    \I__8055\ : InMux
    port map (
            O => \N__38788\,
            I => \N__38780\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__38785\,
            I => buf_dds0_7
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__38780\,
            I => buf_dds0_7
        );

    \I__8052\ : InMux
    port map (
            O => \N__38775\,
            I => \N__38765\
        );

    \I__8051\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38765\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38773\,
            I => \N__38759\
        );

    \I__8049\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38754\
        );

    \I__8048\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38754\
        );

    \I__8047\ : CascadeMux
    port map (
            O => \N__38770\,
            I => \N__38739\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__38765\,
            I => \N__38734\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38764\,
            I => \N__38731\
        );

    \I__8044\ : InMux
    port map (
            O => \N__38763\,
            I => \N__38728\
        );

    \I__8043\ : InMux
    port map (
            O => \N__38762\,
            I => \N__38725\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__38759\,
            I => \N__38722\
        );

    \I__8041\ : LocalMux
    port map (
            O => \N__38754\,
            I => \N__38719\
        );

    \I__8040\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38712\
        );

    \I__8039\ : InMux
    port map (
            O => \N__38752\,
            I => \N__38712\
        );

    \I__8038\ : InMux
    port map (
            O => \N__38751\,
            I => \N__38712\
        );

    \I__8037\ : InMux
    port map (
            O => \N__38750\,
            I => \N__38709\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38749\,
            I => \N__38706\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38748\,
            I => \N__38701\
        );

    \I__8034\ : InMux
    port map (
            O => \N__38747\,
            I => \N__38701\
        );

    \I__8033\ : InMux
    port map (
            O => \N__38746\,
            I => \N__38696\
        );

    \I__8032\ : InMux
    port map (
            O => \N__38745\,
            I => \N__38696\
        );

    \I__8031\ : InMux
    port map (
            O => \N__38744\,
            I => \N__38693\
        );

    \I__8030\ : InMux
    port map (
            O => \N__38743\,
            I => \N__38688\
        );

    \I__8029\ : InMux
    port map (
            O => \N__38742\,
            I => \N__38688\
        );

    \I__8028\ : InMux
    port map (
            O => \N__38739\,
            I => \N__38685\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38738\,
            I => \N__38680\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38737\,
            I => \N__38680\
        );

    \I__8025\ : Span4Mux_h
    port map (
            O => \N__38734\,
            I => \N__38673\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__38731\,
            I => \N__38673\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__38728\,
            I => \N__38673\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38725\,
            I => \N__38670\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__38722\,
            I => \N__38665\
        );

    \I__8020\ : Span4Mux_h
    port map (
            O => \N__38719\,
            I => \N__38665\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__38712\,
            I => \N__38662\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__38709\,
            I => \N__38659\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__38706\,
            I => \N__38654\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38701\,
            I => \N__38654\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38696\,
            I => \N__38651\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__38693\,
            I => \N__38644\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__38688\,
            I => \N__38644\
        );

    \I__8012\ : LocalMux
    port map (
            O => \N__38685\,
            I => \N__38644\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__38680\,
            I => \N__38641\
        );

    \I__8010\ : Span4Mux_v
    port map (
            O => \N__38673\,
            I => \N__38635\
        );

    \I__8009\ : Span4Mux_h
    port map (
            O => \N__38670\,
            I => \N__38635\
        );

    \I__8008\ : Span4Mux_h
    port map (
            O => \N__38665\,
            I => \N__38628\
        );

    \I__8007\ : Span4Mux_v
    port map (
            O => \N__38662\,
            I => \N__38628\
        );

    \I__8006\ : Span4Mux_h
    port map (
            O => \N__38659\,
            I => \N__38628\
        );

    \I__8005\ : Span4Mux_h
    port map (
            O => \N__38654\,
            I => \N__38619\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__38651\,
            I => \N__38619\
        );

    \I__8003\ : Span4Mux_v
    port map (
            O => \N__38644\,
            I => \N__38619\
        );

    \I__8002\ : Span4Mux_h
    port map (
            O => \N__38641\,
            I => \N__38619\
        );

    \I__8001\ : InMux
    port map (
            O => \N__38640\,
            I => \N__38616\
        );

    \I__8000\ : Odrv4
    port map (
            O => \N__38635\,
            I => n21079
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__38628\,
            I => n21079
        );

    \I__7998\ : Odrv4
    port map (
            O => \N__38619\,
            I => n21079
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__38616\,
            I => n21079
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__38607\,
            I => \N__38603\
        );

    \I__7995\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38579\
        );

    \I__7994\ : InMux
    port map (
            O => \N__38603\,
            I => \N__38574\
        );

    \I__7993\ : InMux
    port map (
            O => \N__38602\,
            I => \N__38574\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38601\,
            I => \N__38571\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38600\,
            I => \N__38565\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38565\
        );

    \I__7989\ : InMux
    port map (
            O => \N__38598\,
            I => \N__38554\
        );

    \I__7988\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38544\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38544\
        );

    \I__7986\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38544\
        );

    \I__7985\ : InMux
    port map (
            O => \N__38594\,
            I => \N__38533\
        );

    \I__7984\ : InMux
    port map (
            O => \N__38593\,
            I => \N__38533\
        );

    \I__7983\ : InMux
    port map (
            O => \N__38592\,
            I => \N__38533\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38591\,
            I => \N__38533\
        );

    \I__7981\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38533\
        );

    \I__7980\ : InMux
    port map (
            O => \N__38589\,
            I => \N__38528\
        );

    \I__7979\ : InMux
    port map (
            O => \N__38588\,
            I => \N__38528\
        );

    \I__7978\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38515\
        );

    \I__7977\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38515\
        );

    \I__7976\ : InMux
    port map (
            O => \N__38585\,
            I => \N__38515\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38584\,
            I => \N__38515\
        );

    \I__7974\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38515\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38582\,
            I => \N__38515\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38579\,
            I => \N__38510\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__38574\,
            I => \N__38510\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38507\
        );

    \I__7969\ : InMux
    port map (
            O => \N__38570\,
            I => \N__38497\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38494\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__38564\,
            I => \N__38491\
        );

    \I__7966\ : InMux
    port map (
            O => \N__38563\,
            I => \N__38488\
        );

    \I__7965\ : InMux
    port map (
            O => \N__38562\,
            I => \N__38481\
        );

    \I__7964\ : InMux
    port map (
            O => \N__38561\,
            I => \N__38481\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38481\
        );

    \I__7962\ : InMux
    port map (
            O => \N__38559\,
            I => \N__38474\
        );

    \I__7961\ : InMux
    port map (
            O => \N__38558\,
            I => \N__38474\
        );

    \I__7960\ : InMux
    port map (
            O => \N__38557\,
            I => \N__38474\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__38554\,
            I => \N__38471\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38553\,
            I => \N__38468\
        );

    \I__7957\ : InMux
    port map (
            O => \N__38552\,
            I => \N__38463\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38463\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__38544\,
            I => \N__38460\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__38533\,
            I => \N__38443\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38528\,
            I => \N__38438\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__38515\,
            I => \N__38438\
        );

    \I__7951\ : Span4Mux_v
    port map (
            O => \N__38510\,
            I => \N__38435\
        );

    \I__7950\ : Span4Mux_v
    port map (
            O => \N__38507\,
            I => \N__38432\
        );

    \I__7949\ : InMux
    port map (
            O => \N__38506\,
            I => \N__38427\
        );

    \I__7948\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38427\
        );

    \I__7947\ : InMux
    port map (
            O => \N__38504\,
            I => \N__38422\
        );

    \I__7946\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38422\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38502\,
            I => \N__38415\
        );

    \I__7944\ : InMux
    port map (
            O => \N__38501\,
            I => \N__38415\
        );

    \I__7943\ : InMux
    port map (
            O => \N__38500\,
            I => \N__38415\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__38497\,
            I => \N__38412\
        );

    \I__7941\ : Span4Mux_v
    port map (
            O => \N__38494\,
            I => \N__38409\
        );

    \I__7940\ : InMux
    port map (
            O => \N__38491\,
            I => \N__38394\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__38488\,
            I => \N__38385\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__38481\,
            I => \N__38385\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__38474\,
            I => \N__38385\
        );

    \I__7936\ : Span4Mux_h
    port map (
            O => \N__38471\,
            I => \N__38385\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__38468\,
            I => \N__38378\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__38463\,
            I => \N__38378\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__38460\,
            I => \N__38378\
        );

    \I__7932\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38371\
        );

    \I__7931\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38371\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38371\
        );

    \I__7929\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38364\
        );

    \I__7928\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38364\
        );

    \I__7927\ : InMux
    port map (
            O => \N__38454\,
            I => \N__38364\
        );

    \I__7926\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38353\
        );

    \I__7925\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38353\
        );

    \I__7924\ : InMux
    port map (
            O => \N__38451\,
            I => \N__38353\
        );

    \I__7923\ : InMux
    port map (
            O => \N__38450\,
            I => \N__38353\
        );

    \I__7922\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38353\
        );

    \I__7921\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38348\
        );

    \I__7920\ : InMux
    port map (
            O => \N__38447\,
            I => \N__38348\
        );

    \I__7919\ : InMux
    port map (
            O => \N__38446\,
            I => \N__38345\
        );

    \I__7918\ : Sp12to4
    port map (
            O => \N__38443\,
            I => \N__38342\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__38438\,
            I => \N__38335\
        );

    \I__7916\ : Span4Mux_v
    port map (
            O => \N__38435\,
            I => \N__38335\
        );

    \I__7915\ : Span4Mux_h
    port map (
            O => \N__38432\,
            I => \N__38335\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__38427\,
            I => \N__38324\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__38422\,
            I => \N__38324\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__38415\,
            I => \N__38324\
        );

    \I__7911\ : Sp12to4
    port map (
            O => \N__38412\,
            I => \N__38324\
        );

    \I__7910\ : Sp12to4
    port map (
            O => \N__38409\,
            I => \N__38324\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38408\,
            I => \N__38317\
        );

    \I__7908\ : InMux
    port map (
            O => \N__38407\,
            I => \N__38317\
        );

    \I__7907\ : InMux
    port map (
            O => \N__38406\,
            I => \N__38317\
        );

    \I__7906\ : InMux
    port map (
            O => \N__38405\,
            I => \N__38308\
        );

    \I__7905\ : InMux
    port map (
            O => \N__38404\,
            I => \N__38308\
        );

    \I__7904\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38308\
        );

    \I__7903\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38308\
        );

    \I__7902\ : InMux
    port map (
            O => \N__38401\,
            I => \N__38297\
        );

    \I__7901\ : InMux
    port map (
            O => \N__38400\,
            I => \N__38297\
        );

    \I__7900\ : InMux
    port map (
            O => \N__38399\,
            I => \N__38297\
        );

    \I__7899\ : InMux
    port map (
            O => \N__38398\,
            I => \N__38297\
        );

    \I__7898\ : InMux
    port map (
            O => \N__38397\,
            I => \N__38297\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__38394\,
            I => \N__38288\
        );

    \I__7896\ : Span4Mux_v
    port map (
            O => \N__38385\,
            I => \N__38288\
        );

    \I__7895\ : Span4Mux_h
    port map (
            O => \N__38378\,
            I => \N__38288\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38288\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__38364\,
            I => adc_state_0
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__38353\,
            I => adc_state_0
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__38348\,
            I => adc_state_0
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__38345\,
            I => adc_state_0
        );

    \I__7889\ : Odrv12
    port map (
            O => \N__38342\,
            I => adc_state_0
        );

    \I__7888\ : Odrv4
    port map (
            O => \N__38335\,
            I => adc_state_0
        );

    \I__7887\ : Odrv12
    port map (
            O => \N__38324\,
            I => adc_state_0
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__38317\,
            I => adc_state_0
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__38308\,
            I => adc_state_0
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__38297\,
            I => adc_state_0
        );

    \I__7883\ : Odrv4
    port map (
            O => \N__38288\,
            I => adc_state_0
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__38265\,
            I => \N__38260\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__38264\,
            I => \N__38257\
        );

    \I__7880\ : InMux
    port map (
            O => \N__38263\,
            I => \N__38254\
        );

    \I__7879\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38251\
        );

    \I__7878\ : InMux
    port map (
            O => \N__38257\,
            I => \N__38248\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__38254\,
            I => \N__38245\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__38251\,
            I => cmd_rdadctmp_18
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__38248\,
            I => cmd_rdadctmp_18
        );

    \I__7874\ : Odrv12
    port map (
            O => \N__38245\,
            I => cmd_rdadctmp_18
        );

    \I__7873\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38233\
        );

    \I__7872\ : InMux
    port map (
            O => \N__38237\,
            I => \N__38230\
        );

    \I__7871\ : CascadeMux
    port map (
            O => \N__38236\,
            I => \N__38227\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__38233\,
            I => \N__38224\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__38230\,
            I => \N__38221\
        );

    \I__7868\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38218\
        );

    \I__7867\ : Span4Mux_v
    port map (
            O => \N__38224\,
            I => \N__38215\
        );

    \I__7866\ : Span12Mux_s9_v
    port map (
            O => \N__38221\,
            I => \N__38212\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__38218\,
            I => buf_adcdata_iac_10
        );

    \I__7864\ : Odrv4
    port map (
            O => \N__38215\,
            I => buf_adcdata_iac_10
        );

    \I__7863\ : Odrv12
    port map (
            O => \N__38212\,
            I => buf_adcdata_iac_10
        );

    \I__7862\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38202\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__38202\,
            I => n8_adj_1564
        );

    \I__7860\ : InMux
    port map (
            O => \N__38199\,
            I => \N__38196\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__38196\,
            I => \N__38192\
        );

    \I__7858\ : InMux
    port map (
            O => \N__38195\,
            I => \N__38189\
        );

    \I__7857\ : Odrv4
    port map (
            O => \N__38192\,
            I => n7_adj_1563
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__38189\,
            I => n7_adj_1563
        );

    \I__7855\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38179\
        );

    \I__7854\ : InMux
    port map (
            O => \N__38183\,
            I => \N__38176\
        );

    \I__7853\ : InMux
    port map (
            O => \N__38182\,
            I => \N__38173\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__38179\,
            I => \N__38168\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__38176\,
            I => \N__38168\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__38173\,
            I => data_index_4
        );

    \I__7849\ : Odrv4
    port map (
            O => \N__38168\,
            I => data_index_4
        );

    \I__7848\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38160\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__38160\,
            I => \N__38157\
        );

    \I__7846\ : Span4Mux_v
    port map (
            O => \N__38157\,
            I => \N__38154\
        );

    \I__7845\ : Odrv4
    port map (
            O => \N__38154\,
            I => n11611
        );

    \I__7844\ : SRMux
    port map (
            O => \N__38151\,
            I => \N__38146\
        );

    \I__7843\ : SRMux
    port map (
            O => \N__38150\,
            I => \N__38143\
        );

    \I__7842\ : SRMux
    port map (
            O => \N__38149\,
            I => \N__38140\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__38146\,
            I => \N__38136\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__38143\,
            I => \N__38133\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38130\
        );

    \I__7838\ : SRMux
    port map (
            O => \N__38139\,
            I => \N__38127\
        );

    \I__7837\ : Span4Mux_h
    port map (
            O => \N__38136\,
            I => \N__38124\
        );

    \I__7836\ : Span4Mux_v
    port map (
            O => \N__38133\,
            I => \N__38121\
        );

    \I__7835\ : Span4Mux_h
    port map (
            O => \N__38130\,
            I => \N__38118\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__38115\
        );

    \I__7833\ : Odrv4
    port map (
            O => \N__38124\,
            I => n14907
        );

    \I__7832\ : Odrv4
    port map (
            O => \N__38121\,
            I => n14907
        );

    \I__7831\ : Odrv4
    port map (
            O => \N__38118\,
            I => n14907
        );

    \I__7830\ : Odrv4
    port map (
            O => \N__38115\,
            I => n14907
        );

    \I__7829\ : InMux
    port map (
            O => \N__38106\,
            I => \bfn_14_15_0_\
        );

    \I__7828\ : InMux
    port map (
            O => \N__38103\,
            I => n19804
        );

    \I__7827\ : InMux
    port map (
            O => \N__38100\,
            I => n19805
        );

    \I__7826\ : InMux
    port map (
            O => \N__38097\,
            I => \N__38092\
        );

    \I__7825\ : InMux
    port map (
            O => \N__38096\,
            I => \N__38089\
        );

    \I__7824\ : InMux
    port map (
            O => \N__38095\,
            I => \N__38086\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__38092\,
            I => data_index_3
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__38089\,
            I => data_index_3
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__38086\,
            I => data_index_3
        );

    \I__7820\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38075\
        );

    \I__7819\ : InMux
    port map (
            O => \N__38078\,
            I => \N__38072\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__38075\,
            I => n7_adj_1565
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__38072\,
            I => n7_adj_1565
        );

    \I__7816\ : InMux
    port map (
            O => \N__38067\,
            I => n19806
        );

    \I__7815\ : InMux
    port map (
            O => \N__38064\,
            I => n19807
        );

    \I__7814\ : InMux
    port map (
            O => \N__38061\,
            I => n19808
        );

    \I__7813\ : InMux
    port map (
            O => \N__38058\,
            I => \N__38054\
        );

    \I__7812\ : InMux
    port map (
            O => \N__38057\,
            I => \N__38051\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__38054\,
            I => \N__38045\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__38051\,
            I => \N__38045\
        );

    \I__7809\ : InMux
    port map (
            O => \N__38050\,
            I => \N__38042\
        );

    \I__7808\ : Span4Mux_h
    port map (
            O => \N__38045\,
            I => \N__38039\
        );

    \I__7807\ : LocalMux
    port map (
            O => \N__38042\,
            I => data_index_6
        );

    \I__7806\ : Odrv4
    port map (
            O => \N__38039\,
            I => data_index_6
        );

    \I__7805\ : CascadeMux
    port map (
            O => \N__38034\,
            I => \N__38030\
        );

    \I__7804\ : InMux
    port map (
            O => \N__38033\,
            I => \N__38027\
        );

    \I__7803\ : InMux
    port map (
            O => \N__38030\,
            I => \N__38024\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__38027\,
            I => \N__38021\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__38024\,
            I => \N__38018\
        );

    \I__7800\ : Odrv12
    port map (
            O => \N__38021\,
            I => n7_adj_1561
        );

    \I__7799\ : Odrv4
    port map (
            O => \N__38018\,
            I => n7_adj_1561
        );

    \I__7798\ : InMux
    port map (
            O => \N__38013\,
            I => n19809
        );

    \I__7797\ : InMux
    port map (
            O => \N__38010\,
            I => \N__38005\
        );

    \I__7796\ : InMux
    port map (
            O => \N__38009\,
            I => \N__38002\
        );

    \I__7795\ : InMux
    port map (
            O => \N__38008\,
            I => \N__37999\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__38005\,
            I => \N__37994\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__38002\,
            I => \N__37994\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37999\,
            I => data_index_7
        );

    \I__7791\ : Odrv12
    port map (
            O => \N__37994\,
            I => data_index_7
        );

    \I__7790\ : InMux
    port map (
            O => \N__37989\,
            I => \N__37983\
        );

    \I__7789\ : InMux
    port map (
            O => \N__37988\,
            I => \N__37983\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__7787\ : Odrv4
    port map (
            O => \N__37980\,
            I => n7_adj_1559
        );

    \I__7786\ : InMux
    port map (
            O => \N__37977\,
            I => n19810
        );

    \I__7785\ : InMux
    port map (
            O => \N__37974\,
            I => \bfn_14_16_0_\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37971\,
            I => \bfn_14_14_0_\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37968\,
            I => n19782
        );

    \I__7782\ : InMux
    port map (
            O => \N__37965\,
            I => n19783
        );

    \I__7781\ : InMux
    port map (
            O => \N__37962\,
            I => \N__37959\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__37959\,
            I => \N__37956\
        );

    \I__7779\ : Span4Mux_h
    port map (
            O => \N__37956\,
            I => \N__37951\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37955\,
            I => \N__37948\
        );

    \I__7777\ : InMux
    port map (
            O => \N__37954\,
            I => \N__37945\
        );

    \I__7776\ : Span4Mux_v
    port map (
            O => \N__37951\,
            I => \N__37942\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__37948\,
            I => \N__37939\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37945\,
            I => data_cntvec_11
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__37942\,
            I => data_cntvec_11
        );

    \I__7772\ : Odrv12
    port map (
            O => \N__37939\,
            I => data_cntvec_11
        );

    \I__7771\ : InMux
    port map (
            O => \N__37932\,
            I => n19784
        );

    \I__7770\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37926\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__37926\,
            I => \N__37922\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37925\,
            I => \N__37919\
        );

    \I__7767\ : Span4Mux_v
    port map (
            O => \N__37922\,
            I => \N__37916\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37919\,
            I => data_cntvec_12
        );

    \I__7765\ : Odrv4
    port map (
            O => \N__37916\,
            I => data_cntvec_12
        );

    \I__7764\ : InMux
    port map (
            O => \N__37911\,
            I => n19785
        );

    \I__7763\ : InMux
    port map (
            O => \N__37908\,
            I => \N__37905\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37905\,
            I => \N__37901\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37898\
        );

    \I__7760\ : Span4Mux_h
    port map (
            O => \N__37901\,
            I => \N__37895\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__37898\,
            I => data_cntvec_13
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__37895\,
            I => data_cntvec_13
        );

    \I__7757\ : InMux
    port map (
            O => \N__37890\,
            I => n19786
        );

    \I__7756\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37884\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__37884\,
            I => \N__37880\
        );

    \I__7754\ : InMux
    port map (
            O => \N__37883\,
            I => \N__37877\
        );

    \I__7753\ : Span12Mux_v
    port map (
            O => \N__37880\,
            I => \N__37874\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37877\,
            I => data_cntvec_14
        );

    \I__7751\ : Odrv12
    port map (
            O => \N__37874\,
            I => data_cntvec_14
        );

    \I__7750\ : InMux
    port map (
            O => \N__37869\,
            I => n19787
        );

    \I__7749\ : InMux
    port map (
            O => \N__37866\,
            I => n19788
        );

    \I__7748\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37860\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__37860\,
            I => \N__37856\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37859\,
            I => \N__37853\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__37856\,
            I => \N__37850\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__37853\,
            I => data_cntvec_15
        );

    \I__7743\ : Odrv4
    port map (
            O => \N__37850\,
            I => data_cntvec_15
        );

    \I__7742\ : CEMux
    port map (
            O => \N__37845\,
            I => \N__37839\
        );

    \I__7741\ : CEMux
    port map (
            O => \N__37844\,
            I => \N__37836\
        );

    \I__7740\ : CEMux
    port map (
            O => \N__37843\,
            I => \N__37833\
        );

    \I__7739\ : CEMux
    port map (
            O => \N__37842\,
            I => \N__37830\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37839\,
            I => \N__37827\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__37836\,
            I => \N__37824\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37833\,
            I => \N__37821\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__37830\,
            I => \N__37818\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__37827\,
            I => \N__37815\
        );

    \I__7733\ : Span4Mux_h
    port map (
            O => \N__37824\,
            I => \N__37812\
        );

    \I__7732\ : Span4Mux_h
    port map (
            O => \N__37821\,
            I => \N__37809\
        );

    \I__7731\ : Span4Mux_h
    port map (
            O => \N__37818\,
            I => \N__37805\
        );

    \I__7730\ : Span4Mux_v
    port map (
            O => \N__37815\,
            I => \N__37802\
        );

    \I__7729\ : Span4Mux_h
    port map (
            O => \N__37812\,
            I => \N__37797\
        );

    \I__7728\ : Span4Mux_h
    port map (
            O => \N__37809\,
            I => \N__37797\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37794\
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__37805\,
            I => n11933
        );

    \I__7725\ : Odrv4
    port map (
            O => \N__37802\,
            I => n11933
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__37797\,
            I => n11933
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__37794\,
            I => n11933
        );

    \I__7722\ : CascadeMux
    port map (
            O => \N__37785\,
            I => \N__37781\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__37784\,
            I => \N__37776\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37781\,
            I => \N__37773\
        );

    \I__7719\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37766\
        );

    \I__7718\ : InMux
    port map (
            O => \N__37779\,
            I => \N__37766\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37776\,
            I => \N__37763\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__37773\,
            I => \N__37760\
        );

    \I__7715\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37757\
        );

    \I__7714\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37754\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__37766\,
            I => \N__37751\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37748\
        );

    \I__7711\ : Sp12to4
    port map (
            O => \N__37760\,
            I => \N__37743\
        );

    \I__7710\ : LocalMux
    port map (
            O => \N__37757\,
            I => \N__37743\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__37754\,
            I => \N__37736\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__37751\,
            I => \N__37736\
        );

    \I__7707\ : Span4Mux_h
    port map (
            O => \N__37748\,
            I => \N__37736\
        );

    \I__7706\ : Span12Mux_v
    port map (
            O => \N__37743\,
            I => \N__37733\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__37736\,
            I => \iac_raw_buf_N_776\
        );

    \I__7704\ : Odrv12
    port map (
            O => \N__37733\,
            I => \iac_raw_buf_N_776\
        );

    \I__7703\ : InMux
    port map (
            O => \N__37728\,
            I => n19774
        );

    \I__7702\ : InMux
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__37722\,
            I => \N__37718\
        );

    \I__7700\ : InMux
    port map (
            O => \N__37721\,
            I => \N__37714\
        );

    \I__7699\ : Span4Mux_v
    port map (
            O => \N__37718\,
            I => \N__37711\
        );

    \I__7698\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37708\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__37714\,
            I => data_cntvec_2
        );

    \I__7696\ : Odrv4
    port map (
            O => \N__37711\,
            I => data_cntvec_2
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__37708\,
            I => data_cntvec_2
        );

    \I__7694\ : InMux
    port map (
            O => \N__37701\,
            I => n19775
        );

    \I__7693\ : InMux
    port map (
            O => \N__37698\,
            I => n19776
        );

    \I__7692\ : InMux
    port map (
            O => \N__37695\,
            I => \N__37692\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37692\,
            I => \N__37687\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37684\
        );

    \I__7689\ : InMux
    port map (
            O => \N__37690\,
            I => \N__37681\
        );

    \I__7688\ : Span4Mux_h
    port map (
            O => \N__37687\,
            I => \N__37678\
        );

    \I__7687\ : LocalMux
    port map (
            O => \N__37684\,
            I => data_cntvec_4
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__37681\,
            I => data_cntvec_4
        );

    \I__7685\ : Odrv4
    port map (
            O => \N__37678\,
            I => data_cntvec_4
        );

    \I__7684\ : InMux
    port map (
            O => \N__37671\,
            I => n19777
        );

    \I__7683\ : InMux
    port map (
            O => \N__37668\,
            I => \N__37664\
        );

    \I__7682\ : InMux
    port map (
            O => \N__37667\,
            I => \N__37661\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__37664\,
            I => \N__37657\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__37661\,
            I => \N__37654\
        );

    \I__7679\ : InMux
    port map (
            O => \N__37660\,
            I => \N__37651\
        );

    \I__7678\ : Span4Mux_h
    port map (
            O => \N__37657\,
            I => \N__37648\
        );

    \I__7677\ : Span4Mux_h
    port map (
            O => \N__37654\,
            I => \N__37645\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__37651\,
            I => data_cntvec_5
        );

    \I__7675\ : Odrv4
    port map (
            O => \N__37648\,
            I => data_cntvec_5
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__37645\,
            I => data_cntvec_5
        );

    \I__7673\ : InMux
    port map (
            O => \N__37638\,
            I => n19778
        );

    \I__7672\ : InMux
    port map (
            O => \N__37635\,
            I => n19779
        );

    \I__7671\ : InMux
    port map (
            O => \N__37632\,
            I => n19780
        );

    \I__7670\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37626\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__37626\,
            I => \N__37623\
        );

    \I__7668\ : Span4Mux_h
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__37617\,
            I => n22380
        );

    \I__7665\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37611\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37611\,
            I => \N__37608\
        );

    \I__7663\ : Span4Mux_v
    port map (
            O => \N__37608\,
            I => \N__37605\
        );

    \I__7662\ : Odrv4
    port map (
            O => \N__37605\,
            I => n30_adj_1679
        );

    \I__7661\ : CascadeMux
    port map (
            O => \N__37602\,
            I => \n8_adj_1689_cascade_\
        );

    \I__7660\ : CascadeMux
    port map (
            O => \N__37599\,
            I => \n26_adj_1595_cascade_\
        );

    \I__7659\ : CEMux
    port map (
            O => \N__37596\,
            I => \N__37593\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__37593\,
            I => n18_adj_1615
        );

    \I__7657\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37586\
        );

    \I__7656\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37583\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__37586\,
            I => \N__37579\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__37583\,
            I => \N__37576\
        );

    \I__7653\ : CascadeMux
    port map (
            O => \N__37582\,
            I => \N__37573\
        );

    \I__7652\ : Span4Mux_h
    port map (
            O => \N__37579\,
            I => \N__37567\
        );

    \I__7651\ : Span4Mux_h
    port map (
            O => \N__37576\,
            I => \N__37564\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37573\,
            I => \N__37557\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37572\,
            I => \N__37557\
        );

    \I__7648\ : InMux
    port map (
            O => \N__37571\,
            I => \N__37557\
        );

    \I__7647\ : InMux
    port map (
            O => \N__37570\,
            I => \N__37554\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__37567\,
            I => n16818
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__37564\,
            I => n16818
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37557\,
            I => n16818
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__37554\,
            I => n16818
        );

    \I__7642\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37542\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__37542\,
            I => n21714
        );

    \I__7640\ : CascadeMux
    port map (
            O => \N__37539\,
            I => \n7_cascade_\
        );

    \I__7639\ : InMux
    port map (
            O => \N__37536\,
            I => \N__37533\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37533\,
            I => \N__37528\
        );

    \I__7637\ : InMux
    port map (
            O => \N__37532\,
            I => \N__37525\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37531\,
            I => \N__37519\
        );

    \I__7635\ : Span4Mux_v
    port map (
            O => \N__37528\,
            I => \N__37514\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__37525\,
            I => \N__37514\
        );

    \I__7633\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37509\
        );

    \I__7632\ : InMux
    port map (
            O => \N__37523\,
            I => \N__37509\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37506\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__37519\,
            I => \N__37503\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__37514\,
            I => \N__37498\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__37509\,
            I => \N__37498\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__37506\,
            I => \N__37493\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__37503\,
            I => \N__37488\
        );

    \I__7625\ : Span4Mux_h
    port map (
            O => \N__37498\,
            I => \N__37488\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37483\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37496\,
            I => \N__37483\
        );

    \I__7622\ : Odrv12
    port map (
            O => \N__37493\,
            I => n12107
        );

    \I__7621\ : Odrv4
    port map (
            O => \N__37488\,
            I => n12107
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__37483\,
            I => n12107
        );

    \I__7619\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37473\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__37473\,
            I => \N__37469\
        );

    \I__7617\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37466\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__37469\,
            I => \N__37461\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37466\,
            I => \N__37461\
        );

    \I__7614\ : Span4Mux_v
    port map (
            O => \N__37461\,
            I => \N__37458\
        );

    \I__7613\ : Sp12to4
    port map (
            O => \N__37458\,
            I => \N__37455\
        );

    \I__7612\ : Odrv12
    port map (
            O => \N__37455\,
            I => n14_adj_1544
        );

    \I__7611\ : InMux
    port map (
            O => \N__37452\,
            I => \N__37449\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37449\,
            I => \N__37446\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__37446\,
            I => \N__37442\
        );

    \I__7608\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37439\
        );

    \I__7607\ : Sp12to4
    port map (
            O => \N__37442\,
            I => \N__37436\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__37439\,
            I => n14_adj_1575
        );

    \I__7605\ : Odrv12
    port map (
            O => \N__37436\,
            I => n14_adj_1575
        );

    \I__7604\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37428\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__37428\,
            I => \N__37425\
        );

    \I__7602\ : Odrv12
    port map (
            O => \N__37425\,
            I => n19_adj_1666
        );

    \I__7601\ : CascadeMux
    port map (
            O => \N__37422\,
            I => \N__37419\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37419\,
            I => \N__37416\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__37416\,
            I => n20_adj_1667
        );

    \I__7598\ : InMux
    port map (
            O => \N__37413\,
            I => \N__37410\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__37410\,
            I => n16_adj_1664
        );

    \I__7596\ : InMux
    port map (
            O => \N__37407\,
            I => \N__37404\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__37404\,
            I => \N__37401\
        );

    \I__7594\ : Odrv12
    port map (
            O => \N__37401\,
            I => n17_adj_1665
        );

    \I__7593\ : CascadeMux
    port map (
            O => \N__37398\,
            I => \n22413_cascade_\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__7591\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__7589\ : Span4Mux_v
    port map (
            O => \N__37386\,
            I => \N__37383\
        );

    \I__7588\ : Odrv4
    port map (
            O => \N__37383\,
            I => n21671
        );

    \I__7587\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37377\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__7585\ : Span4Mux_v
    port map (
            O => \N__37374\,
            I => \N__37371\
        );

    \I__7584\ : Span4Mux_h
    port map (
            O => \N__37371\,
            I => \N__37368\
        );

    \I__7583\ : Odrv4
    port map (
            O => \N__37368\,
            I => n23_adj_1668
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__37365\,
            I => \n22569_cascade_\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37359\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__37359\,
            I => n21702
        );

    \I__7579\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37353\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__37353\,
            I => n22416
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__37350\,
            I => \n22572_cascade_\
        );

    \I__7576\ : CascadeMux
    port map (
            O => \N__37347\,
            I => \n30_adj_1669_cascade_\
        );

    \I__7575\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37341\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__37341\,
            I => \N__37338\
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__37338\,
            I => n22404
        );

    \I__7572\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37332\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__37329\,
            I => \N__37326\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__37326\,
            I => n19_adj_1673
        );

    \I__7568\ : CascadeMux
    port map (
            O => \N__37323\,
            I => \N__37320\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37317\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__37317\,
            I => n20_adj_1674
        );

    \I__7565\ : InMux
    port map (
            O => \N__37314\,
            I => \N__37304\
        );

    \I__7564\ : InMux
    port map (
            O => \N__37313\,
            I => \N__37304\
        );

    \I__7563\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37304\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37311\,
            I => \N__37301\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__37304\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37301\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__7559\ : InMux
    port map (
            O => \N__37296\,
            I => \N__37289\
        );

    \I__7558\ : InMux
    port map (
            O => \N__37295\,
            I => \N__37289\
        );

    \I__7557\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37286\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__37289\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__37286\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__37281\,
            I => \N__37278\
        );

    \I__7553\ : InMux
    port map (
            O => \N__37278\,
            I => \N__37265\
        );

    \I__7552\ : InMux
    port map (
            O => \N__37277\,
            I => \N__37265\
        );

    \I__7551\ : InMux
    port map (
            O => \N__37276\,
            I => \N__37265\
        );

    \I__7550\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37265\
        );

    \I__7549\ : InMux
    port map (
            O => \N__37274\,
            I => \N__37262\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__37265\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__37262\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__7546\ : CascadeMux
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__7545\ : InMux
    port map (
            O => \N__37254\,
            I => \N__37251\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__37251\,
            I => \N__37246\
        );

    \I__7543\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37243\
        );

    \I__7542\ : InMux
    port map (
            O => \N__37249\,
            I => \N__37240\
        );

    \I__7541\ : Span4Mux_h
    port map (
            O => \N__37246\,
            I => \N__37237\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__37243\,
            I => \N__37234\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__37240\,
            I => \N__37231\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__37237\,
            I => \N__37228\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__37234\,
            I => \N__37225\
        );

    \I__7536\ : Span4Mux_v
    port map (
            O => \N__37231\,
            I => \N__37222\
        );

    \I__7535\ : Span4Mux_v
    port map (
            O => \N__37228\,
            I => \N__37219\
        );

    \I__7534\ : Span4Mux_h
    port map (
            O => \N__37225\,
            I => \N__37216\
        );

    \I__7533\ : Span4Mux_h
    port map (
            O => \N__37222\,
            I => \N__37213\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__37219\,
            I => n14_adj_1579
        );

    \I__7531\ : Odrv4
    port map (
            O => \N__37216\,
            I => n14_adj_1579
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__37213\,
            I => n14_adj_1579
        );

    \I__7529\ : InMux
    port map (
            O => \N__37206\,
            I => \N__37203\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__37203\,
            I => \N__37200\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__37200\,
            I => \N__37197\
        );

    \I__7526\ : Span4Mux_h
    port map (
            O => \N__37197\,
            I => \N__37193\
        );

    \I__7525\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37190\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__37193\,
            I => \N__37187\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__37190\,
            I => n14_adj_1572
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__37187\,
            I => n14_adj_1572
        );

    \I__7521\ : InMux
    port map (
            O => \N__37182\,
            I => \N__37179\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__37179\,
            I => \N__37176\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__37176\,
            I => n4_adj_1637
        );

    \I__7518\ : CascadeMux
    port map (
            O => \N__37173\,
            I => \comm_spi.imosi_cascade_\
        );

    \I__7517\ : SRMux
    port map (
            O => \N__37170\,
            I => \N__37167\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__37167\,
            I => \N__37164\
        );

    \I__7515\ : Span4Mux_h
    port map (
            O => \N__37164\,
            I => \N__37161\
        );

    \I__7514\ : Odrv4
    port map (
            O => \N__37161\,
            I => \comm_spi.DOUT_7__N_786\
        );

    \I__7513\ : SRMux
    port map (
            O => \N__37158\,
            I => \N__37155\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__37155\,
            I => \N__37152\
        );

    \I__7511\ : Odrv12
    port map (
            O => \N__37152\,
            I => \comm_spi.imosi_N_792\
        );

    \I__7510\ : CascadeMux
    port map (
            O => \N__37149\,
            I => \n12_adj_1542_cascade_\
        );

    \I__7509\ : CascadeMux
    port map (
            O => \N__37146\,
            I => \n19986_cascade_\
        );

    \I__7508\ : InMux
    port map (
            O => \N__37143\,
            I => \N__37140\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__37140\,
            I => n30_adj_1530
        );

    \I__7506\ : InMux
    port map (
            O => \N__37137\,
            I => \N__37134\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__37134\,
            I => n33
        );

    \I__7504\ : CascadeMux
    port map (
            O => \N__37131\,
            I => \n34_cascade_\
        );

    \I__7503\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37125\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__37125\,
            I => n31
        );

    \I__7501\ : CascadeMux
    port map (
            O => \N__37122\,
            I => \n49_cascade_\
        );

    \I__7500\ : InMux
    port map (
            O => \N__37119\,
            I => \N__37116\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__37116\,
            I => n32
        );

    \I__7498\ : InMux
    port map (
            O => \N__37113\,
            I => \N__37110\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__37110\,
            I => \N__37106\
        );

    \I__7496\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37103\
        );

    \I__7495\ : Span4Mux_h
    port map (
            O => \N__37106\,
            I => \N__37100\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__37103\,
            I => acadc_skipcnt_13
        );

    \I__7493\ : Odrv4
    port map (
            O => \N__37100\,
            I => acadc_skipcnt_13
        );

    \I__7492\ : InMux
    port map (
            O => \N__37095\,
            I => n19801
        );

    \I__7491\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37089\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__37089\,
            I => \N__37086\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__37086\,
            I => \N__37082\
        );

    \I__7488\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37079\
        );

    \I__7487\ : Sp12to4
    port map (
            O => \N__37082\,
            I => \N__37076\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__37079\,
            I => acadc_skipcnt_14
        );

    \I__7485\ : Odrv12
    port map (
            O => \N__37076\,
            I => acadc_skipcnt_14
        );

    \I__7484\ : InMux
    port map (
            O => \N__37071\,
            I => n19802
        );

    \I__7483\ : InMux
    port map (
            O => \N__37068\,
            I => n19803
        );

    \I__7482\ : CascadeMux
    port map (
            O => \N__37065\,
            I => \N__37062\
        );

    \I__7481\ : InMux
    port map (
            O => \N__37062\,
            I => \N__37059\
        );

    \I__7480\ : LocalMux
    port map (
            O => \N__37059\,
            I => \N__37055\
        );

    \I__7479\ : InMux
    port map (
            O => \N__37058\,
            I => \N__37052\
        );

    \I__7478\ : Span12Mux_v
    port map (
            O => \N__37055\,
            I => \N__37049\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__37052\,
            I => acadc_skipcnt_15
        );

    \I__7476\ : Odrv12
    port map (
            O => \N__37049\,
            I => acadc_skipcnt_15
        );

    \I__7475\ : CEMux
    port map (
            O => \N__37044\,
            I => \N__37039\
        );

    \I__7474\ : CEMux
    port map (
            O => \N__37043\,
            I => \N__37036\
        );

    \I__7473\ : CEMux
    port map (
            O => \N__37042\,
            I => \N__37032\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__37039\,
            I => \N__37027\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__37036\,
            I => \N__37027\
        );

    \I__7470\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37024\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__37032\,
            I => \N__37021\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__37027\,
            I => \N__37018\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__37024\,
            I => \N__37015\
        );

    \I__7466\ : Span4Mux_v
    port map (
            O => \N__37021\,
            I => \N__37010\
        );

    \I__7465\ : Span4Mux_h
    port map (
            O => \N__37018\,
            I => \N__37010\
        );

    \I__7464\ : Span4Mux_h
    port map (
            O => \N__37015\,
            I => \N__37007\
        );

    \I__7463\ : Span4Mux_h
    port map (
            O => \N__37010\,
            I => \N__37002\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__37007\,
            I => \N__37002\
        );

    \I__7461\ : Odrv4
    port map (
            O => \N__37002\,
            I => n11989
        );

    \I__7460\ : SRMux
    port map (
            O => \N__36999\,
            I => \N__36995\
        );

    \I__7459\ : SRMux
    port map (
            O => \N__36998\,
            I => \N__36992\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36995\,
            I => \N__36989\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__36992\,
            I => \N__36986\
        );

    \I__7456\ : Span4Mux_v
    port map (
            O => \N__36989\,
            I => \N__36983\
        );

    \I__7455\ : Sp12to4
    port map (
            O => \N__36986\,
            I => \N__36980\
        );

    \I__7454\ : Span4Mux_v
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__7453\ : Odrv12
    port map (
            O => \N__36980\,
            I => n14915
        );

    \I__7452\ : Odrv4
    port map (
            O => \N__36977\,
            I => n14915
        );

    \I__7451\ : InMux
    port map (
            O => \N__36972\,
            I => \N__36967\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36971\,
            I => \N__36964\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36970\,
            I => \N__36961\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__36967\,
            I => \comm_spi.n23083\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__36964\,
            I => \comm_spi.n23083\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__36961\,
            I => \comm_spi.n23083\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__36951\,
            I => \N__36947\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36944\
        );

    \I__7442\ : Span4Mux_h
    port map (
            O => \N__36947\,
            I => \N__36939\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__36944\,
            I => \N__36939\
        );

    \I__7440\ : Span4Mux_v
    port map (
            O => \N__36939\,
            I => \N__36936\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__36936\,
            I => \comm_spi.n14846\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36930\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__36930\,
            I => \N__36926\
        );

    \I__7436\ : InMux
    port map (
            O => \N__36929\,
            I => \N__36923\
        );

    \I__7435\ : Span4Mux_h
    port map (
            O => \N__36926\,
            I => \N__36918\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36923\,
            I => \N__36918\
        );

    \I__7433\ : Span4Mux_v
    port map (
            O => \N__36918\,
            I => \N__36915\
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__36915\,
            I => \comm_spi.n14847\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36908\
        );

    \I__7430\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36905\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__36908\,
            I => \N__36899\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__36905\,
            I => \N__36899\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36904\,
            I => \N__36896\
        );

    \I__7426\ : Odrv4
    port map (
            O => \N__36899\,
            I => \comm_spi.n14808\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36896\,
            I => \comm_spi.n14808\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36891\,
            I => \N__36888\
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__36888\,
            I => \N__36883\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36887\,
            I => \N__36880\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36877\
        );

    \I__7420\ : Span4Mux_v
    port map (
            O => \N__36883\,
            I => \N__36874\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__36880\,
            I => \comm_spi.n14809\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__36877\,
            I => \comm_spi.n14809\
        );

    \I__7417\ : Odrv4
    port map (
            O => \N__36874\,
            I => \comm_spi.n14809\
        );

    \I__7416\ : CascadeMux
    port map (
            O => \N__36867\,
            I => \N__36864\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36860\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36857\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__36860\,
            I => \N__36854\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__36857\,
            I => acadc_skipcnt_5
        );

    \I__7411\ : Odrv4
    port map (
            O => \N__36854\,
            I => acadc_skipcnt_5
        );

    \I__7410\ : InMux
    port map (
            O => \N__36849\,
            I => n19793
        );

    \I__7409\ : CascadeMux
    port map (
            O => \N__36846\,
            I => \N__36843\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36843\,
            I => \N__36839\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36842\,
            I => \N__36836\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36839\,
            I => \N__36833\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__36836\,
            I => acadc_skipcnt_6
        );

    \I__7404\ : Odrv12
    port map (
            O => \N__36833\,
            I => acadc_skipcnt_6
        );

    \I__7403\ : InMux
    port map (
            O => \N__36828\,
            I => n19794
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__36825\,
            I => \N__36822\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36819\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__36819\,
            I => \N__36815\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36812\
        );

    \I__7398\ : Span4Mux_v
    port map (
            O => \N__36815\,
            I => \N__36809\
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__36812\,
            I => acadc_skipcnt_7
        );

    \I__7396\ : Odrv4
    port map (
            O => \N__36809\,
            I => acadc_skipcnt_7
        );

    \I__7395\ : InMux
    port map (
            O => \N__36804\,
            I => n19795
        );

    \I__7394\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__36798\,
            I => \N__36794\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36797\,
            I => \N__36791\
        );

    \I__7391\ : Span4Mux_h
    port map (
            O => \N__36794\,
            I => \N__36788\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__36791\,
            I => acadc_skipcnt_8
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__36788\,
            I => acadc_skipcnt_8
        );

    \I__7388\ : InMux
    port map (
            O => \N__36783\,
            I => n19796
        );

    \I__7387\ : InMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__36777\,
            I => \N__36773\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36776\,
            I => \N__36770\
        );

    \I__7384\ : Span4Mux_h
    port map (
            O => \N__36773\,
            I => \N__36767\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__36770\,
            I => acadc_skipcnt_9
        );

    \I__7382\ : Odrv4
    port map (
            O => \N__36767\,
            I => acadc_skipcnt_9
        );

    \I__7381\ : InMux
    port map (
            O => \N__36762\,
            I => \bfn_13_20_0_\
        );

    \I__7380\ : InMux
    port map (
            O => \N__36759\,
            I => n19798
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__36756\,
            I => \N__36753\
        );

    \I__7378\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36750\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__7376\ : Sp12to4
    port map (
            O => \N__36747\,
            I => \N__36743\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36740\
        );

    \I__7374\ : Span12Mux_v
    port map (
            O => \N__36743\,
            I => \N__36737\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36740\,
            I => acadc_skipcnt_11
        );

    \I__7372\ : Odrv12
    port map (
            O => \N__36737\,
            I => acadc_skipcnt_11
        );

    \I__7371\ : InMux
    port map (
            O => \N__36732\,
            I => n19799
        );

    \I__7370\ : InMux
    port map (
            O => \N__36729\,
            I => n19800
        );

    \I__7369\ : InMux
    port map (
            O => \N__36726\,
            I => \N__36723\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__36723\,
            I => \N__36720\
        );

    \I__7367\ : Span4Mux_v
    port map (
            O => \N__36720\,
            I => \N__36716\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36713\
        );

    \I__7365\ : Span4Mux_h
    port map (
            O => \N__36716\,
            I => \N__36710\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__36713\,
            I => acadc_skipcnt_1
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__36710\,
            I => acadc_skipcnt_1
        );

    \I__7362\ : InMux
    port map (
            O => \N__36705\,
            I => \bfn_13_19_0_\
        );

    \I__7361\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36699\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__36699\,
            I => \N__36695\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36692\
        );

    \I__7358\ : Span4Mux_h
    port map (
            O => \N__36695\,
            I => \N__36689\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36692\,
            I => acadc_skipcnt_2
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__36689\,
            I => acadc_skipcnt_2
        );

    \I__7355\ : InMux
    port map (
            O => \N__36684\,
            I => n19790
        );

    \I__7354\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36677\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36674\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__36677\,
            I => \N__36671\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__36674\,
            I => \N__36666\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__36671\,
            I => \N__36666\
        );

    \I__7349\ : Odrv4
    port map (
            O => \N__36666\,
            I => acadc_skipcnt_3
        );

    \I__7348\ : InMux
    port map (
            O => \N__36663\,
            I => n19791
        );

    \I__7347\ : CascadeMux
    port map (
            O => \N__36660\,
            I => \N__36657\
        );

    \I__7346\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36654\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__36654\,
            I => \N__36650\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36647\
        );

    \I__7343\ : Span4Mux_v
    port map (
            O => \N__36650\,
            I => \N__36644\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__36647\,
            I => acadc_skipcnt_4
        );

    \I__7341\ : Odrv4
    port map (
            O => \N__36644\,
            I => acadc_skipcnt_4
        );

    \I__7340\ : InMux
    port map (
            O => \N__36639\,
            I => n19792
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__36636\,
            I => \n8_adj_1566_cascade_\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36630\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__36630\,
            I => \N__36627\
        );

    \I__7336\ : Span4Mux_h
    port map (
            O => \N__36627\,
            I => \N__36624\
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__36624\,
            I => \SIG_DDS.tmp_buf_6\
        );

    \I__7334\ : InMux
    port map (
            O => \N__36621\,
            I => \N__36618\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__36618\,
            I => \N__36615\
        );

    \I__7332\ : Odrv4
    port map (
            O => \N__36615\,
            I => \SIG_DDS.tmp_buf_7\
        );

    \I__7331\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36609\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36606\
        );

    \I__7329\ : Span4Mux_h
    port map (
            O => \N__36606\,
            I => \N__36602\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36605\,
            I => \N__36599\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__36602\,
            I => \N__36596\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__36599\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__36596\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__7324\ : InMux
    port map (
            O => \N__36591\,
            I => \N__36588\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36588\,
            I => \N__36585\
        );

    \I__7322\ : Span4Mux_v
    port map (
            O => \N__36585\,
            I => \N__36582\
        );

    \I__7321\ : Span4Mux_h
    port map (
            O => \N__36582\,
            I => \N__36579\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__36579\,
            I => \SIG_DDS.n21744\
        );

    \I__7319\ : InMux
    port map (
            O => \N__36576\,
            I => \N__36573\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__36573\,
            I => \N__36570\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__36570\,
            I => \N__36565\
        );

    \I__7316\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36562\
        );

    \I__7315\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36559\
        );

    \I__7314\ : Span4Mux_h
    port map (
            O => \N__36565\,
            I => \N__36556\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__36562\,
            I => \N__36553\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__36559\,
            I => buf_dds1_7
        );

    \I__7311\ : Odrv4
    port map (
            O => \N__36556\,
            I => buf_dds1_7
        );

    \I__7310\ : Odrv12
    port map (
            O => \N__36553\,
            I => buf_dds1_7
        );

    \I__7309\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36542\
        );

    \I__7308\ : CascadeMux
    port map (
            O => \N__36545\,
            I => \N__36539\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__36542\,
            I => \N__36536\
        );

    \I__7306\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36533\
        );

    \I__7305\ : Span4Mux_v
    port map (
            O => \N__36536\,
            I => \N__36530\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__36533\,
            I => acadc_skipcnt_0
        );

    \I__7303\ : Odrv4
    port map (
            O => \N__36530\,
            I => acadc_skipcnt_0
        );

    \I__7302\ : SRMux
    port map (
            O => \N__36525\,
            I => \N__36522\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__36522\,
            I => \N__36519\
        );

    \I__7300\ : Span4Mux_v
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__36516\,
            I => n21226
        );

    \I__7298\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36507\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36512\,
            I => \N__36507\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36507\,
            I => \N__36504\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__36504\,
            I => n20011
        );

    \I__7294\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36498\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36498\,
            I => \N__36495\
        );

    \I__7292\ : Span4Mux_h
    port map (
            O => \N__36495\,
            I => \N__36492\
        );

    \I__7291\ : Span4Mux_v
    port map (
            O => \N__36492\,
            I => \N__36489\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__36489\,
            I => n19_adj_1616
        );

    \I__7289\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36482\
        );

    \I__7288\ : InMux
    port map (
            O => \N__36485\,
            I => \N__36478\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36482\,
            I => \N__36475\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36481\,
            I => \N__36472\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__36478\,
            I => \N__36467\
        );

    \I__7284\ : Span4Mux_v
    port map (
            O => \N__36475\,
            I => \N__36467\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__36472\,
            I => \N__36462\
        );

    \I__7282\ : Span4Mux_h
    port map (
            O => \N__36467\,
            I => \N__36459\
        );

    \I__7281\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36454\
        );

    \I__7280\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36454\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__36462\,
            I => \N__36451\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__36459\,
            I => \N__36448\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__36454\,
            I => n14_adj_1547
        );

    \I__7276\ : Odrv4
    port map (
            O => \N__36451\,
            I => n14_adj_1547
        );

    \I__7275\ : Odrv4
    port map (
            O => \N__36448\,
            I => n14_adj_1547
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__36441\,
            I => \n8_adj_1564_cascade_\
        );

    \I__7273\ : CascadeMux
    port map (
            O => \N__36438\,
            I => \N__36435\
        );

    \I__7272\ : CascadeBuf
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__7271\ : CascadeMux
    port map (
            O => \N__36432\,
            I => \N__36429\
        );

    \I__7270\ : CascadeBuf
    port map (
            O => \N__36429\,
            I => \N__36426\
        );

    \I__7269\ : CascadeMux
    port map (
            O => \N__36426\,
            I => \N__36423\
        );

    \I__7268\ : CascadeBuf
    port map (
            O => \N__36423\,
            I => \N__36420\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__36420\,
            I => \N__36417\
        );

    \I__7266\ : CascadeBuf
    port map (
            O => \N__36417\,
            I => \N__36414\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__36414\,
            I => \N__36411\
        );

    \I__7264\ : CascadeBuf
    port map (
            O => \N__36411\,
            I => \N__36408\
        );

    \I__7263\ : CascadeMux
    port map (
            O => \N__36408\,
            I => \N__36405\
        );

    \I__7262\ : CascadeBuf
    port map (
            O => \N__36405\,
            I => \N__36402\
        );

    \I__7261\ : CascadeMux
    port map (
            O => \N__36402\,
            I => \N__36399\
        );

    \I__7260\ : CascadeBuf
    port map (
            O => \N__36399\,
            I => \N__36396\
        );

    \I__7259\ : CascadeMux
    port map (
            O => \N__36396\,
            I => \N__36393\
        );

    \I__7258\ : CascadeBuf
    port map (
            O => \N__36393\,
            I => \N__36389\
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__36392\,
            I => \N__36386\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__36389\,
            I => \N__36383\
        );

    \I__7255\ : CascadeBuf
    port map (
            O => \N__36386\,
            I => \N__36380\
        );

    \I__7254\ : CascadeBuf
    port map (
            O => \N__36383\,
            I => \N__36377\
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__36380\,
            I => \N__36374\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__36377\,
            I => \N__36371\
        );

    \I__7251\ : InMux
    port map (
            O => \N__36374\,
            I => \N__36368\
        );

    \I__7250\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36365\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__36368\,
            I => \N__36362\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__36365\,
            I => \N__36359\
        );

    \I__7247\ : Span12Mux_h
    port map (
            O => \N__36362\,
            I => \N__36354\
        );

    \I__7246\ : Span12Mux_h
    port map (
            O => \N__36359\,
            I => \N__36354\
        );

    \I__7245\ : Odrv12
    port map (
            O => \N__36354\,
            I => \data_index_9_N_212_4\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__36351\,
            I => \N__36348\
        );

    \I__7243\ : InMux
    port map (
            O => \N__36348\,
            I => \N__36345\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__36345\,
            I => \N__36341\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__36344\,
            I => \N__36338\
        );

    \I__7240\ : Span4Mux_v
    port map (
            O => \N__36341\,
            I => \N__36335\
        );

    \I__7239\ : InMux
    port map (
            O => \N__36338\,
            I => \N__36332\
        );

    \I__7238\ : Span4Mux_h
    port map (
            O => \N__36335\,
            I => \N__36328\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__36332\,
            I => \N__36325\
        );

    \I__7236\ : InMux
    port map (
            O => \N__36331\,
            I => \N__36322\
        );

    \I__7235\ : Odrv4
    port map (
            O => \N__36328\,
            I => cmd_rdadctmp_9
        );

    \I__7234\ : Odrv4
    port map (
            O => \N__36325\,
            I => cmd_rdadctmp_9
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36322\,
            I => cmd_rdadctmp_9
        );

    \I__7232\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36312\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__36312\,
            I => \N__36309\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__7229\ : Sp12to4
    port map (
            O => \N__36306\,
            I => \N__36303\
        );

    \I__7228\ : Span12Mux_h
    port map (
            O => \N__36303\,
            I => \N__36298\
        );

    \I__7227\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36293\
        );

    \I__7226\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36293\
        );

    \I__7225\ : Odrv12
    port map (
            O => \N__36298\,
            I => buf_adcdata_iac_1
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__36293\,
            I => buf_adcdata_iac_1
        );

    \I__7223\ : InMux
    port map (
            O => \N__36288\,
            I => \N__36284\
        );

    \I__7222\ : InMux
    port map (
            O => \N__36287\,
            I => \N__36281\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__36284\,
            I => \N__36278\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__36281\,
            I => \N__36274\
        );

    \I__7219\ : Span4Mux_h
    port map (
            O => \N__36278\,
            I => \N__36271\
        );

    \I__7218\ : InMux
    port map (
            O => \N__36277\,
            I => \N__36268\
        );

    \I__7217\ : Span4Mux_v
    port map (
            O => \N__36274\,
            I => \N__36263\
        );

    \I__7216\ : Span4Mux_v
    port map (
            O => \N__36271\,
            I => \N__36263\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__36268\,
            I => buf_dds1_12
        );

    \I__7214\ : Odrv4
    port map (
            O => \N__36263\,
            I => buf_dds1_12
        );

    \I__7213\ : InMux
    port map (
            O => \N__36258\,
            I => \N__36253\
        );

    \I__7212\ : InMux
    port map (
            O => \N__36257\,
            I => \N__36250\
        );

    \I__7211\ : InMux
    port map (
            O => \N__36256\,
            I => \N__36247\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__36253\,
            I => \N__36244\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__36250\,
            I => buf_dds0_12
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__36247\,
            I => buf_dds0_12
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__36244\,
            I => buf_dds0_12
        );

    \I__7206\ : CascadeMux
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__7205\ : InMux
    port map (
            O => \N__36234\,
            I => \N__36231\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__36231\,
            I => \N__36228\
        );

    \I__7203\ : Odrv4
    port map (
            O => \N__36228\,
            I => n8_adj_1566
        );

    \I__7202\ : IoInMux
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__36222\,
            I => \N__36219\
        );

    \I__7200\ : Sp12to4
    port map (
            O => \N__36219\,
            I => \N__36216\
        );

    \I__7199\ : Span12Mux_v
    port map (
            O => \N__36216\,
            I => \N__36211\
        );

    \I__7198\ : InMux
    port map (
            O => \N__36215\,
            I => \N__36208\
        );

    \I__7197\ : InMux
    port map (
            O => \N__36214\,
            I => \N__36205\
        );

    \I__7196\ : Odrv12
    port map (
            O => \N__36211\,
            I => \SELIRNG1\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__36208\,
            I => \SELIRNG1\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__36205\,
            I => \SELIRNG1\
        );

    \I__7193\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36193\
        );

    \I__7192\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36190\
        );

    \I__7191\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36187\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__36193\,
            I => \N__36182\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__36190\,
            I => \N__36182\
        );

    \I__7188\ : InMux
    port map (
            O => \N__36187\,
            I => \N__36179\
        );

    \I__7187\ : Span4Mux_h
    port map (
            O => \N__36182\,
            I => \N__36176\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__36179\,
            I => n14_adj_1546
        );

    \I__7185\ : Odrv4
    port map (
            O => \N__36176\,
            I => n14_adj_1546
        );

    \I__7184\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36167\
        );

    \I__7183\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36162\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__36167\,
            I => \N__36159\
        );

    \I__7181\ : CascadeMux
    port map (
            O => \N__36166\,
            I => \N__36156\
        );

    \I__7180\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36153\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__36162\,
            I => \N__36150\
        );

    \I__7178\ : Span4Mux_v
    port map (
            O => \N__36159\,
            I => \N__36147\
        );

    \I__7177\ : InMux
    port map (
            O => \N__36156\,
            I => \N__36144\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__36153\,
            I => \N__36139\
        );

    \I__7175\ : Span4Mux_v
    port map (
            O => \N__36150\,
            I => \N__36139\
        );

    \I__7174\ : Span4Mux_h
    port map (
            O => \N__36147\,
            I => \N__36136\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__36144\,
            I => n14_adj_1549
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__36139\,
            I => n14_adj_1549
        );

    \I__7171\ : Odrv4
    port map (
            O => \N__36136\,
            I => n14_adj_1549
        );

    \I__7170\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36125\
        );

    \I__7169\ : InMux
    port map (
            O => \N__36128\,
            I => \N__36122\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__36125\,
            I => n8_adj_1562
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__36122\,
            I => n8_adj_1562
        );

    \I__7166\ : CascadeMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__7165\ : CascadeBuf
    port map (
            O => \N__36114\,
            I => \N__36111\
        );

    \I__7164\ : CascadeMux
    port map (
            O => \N__36111\,
            I => \N__36108\
        );

    \I__7163\ : CascadeBuf
    port map (
            O => \N__36108\,
            I => \N__36105\
        );

    \I__7162\ : CascadeMux
    port map (
            O => \N__36105\,
            I => \N__36102\
        );

    \I__7161\ : CascadeBuf
    port map (
            O => \N__36102\,
            I => \N__36099\
        );

    \I__7160\ : CascadeMux
    port map (
            O => \N__36099\,
            I => \N__36096\
        );

    \I__7159\ : CascadeBuf
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__36093\,
            I => \N__36090\
        );

    \I__7157\ : CascadeBuf
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__7156\ : CascadeMux
    port map (
            O => \N__36087\,
            I => \N__36084\
        );

    \I__7155\ : CascadeBuf
    port map (
            O => \N__36084\,
            I => \N__36081\
        );

    \I__7154\ : CascadeMux
    port map (
            O => \N__36081\,
            I => \N__36077\
        );

    \I__7153\ : CascadeMux
    port map (
            O => \N__36080\,
            I => \N__36074\
        );

    \I__7152\ : CascadeBuf
    port map (
            O => \N__36077\,
            I => \N__36071\
        );

    \I__7151\ : CascadeBuf
    port map (
            O => \N__36074\,
            I => \N__36068\
        );

    \I__7150\ : CascadeMux
    port map (
            O => \N__36071\,
            I => \N__36065\
        );

    \I__7149\ : CascadeMux
    port map (
            O => \N__36068\,
            I => \N__36062\
        );

    \I__7148\ : CascadeBuf
    port map (
            O => \N__36065\,
            I => \N__36059\
        );

    \I__7147\ : InMux
    port map (
            O => \N__36062\,
            I => \N__36056\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__36059\,
            I => \N__36053\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__36056\,
            I => \N__36050\
        );

    \I__7144\ : CascadeBuf
    port map (
            O => \N__36053\,
            I => \N__36047\
        );

    \I__7143\ : Span4Mux_h
    port map (
            O => \N__36050\,
            I => \N__36044\
        );

    \I__7142\ : CascadeMux
    port map (
            O => \N__36047\,
            I => \N__36041\
        );

    \I__7141\ : Span4Mux_v
    port map (
            O => \N__36044\,
            I => \N__36038\
        );

    \I__7140\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36035\
        );

    \I__7139\ : Span4Mux_v
    port map (
            O => \N__36038\,
            I => \N__36032\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__36029\
        );

    \I__7137\ : Sp12to4
    port map (
            O => \N__36032\,
            I => \N__36024\
        );

    \I__7136\ : Span12Mux_s11_v
    port map (
            O => \N__36029\,
            I => \N__36024\
        );

    \I__7135\ : Odrv12
    port map (
            O => \N__36024\,
            I => \data_index_9_N_212_6\
        );

    \I__7134\ : InMux
    port map (
            O => \N__36021\,
            I => \N__36018\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__36018\,
            I => n17_adj_1553
        );

    \I__7132\ : IoInMux
    port map (
            O => \N__36015\,
            I => \N__36012\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__36012\,
            I => \N__36009\
        );

    \I__7130\ : Span4Mux_s0_h
    port map (
            O => \N__36009\,
            I => \N__36006\
        );

    \I__7129\ : Span4Mux_v
    port map (
            O => \N__36006\,
            I => \N__36003\
        );

    \I__7128\ : Span4Mux_v
    port map (
            O => \N__36003\,
            I => \N__36000\
        );

    \I__7127\ : Span4Mux_h
    port map (
            O => \N__36000\,
            I => \N__35997\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__35997\,
            I => \N__35993\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35990\
        );

    \I__7124\ : Span4Mux_h
    port map (
            O => \N__35993\,
            I => \N__35984\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__35990\,
            I => \N__35984\
        );

    \I__7122\ : CascadeMux
    port map (
            O => \N__35989\,
            I => \N__35981\
        );

    \I__7121\ : Span4Mux_h
    port map (
            O => \N__35984\,
            I => \N__35978\
        );

    \I__7120\ : InMux
    port map (
            O => \N__35981\,
            I => \N__35975\
        );

    \I__7119\ : Span4Mux_v
    port map (
            O => \N__35978\,
            I => \N__35972\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__35975\,
            I => \AMPV_POW\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__35972\,
            I => \AMPV_POW\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__35967\,
            I => \N__35964\
        );

    \I__7115\ : CascadeBuf
    port map (
            O => \N__35964\,
            I => \N__35961\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__35961\,
            I => \N__35958\
        );

    \I__7113\ : CascadeBuf
    port map (
            O => \N__35958\,
            I => \N__35955\
        );

    \I__7112\ : CascadeMux
    port map (
            O => \N__35955\,
            I => \N__35952\
        );

    \I__7111\ : CascadeBuf
    port map (
            O => \N__35952\,
            I => \N__35949\
        );

    \I__7110\ : CascadeMux
    port map (
            O => \N__35949\,
            I => \N__35946\
        );

    \I__7109\ : CascadeBuf
    port map (
            O => \N__35946\,
            I => \N__35943\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__35943\,
            I => \N__35940\
        );

    \I__7107\ : CascadeBuf
    port map (
            O => \N__35940\,
            I => \N__35937\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__35937\,
            I => \N__35934\
        );

    \I__7105\ : CascadeBuf
    port map (
            O => \N__35934\,
            I => \N__35931\
        );

    \I__7104\ : CascadeMux
    port map (
            O => \N__35931\,
            I => \N__35928\
        );

    \I__7103\ : CascadeBuf
    port map (
            O => \N__35928\,
            I => \N__35925\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__35925\,
            I => \N__35922\
        );

    \I__7101\ : CascadeBuf
    port map (
            O => \N__35922\,
            I => \N__35918\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__35921\,
            I => \N__35915\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__35918\,
            I => \N__35912\
        );

    \I__7098\ : CascadeBuf
    port map (
            O => \N__35915\,
            I => \N__35909\
        );

    \I__7097\ : CascadeBuf
    port map (
            O => \N__35912\,
            I => \N__35906\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__35909\,
            I => \N__35903\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__35906\,
            I => \N__35900\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35897\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35894\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35897\,
            I => \N__35891\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35894\,
            I => \N__35888\
        );

    \I__7090\ : Span12Mux_h
    port map (
            O => \N__35891\,
            I => \N__35883\
        );

    \I__7089\ : Span12Mux_h
    port map (
            O => \N__35888\,
            I => \N__35883\
        );

    \I__7088\ : Odrv12
    port map (
            O => \N__35883\,
            I => \data_index_9_N_212_3\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35877\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35877\,
            I => \N__35867\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__35876\,
            I => \N__35862\
        );

    \I__7084\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35852\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35874\,
            I => \N__35852\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35873\,
            I => \N__35852\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35872\,
            I => \N__35847\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35871\,
            I => \N__35847\
        );

    \I__7079\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35844\
        );

    \I__7078\ : Span12Mux_h
    port map (
            O => \N__35867\,
            I => \N__35841\
        );

    \I__7077\ : InMux
    port map (
            O => \N__35866\,
            I => \N__35834\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35834\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35834\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35829\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35829\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35826\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__35852\,
            I => eis_state_1
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35847\,
            I => eis_state_1
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__35844\,
            I => eis_state_1
        );

    \I__7068\ : Odrv12
    port map (
            O => \N__35841\,
            I => eis_state_1
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__35834\,
            I => eis_state_1
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35829\,
            I => eis_state_1
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__35826\,
            I => eis_state_1
        );

    \I__7064\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35808\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__35808\,
            I => \N__35804\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35807\,
            I => \N__35801\
        );

    \I__7061\ : Span4Mux_v
    port map (
            O => \N__35804\,
            I => \N__35795\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__35801\,
            I => \N__35795\
        );

    \I__7059\ : InMux
    port map (
            O => \N__35800\,
            I => \N__35788\
        );

    \I__7058\ : Sp12to4
    port map (
            O => \N__35795\,
            I => \N__35785\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__35794\,
            I => \N__35778\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35793\,
            I => \N__35768\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35792\,
            I => \N__35768\
        );

    \I__7054\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35768\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__35788\,
            I => \N__35763\
        );

    \I__7052\ : Span12Mux_v
    port map (
            O => \N__35785\,
            I => \N__35763\
        );

    \I__7051\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35752\
        );

    \I__7050\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35752\
        );

    \I__7049\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35752\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35752\
        );

    \I__7047\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35752\
        );

    \I__7046\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35745\
        );

    \I__7045\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35745\
        );

    \I__7044\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35745\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__35768\,
            I => eis_state_2
        );

    \I__7042\ : Odrv12
    port map (
            O => \N__35763\,
            I => eis_state_2
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35752\,
            I => eis_state_2
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__35745\,
            I => eis_state_2
        );

    \I__7039\ : InMux
    port map (
            O => \N__35736\,
            I => \N__35728\
        );

    \I__7038\ : SRMux
    port map (
            O => \N__35735\,
            I => \N__35725\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35734\,
            I => \N__35720\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35733\,
            I => \N__35720\
        );

    \I__7035\ : SRMux
    port map (
            O => \N__35732\,
            I => \N__35717\
        );

    \I__7034\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35714\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__35728\,
            I => \N__35711\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__35725\,
            I => \N__35703\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__35720\,
            I => \N__35698\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35717\,
            I => \N__35698\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35714\,
            I => \N__35695\
        );

    \I__7028\ : Span4Mux_h
    port map (
            O => \N__35711\,
            I => \N__35692\
        );

    \I__7027\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35689\
        );

    \I__7026\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35686\
        );

    \I__7025\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35681\
        );

    \I__7024\ : InMux
    port map (
            O => \N__35707\,
            I => \N__35681\
        );

    \I__7023\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35678\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__35703\,
            I => \N__35675\
        );

    \I__7021\ : Span12Mux_h
    port map (
            O => \N__35698\,
            I => \N__35672\
        );

    \I__7020\ : Span4Mux_v
    port map (
            O => \N__35695\,
            I => \N__35667\
        );

    \I__7019\ : Span4Mux_v
    port map (
            O => \N__35692\,
            I => \N__35667\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__35689\,
            I => \N__35664\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__35686\,
            I => \N__35661\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__35681\,
            I => \N__35658\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35678\,
            I => acadc_rst
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__35675\,
            I => acadc_rst
        );

    \I__7013\ : Odrv12
    port map (
            O => \N__35672\,
            I => acadc_rst
        );

    \I__7012\ : Odrv4
    port map (
            O => \N__35667\,
            I => acadc_rst
        );

    \I__7011\ : Odrv12
    port map (
            O => \N__35664\,
            I => acadc_rst
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__35661\,
            I => acadc_rst
        );

    \I__7009\ : Odrv4
    port map (
            O => \N__35658\,
            I => acadc_rst
        );

    \I__7008\ : InMux
    port map (
            O => \N__35643\,
            I => \N__35640\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__35640\,
            I => n66
        );

    \I__7006\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35634\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__35634\,
            I => \N__35631\
        );

    \I__7004\ : Span4Mux_h
    port map (
            O => \N__35631\,
            I => \N__35626\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35623\
        );

    \I__7002\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35620\
        );

    \I__7001\ : Span4Mux_h
    port map (
            O => \N__35626\,
            I => \N__35617\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__35623\,
            I => \N__35614\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__35620\,
            I => buf_dds1_14
        );

    \I__6998\ : Odrv4
    port map (
            O => \N__35617\,
            I => buf_dds1_14
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__35614\,
            I => buf_dds1_14
        );

    \I__6996\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35604\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35599\
        );

    \I__6994\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35596\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__35602\,
            I => \N__35593\
        );

    \I__6992\ : Span4Mux_v
    port map (
            O => \N__35599\,
            I => \N__35590\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35587\
        );

    \I__6990\ : InMux
    port map (
            O => \N__35593\,
            I => \N__35584\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__35590\,
            I => \N__35581\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__35587\,
            I => \N__35578\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__35584\,
            I => buf_dds1_1
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__35581\,
            I => buf_dds1_1
        );

    \I__6985\ : Odrv4
    port map (
            O => \N__35578\,
            I => buf_dds1_1
        );

    \I__6984\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35562\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35562\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35562\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35562\,
            I => \N__35552\
        );

    \I__6980\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35547\
        );

    \I__6979\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35547\
        );

    \I__6978\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35544\
        );

    \I__6977\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35539\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35539\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__35556\,
            I => \N__35534\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35530\
        );

    \I__6973\ : Span4Mux_v
    port map (
            O => \N__35552\,
            I => \N__35525\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35525\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__35544\,
            I => \N__35520\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35520\
        );

    \I__6969\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35511\
        );

    \I__6968\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35511\
        );

    \I__6967\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35511\
        );

    \I__6966\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35511\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__35530\,
            I => \N__35505\
        );

    \I__6964\ : Span4Mux_v
    port map (
            O => \N__35525\,
            I => \N__35502\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__35520\,
            I => \N__35499\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__35511\,
            I => \N__35496\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35489\
        );

    \I__6960\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35489\
        );

    \I__6959\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35489\
        );

    \I__6958\ : Odrv12
    port map (
            O => \N__35505\,
            I => n12662
        );

    \I__6957\ : Odrv4
    port map (
            O => \N__35502\,
            I => n12662
        );

    \I__6956\ : Odrv4
    port map (
            O => \N__35499\,
            I => n12662
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__35496\,
            I => n12662
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__35489\,
            I => n12662
        );

    \I__6953\ : CascadeMux
    port map (
            O => \N__35478\,
            I => \N__35475\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35472\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__35472\,
            I => \N__35469\
        );

    \I__6950\ : Span4Mux_h
    port map (
            O => \N__35469\,
            I => \N__35466\
        );

    \I__6949\ : Odrv4
    port map (
            O => \N__35466\,
            I => n5_adj_1536
        );

    \I__6948\ : CascadeMux
    port map (
            O => \N__35463\,
            I => \n7_adj_1650_cascade_\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35460\,
            I => \N__35457\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__35457\,
            I => \N__35453\
        );

    \I__6945\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35450\
        );

    \I__6944\ : Span4Mux_v
    port map (
            O => \N__35453\,
            I => \N__35445\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__35450\,
            I => \N__35445\
        );

    \I__6942\ : Odrv4
    port map (
            O => \N__35445\,
            I => n12
        );

    \I__6941\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35439\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__35439\,
            I => \N__35436\
        );

    \I__6939\ : Span4Mux_h
    port map (
            O => \N__35436\,
            I => \N__35433\
        );

    \I__6938\ : Odrv4
    port map (
            O => \N__35433\,
            I => n16_adj_1645
        );

    \I__6937\ : CascadeMux
    port map (
            O => \N__35430\,
            I => \n22641_cascade_\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35424\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35424\,
            I => \N__35420\
        );

    \I__6934\ : CascadeMux
    port map (
            O => \N__35423\,
            I => \N__35417\
        );

    \I__6933\ : Span4Mux_v
    port map (
            O => \N__35420\,
            I => \N__35414\
        );

    \I__6932\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35411\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__35414\,
            I => \N__35408\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__35411\,
            I => data_idxvec_2
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__35408\,
            I => data_idxvec_2
        );

    \I__6928\ : CascadeMux
    port map (
            O => \N__35403\,
            I => \n26_adj_1647_cascade_\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35397\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__35397\,
            I => \N__35394\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__35394\,
            I => \N__35389\
        );

    \I__6924\ : InMux
    port map (
            O => \N__35393\,
            I => \N__35384\
        );

    \I__6923\ : InMux
    port map (
            O => \N__35392\,
            I => \N__35384\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__35389\,
            I => \acadc_skipCount_2\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__35384\,
            I => \acadc_skipCount_2\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__35379\,
            I => \n22383_cascade_\
        );

    \I__6919\ : InMux
    port map (
            O => \N__35376\,
            I => \N__35371\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__35375\,
            I => \N__35368\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__35374\,
            I => \N__35365\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__35371\,
            I => \N__35362\
        );

    \I__6915\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35357\
        );

    \I__6914\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35357\
        );

    \I__6913\ : Odrv12
    port map (
            O => \N__35362\,
            I => req_data_cnt_2
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__35357\,
            I => req_data_cnt_2
        );

    \I__6911\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35349\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__35349\,
            I => n22644
        );

    \I__6909\ : CascadeMux
    port map (
            O => \N__35346\,
            I => \n22386_cascade_\
        );

    \I__6908\ : CascadeMux
    port map (
            O => \N__35343\,
            I => \n30_adj_1648_cascade_\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__35340\,
            I => \N__35337\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35332\
        );

    \I__6905\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35329\
        );

    \I__6904\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35326\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__35332\,
            I => \N__35323\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__35329\,
            I => req_data_cnt_4
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__35326\,
            I => req_data_cnt_4
        );

    \I__6900\ : Odrv4
    port map (
            O => \N__35323\,
            I => req_data_cnt_4
        );

    \I__6899\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35313\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__35313\,
            I => n18_adj_1644
        );

    \I__6897\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35306\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__35309\,
            I => \N__35303\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__35306\,
            I => \N__35300\
        );

    \I__6894\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35296\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__35300\,
            I => \N__35293\
        );

    \I__6892\ : InMux
    port map (
            O => \N__35299\,
            I => \N__35290\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__35296\,
            I => \N__35287\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__35293\,
            I => buf_dds0_13
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__35290\,
            I => buf_dds0_13
        );

    \I__6888\ : Odrv4
    port map (
            O => \N__35287\,
            I => buf_dds0_13
        );

    \I__6887\ : CascadeMux
    port map (
            O => \N__35280\,
            I => \N__35276\
        );

    \I__6886\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35273\
        );

    \I__6885\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35270\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35267\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__35270\,
            I => \N__35264\
        );

    \I__6882\ : Span4Mux_h
    port map (
            O => \N__35267\,
            I => \N__35261\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__35264\,
            I => n9269
        );

    \I__6880\ : Odrv4
    port map (
            O => \N__35261\,
            I => n9269
        );

    \I__6879\ : CascadeMux
    port map (
            O => \N__35256\,
            I => \n12082_cascade_\
        );

    \I__6878\ : InMux
    port map (
            O => \N__35253\,
            I => \N__35250\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__6876\ : Span4Mux_h
    port map (
            O => \N__35247\,
            I => \N__35243\
        );

    \I__6875\ : InMux
    port map (
            O => \N__35246\,
            I => \N__35240\
        );

    \I__6874\ : Span4Mux_h
    port map (
            O => \N__35243\,
            I => \N__35237\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__35240\,
            I => \N__35234\
        );

    \I__6872\ : Span4Mux_v
    port map (
            O => \N__35237\,
            I => \N__35231\
        );

    \I__6871\ : Odrv4
    port map (
            O => \N__35234\,
            I => n14_adj_1573
        );

    \I__6870\ : Odrv4
    port map (
            O => \N__35231\,
            I => n14_adj_1573
        );

    \I__6869\ : SRMux
    port map (
            O => \N__35226\,
            I => \N__35223\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__35223\,
            I => \N__35220\
        );

    \I__6867\ : Span4Mux_v
    port map (
            O => \N__35220\,
            I => \N__35217\
        );

    \I__6866\ : Odrv4
    port map (
            O => \N__35217\,
            I => \comm_spi.data_tx_7__N_817\
        );

    \I__6865\ : CascadeMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__6864\ : InMux
    port map (
            O => \N__35211\,
            I => \N__35207\
        );

    \I__6863\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35203\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__35207\,
            I => \N__35200\
        );

    \I__6861\ : InMux
    port map (
            O => \N__35206\,
            I => \N__35197\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__35203\,
            I => \N__35192\
        );

    \I__6859\ : Span4Mux_v
    port map (
            O => \N__35200\,
            I => \N__35192\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__35197\,
            I => req_data_cnt_10
        );

    \I__6857\ : Odrv4
    port map (
            O => \N__35192\,
            I => req_data_cnt_10
        );

    \I__6856\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35184\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__35184\,
            I => \N__35181\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__35181\,
            I => \N__35178\
        );

    \I__6853\ : Odrv4
    port map (
            O => \N__35178\,
            I => n19_adj_1646
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__35175\,
            I => \N__35172\
        );

    \I__6851\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35169\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__35169\,
            I => \N__35166\
        );

    \I__6849\ : Span4Mux_v
    port map (
            O => \N__35166\,
            I => \N__35163\
        );

    \I__6848\ : Span4Mux_h
    port map (
            O => \N__35163\,
            I => \N__35160\
        );

    \I__6847\ : Sp12to4
    port map (
            O => \N__35160\,
            I => \N__35156\
        );

    \I__6846\ : InMux
    port map (
            O => \N__35159\,
            I => \N__35153\
        );

    \I__6845\ : Odrv12
    port map (
            O => \N__35156\,
            I => \buf_readRTD_2\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__35153\,
            I => \buf_readRTD_2\
        );

    \I__6843\ : InMux
    port map (
            O => \N__35148\,
            I => \N__35145\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__35145\,
            I => \N__35141\
        );

    \I__6841\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35138\
        );

    \I__6840\ : Span4Mux_h
    port map (
            O => \N__35141\,
            I => \N__35135\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__35138\,
            I => secclk_cnt_9
        );

    \I__6838\ : Odrv4
    port map (
            O => \N__35135\,
            I => secclk_cnt_9
        );

    \I__6837\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35126\
        );

    \I__6836\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35123\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__35126\,
            I => \N__35120\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__35123\,
            I => secclk_cnt_17
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__35120\,
            I => secclk_cnt_17
        );

    \I__6832\ : InMux
    port map (
            O => \N__35115\,
            I => \N__35112\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__35112\,
            I => n10
        );

    \I__6830\ : InMux
    port map (
            O => \N__35109\,
            I => \N__35106\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__6828\ : Span4Mux_v
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__6827\ : Span4Mux_h
    port map (
            O => \N__35100\,
            I => \N__35097\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__35097\,
            I => n19_adj_1683
        );

    \I__6825\ : CascadeMux
    port map (
            O => \N__35094\,
            I => \N__35091\
        );

    \I__6824\ : InMux
    port map (
            O => \N__35091\,
            I => \N__35088\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__35088\,
            I => \N__35085\
        );

    \I__6822\ : Span4Mux_h
    port map (
            O => \N__35085\,
            I => \N__35082\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__35082\,
            I => \N__35079\
        );

    \I__6820\ : Odrv4
    port map (
            O => \N__35079\,
            I => n20_adj_1684
        );

    \I__6819\ : InMux
    port map (
            O => \N__35076\,
            I => \N__35073\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__35073\,
            I => \N__35070\
        );

    \I__6817\ : Span4Mux_v
    port map (
            O => \N__35070\,
            I => \N__35066\
        );

    \I__6816\ : CascadeMux
    port map (
            O => \N__35069\,
            I => \N__35063\
        );

    \I__6815\ : Span4Mux_h
    port map (
            O => \N__35066\,
            I => \N__35060\
        );

    \I__6814\ : InMux
    port map (
            O => \N__35063\,
            I => \N__35057\
        );

    \I__6813\ : Odrv4
    port map (
            O => \N__35060\,
            I => buf_adcdata_vdc_11
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__35057\,
            I => buf_adcdata_vdc_11
        );

    \I__6811\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35049\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__35049\,
            I => \N__35046\
        );

    \I__6809\ : Sp12to4
    port map (
            O => \N__35046\,
            I => \N__35041\
        );

    \I__6808\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35038\
        );

    \I__6807\ : InMux
    port map (
            O => \N__35044\,
            I => \N__35035\
        );

    \I__6806\ : Span12Mux_v
    port map (
            O => \N__35041\,
            I => \N__35030\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__35038\,
            I => \N__35030\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__35035\,
            I => buf_adcdata_vac_11
        );

    \I__6803\ : Odrv12
    port map (
            O => \N__35030\,
            I => buf_adcdata_vac_11
        );

    \I__6802\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__35022\,
            I => \N__35018\
        );

    \I__6800\ : InMux
    port map (
            O => \N__35021\,
            I => \N__35015\
        );

    \I__6799\ : Odrv12
    port map (
            O => \N__35018\,
            I => \buf_readRTD_12\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__35015\,
            I => \buf_readRTD_12\
        );

    \I__6797\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35005\
        );

    \I__6796\ : InMux
    port map (
            O => \N__35009\,
            I => \N__35000\
        );

    \I__6795\ : InMux
    port map (
            O => \N__35008\,
            I => \N__35000\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__35005\,
            I => \N__34993\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__35000\,
            I => \N__34993\
        );

    \I__6792\ : CascadeMux
    port map (
            O => \N__34999\,
            I => \N__34990\
        );

    \I__6791\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34987\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__34993\,
            I => \N__34984\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34990\,
            I => \N__34981\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34978\
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__34984\,
            I => \buf_cfgRTD_4\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34981\,
            I => \buf_cfgRTD_4\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__34978\,
            I => \buf_cfgRTD_4\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34968\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__34968\,
            I => \N__34964\
        );

    \I__6782\ : CascadeMux
    port map (
            O => \N__34967\,
            I => \N__34961\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__34964\,
            I => \N__34957\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34954\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34951\
        );

    \I__6778\ : Span4Mux_h
    port map (
            O => \N__34957\,
            I => \N__34948\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__34954\,
            I => buf_dds1_13
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__34951\,
            I => buf_dds1_13
        );

    \I__6775\ : Odrv4
    port map (
            O => \N__34948\,
            I => buf_dds1_13
        );

    \I__6774\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34934\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34940\,
            I => \N__34934\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34931\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__34934\,
            I => \N__34928\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__34931\,
            I => \N__34923\
        );

    \I__6769\ : Span4Mux_v
    port map (
            O => \N__34928\,
            I => \N__34923\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__34920\,
            I => \N__34915\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34919\,
            I => \N__34912\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34918\,
            I => \N__34909\
        );

    \I__6764\ : Odrv4
    port map (
            O => \N__34915\,
            I => \buf_cfgRTD_5\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__34912\,
            I => \buf_cfgRTD_5\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__34909\,
            I => \buf_cfgRTD_5\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34902\,
            I => \N__34899\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34899\,
            I => \N__34896\
        );

    \I__6759\ : Span4Mux_h
    port map (
            O => \N__34896\,
            I => \N__34893\
        );

    \I__6758\ : Span4Mux_h
    port map (
            O => \N__34893\,
            I => \N__34889\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34886\
        );

    \I__6756\ : Odrv4
    port map (
            O => \N__34889\,
            I => \buf_readRTD_13\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__34886\,
            I => \buf_readRTD_13\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34874\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34880\,
            I => \N__34874\
        );

    \I__6752\ : InMux
    port map (
            O => \N__34879\,
            I => \N__34871\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34874\,
            I => req_data_cnt_12
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__34871\,
            I => req_data_cnt_12
        );

    \I__6749\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34863\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34863\,
            I => n22
        );

    \I__6747\ : InMux
    port map (
            O => \N__34860\,
            I => \N__34856\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34859\,
            I => \N__34852\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34856\,
            I => \N__34848\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34845\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__34852\,
            I => \N__34842\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34839\
        );

    \I__6741\ : Span4Mux_v
    port map (
            O => \N__34848\,
            I => \N__34836\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__34845\,
            I => \N__34833\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__34842\,
            I => \N__34830\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34839\,
            I => \N__34827\
        );

    \I__6737\ : Sp12to4
    port map (
            O => \N__34836\,
            I => \N__34822\
        );

    \I__6736\ : Sp12to4
    port map (
            O => \N__34833\,
            I => \N__34822\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__34830\,
            I => \N__34819\
        );

    \I__6734\ : Sp12to4
    port map (
            O => \N__34827\,
            I => \N__34816\
        );

    \I__6733\ : Span12Mux_h
    port map (
            O => \N__34822\,
            I => \N__34813\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__34819\,
            I => n14_adj_1548
        );

    \I__6731\ : Odrv12
    port map (
            O => \N__34816\,
            I => n14_adj_1548
        );

    \I__6730\ : Odrv12
    port map (
            O => \N__34813\,
            I => n14_adj_1548
        );

    \I__6729\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34801\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34805\,
            I => \N__34798\
        );

    \I__6727\ : InMux
    port map (
            O => \N__34804\,
            I => \N__34795\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__34801\,
            I => \comm_spi.n23095\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__34798\,
            I => \comm_spi.n23095\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__34795\,
            I => \comm_spi.n23095\
        );

    \I__6723\ : SRMux
    port map (
            O => \N__34788\,
            I => \N__34785\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__34785\,
            I => \N__34782\
        );

    \I__6721\ : Span4Mux_h
    port map (
            O => \N__34782\,
            I => \N__34779\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__34779\,
            I => \comm_spi.data_tx_7__N_807\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34773\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__34773\,
            I => \N__34770\
        );

    \I__6717\ : Span4Mux_h
    port map (
            O => \N__34770\,
            I => \N__34765\
        );

    \I__6716\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34760\
        );

    \I__6715\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34760\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__34765\,
            I => req_data_cnt_13
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__34760\,
            I => req_data_cnt_13
        );

    \I__6712\ : InMux
    port map (
            O => \N__34755\,
            I => \ADC_VDC.n19924\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34747\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34751\,
            I => \N__34742\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34750\,
            I => \N__34742\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__34747\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__34742\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__6706\ : SRMux
    port map (
            O => \N__34737\,
            I => \N__34734\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__6704\ : Odrv4
    port map (
            O => \N__34731\,
            I => \ADC_VDC.n15273\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__34728\,
            I => \N__34725\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34722\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__34722\,
            I => \N__34719\
        );

    \I__6700\ : Odrv4
    port map (
            O => \N__34719\,
            I => n21_adj_1594
        );

    \I__6699\ : SRMux
    port map (
            O => \N__34716\,
            I => \N__34711\
        );

    \I__6698\ : SRMux
    port map (
            O => \N__34715\,
            I => \N__34708\
        );

    \I__6697\ : SRMux
    port map (
            O => \N__34714\,
            I => \N__34705\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__34711\,
            I => \N__34702\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__34708\,
            I => \N__34697\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34697\
        );

    \I__6693\ : Span4Mux_h
    port map (
            O => \N__34702\,
            I => \N__34694\
        );

    \I__6692\ : Sp12to4
    port map (
            O => \N__34697\,
            I => \N__34690\
        );

    \I__6691\ : Span4Mux_h
    port map (
            O => \N__34694\,
            I => \N__34687\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34693\,
            I => \N__34684\
        );

    \I__6689\ : Odrv12
    port map (
            O => \N__34690\,
            I => n14899
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__34687\,
            I => n14899
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__34684\,
            I => n14899
        );

    \I__6686\ : IoInMux
    port map (
            O => \N__34677\,
            I => \N__34674\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34674\,
            I => \N__34671\
        );

    \I__6684\ : IoSpan4Mux
    port map (
            O => \N__34671\,
            I => \N__34668\
        );

    \I__6683\ : Span4Mux_s3_v
    port map (
            O => \N__34668\,
            I => \N__34665\
        );

    \I__6682\ : Sp12to4
    port map (
            O => \N__34665\,
            I => \N__34661\
        );

    \I__6681\ : InMux
    port map (
            O => \N__34664\,
            I => \N__34658\
        );

    \I__6680\ : Span12Mux_h
    port map (
            O => \N__34661\,
            I => \N__34655\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34658\,
            I => \N__34652\
        );

    \I__6678\ : Odrv12
    port map (
            O => \N__34655\,
            I => \TEST_LED\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__34652\,
            I => \TEST_LED\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34647\,
            I => \N__34644\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__34644\,
            I => \N__34640\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34643\,
            I => \N__34637\
        );

    \I__6673\ : Span4Mux_h
    port map (
            O => \N__34640\,
            I => \N__34634\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__34637\,
            I => secclk_cnt_15
        );

    \I__6671\ : Odrv4
    port map (
            O => \N__34634\,
            I => secclk_cnt_15
        );

    \I__6670\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34626\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__34626\,
            I => \N__34622\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34619\
        );

    \I__6667\ : Span4Mux_v
    port map (
            O => \N__34622\,
            I => \N__34616\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__34619\,
            I => secclk_cnt_8
        );

    \I__6665\ : Odrv4
    port map (
            O => \N__34616\,
            I => secclk_cnt_8
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__34611\,
            I => \N__34607\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34610\,
            I => \N__34604\
        );

    \I__6662\ : InMux
    port map (
            O => \N__34607\,
            I => \N__34601\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34596\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__34601\,
            I => \N__34596\
        );

    \I__6659\ : Odrv4
    port map (
            O => \N__34596\,
            I => secclk_cnt_1
        );

    \I__6658\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34589\
        );

    \I__6657\ : InMux
    port map (
            O => \N__34592\,
            I => \N__34586\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34583\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34586\,
            I => secclk_cnt_5
        );

    \I__6654\ : Odrv4
    port map (
            O => \N__34583\,
            I => secclk_cnt_5
        );

    \I__6653\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__34575\,
            I => n25
        );

    \I__6651\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34568\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34565\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__34568\,
            I => \N__34562\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34557\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__34562\,
            I => \N__34557\
        );

    \I__6646\ : Odrv4
    port map (
            O => \N__34557\,
            I => secclk_cnt_18
        );

    \I__6645\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34550\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34547\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__34550\,
            I => \N__34542\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__34547\,
            I => \N__34542\
        );

    \I__6641\ : Odrv4
    port map (
            O => \N__34542\,
            I => secclk_cnt_0
        );

    \I__6640\ : CascadeMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__6639\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34533\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__34533\,
            I => \N__34529\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34526\
        );

    \I__6636\ : Span4Mux_h
    port map (
            O => \N__34529\,
            I => \N__34523\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__34526\,
            I => secclk_cnt_11
        );

    \I__6634\ : Odrv4
    port map (
            O => \N__34523\,
            I => secclk_cnt_11
        );

    \I__6633\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34514\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34511\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__34514\,
            I => \N__34508\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__34511\,
            I => secclk_cnt_4
        );

    \I__6629\ : Odrv12
    port map (
            O => \N__34508\,
            I => secclk_cnt_4
        );

    \I__6628\ : CascadeMux
    port map (
            O => \N__34503\,
            I => \N__34500\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34497\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__34497\,
            I => n28_adj_1554
        );

    \I__6625\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34491\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__34491\,
            I => \N__34488\
        );

    \I__6623\ : Span4Mux_h
    port map (
            O => \N__34488\,
            I => \N__34484\
        );

    \I__6622\ : CascadeMux
    port map (
            O => \N__34487\,
            I => \N__34481\
        );

    \I__6621\ : Span4Mux_v
    port map (
            O => \N__34484\,
            I => \N__34477\
        );

    \I__6620\ : InMux
    port map (
            O => \N__34481\,
            I => \N__34474\
        );

    \I__6619\ : InMux
    port map (
            O => \N__34480\,
            I => \N__34471\
        );

    \I__6618\ : Span4Mux_h
    port map (
            O => \N__34477\,
            I => \N__34466\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34474\,
            I => \N__34466\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__34471\,
            I => req_data_cnt_15
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__34466\,
            I => req_data_cnt_15
        );

    \I__6614\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34458\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__34458\,
            I => n24
        );

    \I__6612\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34452\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__34452\,
            I => \comm_spi.n14822\
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__34449\,
            I => \comm_spi.n23089_cascade_\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__34443\,
            I => \comm_spi.n14823\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__34440\,
            I => \N__34437\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34433\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__34436\,
            I => \N__34430\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__34433\,
            I => \N__34426\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34423\
        );

    \I__6602\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34419\
        );

    \I__6601\ : Span4Mux_v
    port map (
            O => \N__34426\,
            I => \N__34414\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__34423\,
            I => \N__34414\
        );

    \I__6599\ : InMux
    port map (
            O => \N__34422\,
            I => \N__34411\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__34419\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__34414\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__34411\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6595\ : InMux
    port map (
            O => \N__34404\,
            I => \bfn_13_6_0_\
        );

    \I__6594\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34398\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__34398\,
            I => \N__34394\
        );

    \I__6592\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34390\
        );

    \I__6591\ : Span4Mux_h
    port map (
            O => \N__34394\,
            I => \N__34387\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34393\,
            I => \N__34384\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34390\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__34387\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34384\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6586\ : InMux
    port map (
            O => \N__34377\,
            I => \ADC_VDC.n19918\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34370\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34366\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__34370\,
            I => \N__34363\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34360\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__34366\,
            I => \N__34354\
        );

    \I__6580\ : Span4Mux_v
    port map (
            O => \N__34363\,
            I => \N__34354\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__34360\,
            I => \N__34351\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34348\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__34354\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__34351\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34348\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6574\ : InMux
    port map (
            O => \N__34341\,
            I => \ADC_VDC.n19919\
        );

    \I__6573\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34334\
        );

    \I__6572\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34330\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34327\
        );

    \I__6570\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34323\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34318\
        );

    \I__6568\ : Span4Mux_v
    port map (
            O => \N__34327\,
            I => \N__34318\
        );

    \I__6567\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34315\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__34323\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__34318\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__34315\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6563\ : InMux
    port map (
            O => \N__34308\,
            I => \ADC_VDC.n19920\
        );

    \I__6562\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__34302\,
            I => \N__34298\
        );

    \I__6560\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34293\
        );

    \I__6559\ : Span4Mux_h
    port map (
            O => \N__34298\,
            I => \N__34290\
        );

    \I__6558\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34285\
        );

    \I__6557\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34285\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__34293\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__6555\ : Odrv4
    port map (
            O => \N__34290\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__34285\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__6553\ : InMux
    port map (
            O => \N__34278\,
            I => \ADC_VDC.n19921\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__34275\,
            I => \N__34270\
        );

    \I__6551\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34267\
        );

    \I__6550\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34262\
        );

    \I__6549\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34262\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__34267\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__34262\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__6546\ : InMux
    port map (
            O => \N__34257\,
            I => \ADC_VDC.n19922\
        );

    \I__6545\ : InMux
    port map (
            O => \N__34254\,
            I => \N__34249\
        );

    \I__6544\ : InMux
    port map (
            O => \N__34253\,
            I => \N__34244\
        );

    \I__6543\ : InMux
    port map (
            O => \N__34252\,
            I => \N__34244\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__34249\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__34244\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__6540\ : InMux
    port map (
            O => \N__34239\,
            I => \ADC_VDC.n19923\
        );

    \I__6539\ : CascadeMux
    port map (
            O => \N__34236\,
            I => \N__34233\
        );

    \I__6538\ : CascadeBuf
    port map (
            O => \N__34233\,
            I => \N__34230\
        );

    \I__6537\ : CascadeMux
    port map (
            O => \N__34230\,
            I => \N__34227\
        );

    \I__6536\ : CascadeBuf
    port map (
            O => \N__34227\,
            I => \N__34224\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__6534\ : CascadeBuf
    port map (
            O => \N__34221\,
            I => \N__34218\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__34218\,
            I => \N__34215\
        );

    \I__6532\ : CascadeBuf
    port map (
            O => \N__34215\,
            I => \N__34212\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__34212\,
            I => \N__34209\
        );

    \I__6530\ : CascadeBuf
    port map (
            O => \N__34209\,
            I => \N__34206\
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__34206\,
            I => \N__34203\
        );

    \I__6528\ : CascadeBuf
    port map (
            O => \N__34203\,
            I => \N__34200\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__34200\,
            I => \N__34197\
        );

    \I__6526\ : CascadeBuf
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__6525\ : CascadeMux
    port map (
            O => \N__34194\,
            I => \N__34190\
        );

    \I__6524\ : CascadeMux
    port map (
            O => \N__34193\,
            I => \N__34187\
        );

    \I__6523\ : CascadeBuf
    port map (
            O => \N__34190\,
            I => \N__34184\
        );

    \I__6522\ : CascadeBuf
    port map (
            O => \N__34187\,
            I => \N__34181\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__34184\,
            I => \N__34178\
        );

    \I__6520\ : CascadeMux
    port map (
            O => \N__34181\,
            I => \N__34175\
        );

    \I__6519\ : CascadeBuf
    port map (
            O => \N__34178\,
            I => \N__34172\
        );

    \I__6518\ : InMux
    port map (
            O => \N__34175\,
            I => \N__34169\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__34172\,
            I => \N__34166\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__34169\,
            I => \N__34163\
        );

    \I__6515\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34160\
        );

    \I__6514\ : Span4Mux_h
    port map (
            O => \N__34163\,
            I => \N__34157\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__34160\,
            I => \N__34154\
        );

    \I__6512\ : Sp12to4
    port map (
            O => \N__34157\,
            I => \N__34150\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__34154\,
            I => \N__34147\
        );

    \I__6510\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34144\
        );

    \I__6509\ : Span12Mux_v
    port map (
            O => \N__34150\,
            I => \N__34141\
        );

    \I__6508\ : Sp12to4
    port map (
            O => \N__34147\,
            I => \N__34138\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__34144\,
            I => data_count_6
        );

    \I__6506\ : Odrv12
    port map (
            O => \N__34141\,
            I => data_count_6
        );

    \I__6505\ : Odrv12
    port map (
            O => \N__34138\,
            I => data_count_6
        );

    \I__6504\ : InMux
    port map (
            O => \N__34131\,
            I => n19770
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__34128\,
            I => \N__34125\
        );

    \I__6502\ : CascadeBuf
    port map (
            O => \N__34125\,
            I => \N__34122\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__34122\,
            I => \N__34119\
        );

    \I__6500\ : CascadeBuf
    port map (
            O => \N__34119\,
            I => \N__34116\
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__34116\,
            I => \N__34113\
        );

    \I__6498\ : CascadeBuf
    port map (
            O => \N__34113\,
            I => \N__34110\
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__34110\,
            I => \N__34107\
        );

    \I__6496\ : CascadeBuf
    port map (
            O => \N__34107\,
            I => \N__34104\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__34104\,
            I => \N__34101\
        );

    \I__6494\ : CascadeBuf
    port map (
            O => \N__34101\,
            I => \N__34098\
        );

    \I__6493\ : CascadeMux
    port map (
            O => \N__34098\,
            I => \N__34095\
        );

    \I__6492\ : CascadeBuf
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__34092\,
            I => \N__34088\
        );

    \I__6490\ : CascadeMux
    port map (
            O => \N__34091\,
            I => \N__34085\
        );

    \I__6489\ : CascadeBuf
    port map (
            O => \N__34088\,
            I => \N__34082\
        );

    \I__6488\ : CascadeBuf
    port map (
            O => \N__34085\,
            I => \N__34079\
        );

    \I__6487\ : CascadeMux
    port map (
            O => \N__34082\,
            I => \N__34076\
        );

    \I__6486\ : CascadeMux
    port map (
            O => \N__34079\,
            I => \N__34073\
        );

    \I__6485\ : CascadeBuf
    port map (
            O => \N__34076\,
            I => \N__34070\
        );

    \I__6484\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34067\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__34070\,
            I => \N__34064\
        );

    \I__6482\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__34061\
        );

    \I__6481\ : CascadeBuf
    port map (
            O => \N__34064\,
            I => \N__34058\
        );

    \I__6480\ : Span4Mux_h
    port map (
            O => \N__34061\,
            I => \N__34055\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__34058\,
            I => \N__34052\
        );

    \I__6478\ : Span4Mux_h
    port map (
            O => \N__34055\,
            I => \N__34049\
        );

    \I__6477\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34046\
        );

    \I__6476\ : Sp12to4
    port map (
            O => \N__34049\,
            I => \N__34042\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__34039\
        );

    \I__6474\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34036\
        );

    \I__6473\ : Span12Mux_v
    port map (
            O => \N__34042\,
            I => \N__34033\
        );

    \I__6472\ : Span12Mux_s8_v
    port map (
            O => \N__34039\,
            I => \N__34030\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__34036\,
            I => data_count_7
        );

    \I__6470\ : Odrv12
    port map (
            O => \N__34033\,
            I => data_count_7
        );

    \I__6469\ : Odrv12
    port map (
            O => \N__34030\,
            I => data_count_7
        );

    \I__6468\ : InMux
    port map (
            O => \N__34023\,
            I => n19771
        );

    \I__6467\ : CascadeMux
    port map (
            O => \N__34020\,
            I => \N__34017\
        );

    \I__6466\ : CascadeBuf
    port map (
            O => \N__34017\,
            I => \N__34014\
        );

    \I__6465\ : CascadeMux
    port map (
            O => \N__34014\,
            I => \N__34011\
        );

    \I__6464\ : CascadeBuf
    port map (
            O => \N__34011\,
            I => \N__34008\
        );

    \I__6463\ : CascadeMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__6462\ : CascadeBuf
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__6461\ : CascadeMux
    port map (
            O => \N__34002\,
            I => \N__33999\
        );

    \I__6460\ : CascadeBuf
    port map (
            O => \N__33999\,
            I => \N__33996\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__33996\,
            I => \N__33993\
        );

    \I__6458\ : CascadeBuf
    port map (
            O => \N__33993\,
            I => \N__33990\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__33990\,
            I => \N__33987\
        );

    \I__6456\ : CascadeBuf
    port map (
            O => \N__33987\,
            I => \N__33984\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__6454\ : CascadeBuf
    port map (
            O => \N__33981\,
            I => \N__33978\
        );

    \I__6453\ : CascadeMux
    port map (
            O => \N__33978\,
            I => \N__33974\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__33977\,
            I => \N__33971\
        );

    \I__6451\ : CascadeBuf
    port map (
            O => \N__33974\,
            I => \N__33968\
        );

    \I__6450\ : CascadeBuf
    port map (
            O => \N__33971\,
            I => \N__33965\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__33968\,
            I => \N__33962\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__33965\,
            I => \N__33959\
        );

    \I__6447\ : CascadeBuf
    port map (
            O => \N__33962\,
            I => \N__33956\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33953\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__33956\,
            I => \N__33950\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__33953\,
            I => \N__33947\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33950\,
            I => \N__33944\
        );

    \I__6442\ : Span4Mux_v
    port map (
            O => \N__33947\,
            I => \N__33941\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__33944\,
            I => \N__33938\
        );

    \I__6440\ : Sp12to4
    port map (
            O => \N__33941\,
            I => \N__33934\
        );

    \I__6439\ : Span4Mux_v
    port map (
            O => \N__33938\,
            I => \N__33931\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33928\
        );

    \I__6437\ : Span12Mux_h
    port map (
            O => \N__33934\,
            I => \N__33925\
        );

    \I__6436\ : Sp12to4
    port map (
            O => \N__33931\,
            I => \N__33922\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__33928\,
            I => data_count_8
        );

    \I__6434\ : Odrv12
    port map (
            O => \N__33925\,
            I => data_count_8
        );

    \I__6433\ : Odrv12
    port map (
            O => \N__33922\,
            I => data_count_8
        );

    \I__6432\ : InMux
    port map (
            O => \N__33915\,
            I => \bfn_12_19_0_\
        );

    \I__6431\ : InMux
    port map (
            O => \N__33912\,
            I => n19773
        );

    \I__6430\ : CascadeMux
    port map (
            O => \N__33909\,
            I => \N__33906\
        );

    \I__6429\ : CascadeBuf
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__6428\ : CascadeMux
    port map (
            O => \N__33903\,
            I => \N__33900\
        );

    \I__6427\ : CascadeBuf
    port map (
            O => \N__33900\,
            I => \N__33897\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__33897\,
            I => \N__33894\
        );

    \I__6425\ : CascadeBuf
    port map (
            O => \N__33894\,
            I => \N__33891\
        );

    \I__6424\ : CascadeMux
    port map (
            O => \N__33891\,
            I => \N__33888\
        );

    \I__6423\ : CascadeBuf
    port map (
            O => \N__33888\,
            I => \N__33885\
        );

    \I__6422\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33882\
        );

    \I__6421\ : CascadeBuf
    port map (
            O => \N__33882\,
            I => \N__33879\
        );

    \I__6420\ : CascadeMux
    port map (
            O => \N__33879\,
            I => \N__33876\
        );

    \I__6419\ : CascadeBuf
    port map (
            O => \N__33876\,
            I => \N__33873\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__33873\,
            I => \N__33870\
        );

    \I__6417\ : CascadeBuf
    port map (
            O => \N__33870\,
            I => \N__33867\
        );

    \I__6416\ : CascadeMux
    port map (
            O => \N__33867\,
            I => \N__33864\
        );

    \I__6415\ : CascadeBuf
    port map (
            O => \N__33864\,
            I => \N__33860\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__33863\,
            I => \N__33857\
        );

    \I__6413\ : CascadeMux
    port map (
            O => \N__33860\,
            I => \N__33854\
        );

    \I__6412\ : CascadeBuf
    port map (
            O => \N__33857\,
            I => \N__33851\
        );

    \I__6411\ : CascadeBuf
    port map (
            O => \N__33854\,
            I => \N__33848\
        );

    \I__6410\ : CascadeMux
    port map (
            O => \N__33851\,
            I => \N__33845\
        );

    \I__6409\ : CascadeMux
    port map (
            O => \N__33848\,
            I => \N__33842\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33839\
        );

    \I__6407\ : InMux
    port map (
            O => \N__33842\,
            I => \N__33836\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33839\,
            I => \N__33832\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__33836\,
            I => \N__33829\
        );

    \I__6404\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33826\
        );

    \I__6403\ : Span12Mux_h
    port map (
            O => \N__33832\,
            I => \N__33821\
        );

    \I__6402\ : Span12Mux_h
    port map (
            O => \N__33829\,
            I => \N__33821\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__33826\,
            I => data_count_9
        );

    \I__6400\ : Odrv12
    port map (
            O => \N__33821\,
            I => data_count_9
        );

    \I__6399\ : InMux
    port map (
            O => \N__33816\,
            I => \N__33813\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__33813\,
            I => \comm_spi.n23089\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33807\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33807\,
            I => \N__33804\
        );

    \I__6395\ : Span4Mux_v
    port map (
            O => \N__33804\,
            I => \N__33800\
        );

    \I__6394\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33797\
        );

    \I__6393\ : Span4Mux_h
    port map (
            O => \N__33800\,
            I => \N__33791\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33797\,
            I => \N__33791\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33788\
        );

    \I__6390\ : Odrv4
    port map (
            O => \N__33791\,
            I => cmd_rdadctmp_16
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33788\,
            I => cmd_rdadctmp_16
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__33783\,
            I => \N__33780\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33777\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33773\
        );

    \I__6385\ : CascadeMux
    port map (
            O => \N__33776\,
            I => \N__33769\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__33773\,
            I => \N__33766\
        );

    \I__6383\ : InMux
    port map (
            O => \N__33772\,
            I => \N__33761\
        );

    \I__6382\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33761\
        );

    \I__6381\ : Odrv4
    port map (
            O => \N__33766\,
            I => cmd_rdadctmp_17
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__33761\,
            I => cmd_rdadctmp_17
        );

    \I__6379\ : CascadeMux
    port map (
            O => \N__33756\,
            I => \N__33753\
        );

    \I__6378\ : CascadeBuf
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__6377\ : CascadeMux
    port map (
            O => \N__33750\,
            I => \N__33747\
        );

    \I__6376\ : CascadeBuf
    port map (
            O => \N__33747\,
            I => \N__33744\
        );

    \I__6375\ : CascadeMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__6374\ : CascadeBuf
    port map (
            O => \N__33741\,
            I => \N__33738\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__6372\ : CascadeBuf
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__6371\ : CascadeMux
    port map (
            O => \N__33732\,
            I => \N__33729\
        );

    \I__6370\ : CascadeBuf
    port map (
            O => \N__33729\,
            I => \N__33726\
        );

    \I__6369\ : CascadeMux
    port map (
            O => \N__33726\,
            I => \N__33723\
        );

    \I__6368\ : CascadeBuf
    port map (
            O => \N__33723\,
            I => \N__33720\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__33720\,
            I => \N__33717\
        );

    \I__6366\ : CascadeBuf
    port map (
            O => \N__33717\,
            I => \N__33714\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__33714\,
            I => \N__33710\
        );

    \I__6364\ : CascadeMux
    port map (
            O => \N__33713\,
            I => \N__33707\
        );

    \I__6363\ : CascadeBuf
    port map (
            O => \N__33710\,
            I => \N__33704\
        );

    \I__6362\ : CascadeBuf
    port map (
            O => \N__33707\,
            I => \N__33701\
        );

    \I__6361\ : CascadeMux
    port map (
            O => \N__33704\,
            I => \N__33698\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \N__33695\
        );

    \I__6359\ : CascadeBuf
    port map (
            O => \N__33698\,
            I => \N__33692\
        );

    \I__6358\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33689\
        );

    \I__6357\ : CascadeMux
    port map (
            O => \N__33692\,
            I => \N__33686\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33689\,
            I => \N__33683\
        );

    \I__6355\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33680\
        );

    \I__6354\ : Span4Mux_h
    port map (
            O => \N__33683\,
            I => \N__33677\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__33680\,
            I => \N__33674\
        );

    \I__6352\ : Sp12to4
    port map (
            O => \N__33677\,
            I => \N__33670\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__33674\,
            I => \N__33667\
        );

    \I__6350\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33664\
        );

    \I__6349\ : Span12Mux_v
    port map (
            O => \N__33670\,
            I => \N__33659\
        );

    \I__6348\ : Sp12to4
    port map (
            O => \N__33667\,
            I => \N__33659\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__33664\,
            I => data_count_0
        );

    \I__6346\ : Odrv12
    port map (
            O => \N__33659\,
            I => data_count_0
        );

    \I__6345\ : CascadeMux
    port map (
            O => \N__33654\,
            I => \N__33651\
        );

    \I__6344\ : CascadeBuf
    port map (
            O => \N__33651\,
            I => \N__33648\
        );

    \I__6343\ : CascadeMux
    port map (
            O => \N__33648\,
            I => \N__33645\
        );

    \I__6342\ : CascadeBuf
    port map (
            O => \N__33645\,
            I => \N__33642\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__33642\,
            I => \N__33639\
        );

    \I__6340\ : CascadeBuf
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__33636\,
            I => \N__33633\
        );

    \I__6338\ : CascadeBuf
    port map (
            O => \N__33633\,
            I => \N__33630\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__6336\ : CascadeBuf
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__33624\,
            I => \N__33621\
        );

    \I__6334\ : CascadeBuf
    port map (
            O => \N__33621\,
            I => \N__33618\
        );

    \I__6333\ : CascadeMux
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__6332\ : CascadeBuf
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__33612\,
            I => \N__33608\
        );

    \I__6330\ : CascadeMux
    port map (
            O => \N__33611\,
            I => \N__33605\
        );

    \I__6329\ : CascadeBuf
    port map (
            O => \N__33608\,
            I => \N__33602\
        );

    \I__6328\ : CascadeBuf
    port map (
            O => \N__33605\,
            I => \N__33599\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__33602\,
            I => \N__33596\
        );

    \I__6326\ : CascadeMux
    port map (
            O => \N__33599\,
            I => \N__33593\
        );

    \I__6325\ : CascadeBuf
    port map (
            O => \N__33596\,
            I => \N__33590\
        );

    \I__6324\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33587\
        );

    \I__6323\ : CascadeMux
    port map (
            O => \N__33590\,
            I => \N__33584\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__33587\,
            I => \N__33581\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33584\,
            I => \N__33578\
        );

    \I__6320\ : Span4Mux_v
    port map (
            O => \N__33581\,
            I => \N__33575\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__33578\,
            I => \N__33572\
        );

    \I__6318\ : Sp12to4
    port map (
            O => \N__33575\,
            I => \N__33568\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__33572\,
            I => \N__33565\
        );

    \I__6316\ : InMux
    port map (
            O => \N__33571\,
            I => \N__33562\
        );

    \I__6315\ : Span12Mux_h
    port map (
            O => \N__33568\,
            I => \N__33559\
        );

    \I__6314\ : Sp12to4
    port map (
            O => \N__33565\,
            I => \N__33556\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__33562\,
            I => data_count_1
        );

    \I__6312\ : Odrv12
    port map (
            O => \N__33559\,
            I => data_count_1
        );

    \I__6311\ : Odrv12
    port map (
            O => \N__33556\,
            I => data_count_1
        );

    \I__6310\ : InMux
    port map (
            O => \N__33549\,
            I => n19765
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__33546\,
            I => \N__33543\
        );

    \I__6308\ : CascadeBuf
    port map (
            O => \N__33543\,
            I => \N__33540\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__33540\,
            I => \N__33537\
        );

    \I__6306\ : CascadeBuf
    port map (
            O => \N__33537\,
            I => \N__33534\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__6304\ : CascadeBuf
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6303\ : CascadeMux
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__6302\ : CascadeBuf
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__6300\ : CascadeBuf
    port map (
            O => \N__33519\,
            I => \N__33516\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__6298\ : CascadeBuf
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__6297\ : CascadeMux
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__6296\ : CascadeBuf
    port map (
            O => \N__33507\,
            I => \N__33504\
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__6294\ : CascadeBuf
    port map (
            O => \N__33501\,
            I => \N__33497\
        );

    \I__6293\ : CascadeMux
    port map (
            O => \N__33500\,
            I => \N__33494\
        );

    \I__6292\ : CascadeMux
    port map (
            O => \N__33497\,
            I => \N__33491\
        );

    \I__6291\ : CascadeBuf
    port map (
            O => \N__33494\,
            I => \N__33488\
        );

    \I__6290\ : CascadeBuf
    port map (
            O => \N__33491\,
            I => \N__33485\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__33488\,
            I => \N__33482\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__33485\,
            I => \N__33479\
        );

    \I__6287\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33476\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33479\,
            I => \N__33473\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__33476\,
            I => \N__33470\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33473\,
            I => \N__33467\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__33470\,
            I => \N__33464\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__33467\,
            I => \N__33461\
        );

    \I__6281\ : Sp12to4
    port map (
            O => \N__33464\,
            I => \N__33457\
        );

    \I__6280\ : Span4Mux_h
    port map (
            O => \N__33461\,
            I => \N__33454\
        );

    \I__6279\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33451\
        );

    \I__6278\ : Span12Mux_v
    port map (
            O => \N__33457\,
            I => \N__33448\
        );

    \I__6277\ : Span4Mux_h
    port map (
            O => \N__33454\,
            I => \N__33445\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__33451\,
            I => data_count_2
        );

    \I__6275\ : Odrv12
    port map (
            O => \N__33448\,
            I => data_count_2
        );

    \I__6274\ : Odrv4
    port map (
            O => \N__33445\,
            I => data_count_2
        );

    \I__6273\ : InMux
    port map (
            O => \N__33438\,
            I => n19766
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__33435\,
            I => \N__33432\
        );

    \I__6271\ : CascadeBuf
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__33429\,
            I => \N__33426\
        );

    \I__6269\ : CascadeBuf
    port map (
            O => \N__33426\,
            I => \N__33423\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__33423\,
            I => \N__33420\
        );

    \I__6267\ : CascadeBuf
    port map (
            O => \N__33420\,
            I => \N__33417\
        );

    \I__6266\ : CascadeMux
    port map (
            O => \N__33417\,
            I => \N__33414\
        );

    \I__6265\ : CascadeBuf
    port map (
            O => \N__33414\,
            I => \N__33411\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__33411\,
            I => \N__33408\
        );

    \I__6263\ : CascadeBuf
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__6262\ : CascadeMux
    port map (
            O => \N__33405\,
            I => \N__33402\
        );

    \I__6261\ : CascadeBuf
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__6260\ : CascadeMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__6259\ : CascadeBuf
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__6258\ : CascadeMux
    port map (
            O => \N__33393\,
            I => \N__33390\
        );

    \I__6257\ : CascadeBuf
    port map (
            O => \N__33390\,
            I => \N__33386\
        );

    \I__6256\ : CascadeMux
    port map (
            O => \N__33389\,
            I => \N__33383\
        );

    \I__6255\ : CascadeMux
    port map (
            O => \N__33386\,
            I => \N__33380\
        );

    \I__6254\ : CascadeBuf
    port map (
            O => \N__33383\,
            I => \N__33377\
        );

    \I__6253\ : CascadeBuf
    port map (
            O => \N__33380\,
            I => \N__33374\
        );

    \I__6252\ : CascadeMux
    port map (
            O => \N__33377\,
            I => \N__33371\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__33374\,
            I => \N__33368\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33365\
        );

    \I__6249\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33362\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__33365\,
            I => \N__33359\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__33362\,
            I => \N__33356\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__33359\,
            I => \N__33353\
        );

    \I__6245\ : Span4Mux_v
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__33353\,
            I => \N__33346\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__33350\,
            I => \N__33343\
        );

    \I__6242\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33340\
        );

    \I__6241\ : Sp12to4
    port map (
            O => \N__33346\,
            I => \N__33337\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__33343\,
            I => \N__33334\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__33340\,
            I => data_count_3
        );

    \I__6238\ : Odrv12
    port map (
            O => \N__33337\,
            I => data_count_3
        );

    \I__6237\ : Odrv4
    port map (
            O => \N__33334\,
            I => data_count_3
        );

    \I__6236\ : InMux
    port map (
            O => \N__33327\,
            I => n19767
        );

    \I__6235\ : CascadeMux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__6234\ : CascadeBuf
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__6233\ : CascadeMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__6232\ : CascadeBuf
    port map (
            O => \N__33315\,
            I => \N__33312\
        );

    \I__6231\ : CascadeMux
    port map (
            O => \N__33312\,
            I => \N__33309\
        );

    \I__6230\ : CascadeBuf
    port map (
            O => \N__33309\,
            I => \N__33306\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__33306\,
            I => \N__33303\
        );

    \I__6228\ : CascadeBuf
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__6227\ : CascadeMux
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__6226\ : CascadeBuf
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__33294\,
            I => \N__33291\
        );

    \I__6224\ : CascadeBuf
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__33288\,
            I => \N__33285\
        );

    \I__6222\ : CascadeBuf
    port map (
            O => \N__33285\,
            I => \N__33282\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__6220\ : CascadeBuf
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__6219\ : CascadeMux
    port map (
            O => \N__33276\,
            I => \N__33272\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__33275\,
            I => \N__33269\
        );

    \I__6217\ : CascadeBuf
    port map (
            O => \N__33272\,
            I => \N__33266\
        );

    \I__6216\ : CascadeBuf
    port map (
            O => \N__33269\,
            I => \N__33263\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__33266\,
            I => \N__33260\
        );

    \I__6214\ : CascadeMux
    port map (
            O => \N__33263\,
            I => \N__33257\
        );

    \I__6213\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33254\
        );

    \I__6212\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33251\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33248\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__33251\,
            I => \N__33244\
        );

    \I__6209\ : Span4Mux_v
    port map (
            O => \N__33248\,
            I => \N__33241\
        );

    \I__6208\ : InMux
    port map (
            O => \N__33247\,
            I => \N__33238\
        );

    \I__6207\ : Span12Mux_v
    port map (
            O => \N__33244\,
            I => \N__33235\
        );

    \I__6206\ : Sp12to4
    port map (
            O => \N__33241\,
            I => \N__33232\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__33238\,
            I => data_count_4
        );

    \I__6204\ : Odrv12
    port map (
            O => \N__33235\,
            I => data_count_4
        );

    \I__6203\ : Odrv12
    port map (
            O => \N__33232\,
            I => data_count_4
        );

    \I__6202\ : InMux
    port map (
            O => \N__33225\,
            I => n19768
        );

    \I__6201\ : CascadeMux
    port map (
            O => \N__33222\,
            I => \N__33219\
        );

    \I__6200\ : CascadeBuf
    port map (
            O => \N__33219\,
            I => \N__33216\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__33216\,
            I => \N__33213\
        );

    \I__6198\ : CascadeBuf
    port map (
            O => \N__33213\,
            I => \N__33210\
        );

    \I__6197\ : CascadeMux
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__6196\ : CascadeBuf
    port map (
            O => \N__33207\,
            I => \N__33204\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__6194\ : CascadeBuf
    port map (
            O => \N__33201\,
            I => \N__33198\
        );

    \I__6193\ : CascadeMux
    port map (
            O => \N__33198\,
            I => \N__33195\
        );

    \I__6192\ : CascadeBuf
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__6191\ : CascadeMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__6190\ : CascadeBuf
    port map (
            O => \N__33189\,
            I => \N__33186\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__33186\,
            I => \N__33183\
        );

    \I__6188\ : CascadeBuf
    port map (
            O => \N__33183\,
            I => \N__33179\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__33182\,
            I => \N__33176\
        );

    \I__6186\ : CascadeMux
    port map (
            O => \N__33179\,
            I => \N__33173\
        );

    \I__6185\ : CascadeBuf
    port map (
            O => \N__33176\,
            I => \N__33170\
        );

    \I__6184\ : CascadeBuf
    port map (
            O => \N__33173\,
            I => \N__33167\
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__33170\,
            I => \N__33164\
        );

    \I__6182\ : CascadeMux
    port map (
            O => \N__33167\,
            I => \N__33161\
        );

    \I__6181\ : InMux
    port map (
            O => \N__33164\,
            I => \N__33158\
        );

    \I__6180\ : CascadeBuf
    port map (
            O => \N__33161\,
            I => \N__33155\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__33158\,
            I => \N__33152\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__33155\,
            I => \N__33149\
        );

    \I__6177\ : Span4Mux_v
    port map (
            O => \N__33152\,
            I => \N__33146\
        );

    \I__6176\ : InMux
    port map (
            O => \N__33149\,
            I => \N__33143\
        );

    \I__6175\ : Sp12to4
    port map (
            O => \N__33146\,
            I => \N__33139\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__33143\,
            I => \N__33136\
        );

    \I__6173\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33133\
        );

    \I__6172\ : Span12Mux_h
    port map (
            O => \N__33139\,
            I => \N__33130\
        );

    \I__6171\ : Span4Mux_v
    port map (
            O => \N__33136\,
            I => \N__33127\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__33133\,
            I => \N__33120\
        );

    \I__6169\ : Span12Mux_v
    port map (
            O => \N__33130\,
            I => \N__33120\
        );

    \I__6168\ : Sp12to4
    port map (
            O => \N__33127\,
            I => \N__33120\
        );

    \I__6167\ : Odrv12
    port map (
            O => \N__33120\,
            I => data_count_5
        );

    \I__6166\ : InMux
    port map (
            O => \N__33117\,
            I => n19769
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__33114\,
            I => \N__33110\
        );

    \I__6164\ : InMux
    port map (
            O => \N__33113\,
            I => \N__33107\
        );

    \I__6163\ : InMux
    port map (
            O => \N__33110\,
            I => \N__33104\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__33107\,
            I => \N__33101\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__33104\,
            I => \N__33098\
        );

    \I__6160\ : Span4Mux_v
    port map (
            O => \N__33101\,
            I => \N__33092\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__33098\,
            I => \N__33092\
        );

    \I__6158\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33089\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__33092\,
            I => cmd_rdadctmp_21
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__33089\,
            I => cmd_rdadctmp_21
        );

    \I__6155\ : CascadeMux
    port map (
            O => \N__33084\,
            I => \N__33080\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__33083\,
            I => \N__33076\
        );

    \I__6153\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33073\
        );

    \I__6152\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33070\
        );

    \I__6151\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33067\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__33073\,
            I => \N__33064\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33061\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__33067\,
            I => \N__33056\
        );

    \I__6147\ : Span4Mux_v
    port map (
            O => \N__33064\,
            I => \N__33056\
        );

    \I__6146\ : Span12Mux_h
    port map (
            O => \N__33061\,
            I => \N__33053\
        );

    \I__6145\ : Odrv4
    port map (
            O => \N__33056\,
            I => buf_adcdata_iac_13
        );

    \I__6144\ : Odrv12
    port map (
            O => \N__33053\,
            I => buf_adcdata_iac_13
        );

    \I__6143\ : InMux
    port map (
            O => \N__33048\,
            I => \N__33045\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__33042\
        );

    \I__6141\ : Span12Mux_h
    port map (
            O => \N__33042\,
            I => \N__33037\
        );

    \I__6140\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33032\
        );

    \I__6139\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33032\
        );

    \I__6138\ : Odrv12
    port map (
            O => \N__33037\,
            I => \acadc_skipCount_13\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__33032\,
            I => \acadc_skipCount_13\
        );

    \I__6136\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33024\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__33020\
        );

    \I__6134\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33017\
        );

    \I__6133\ : Sp12to4
    port map (
            O => \N__33020\,
            I => \N__33013\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__33017\,
            I => \N__33010\
        );

    \I__6131\ : InMux
    port map (
            O => \N__33016\,
            I => \N__33007\
        );

    \I__6130\ : Span12Mux_v
    port map (
            O => \N__33013\,
            I => \N__33004\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__33010\,
            I => buf_dds0_5
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__33007\,
            I => buf_dds0_5
        );

    \I__6127\ : Odrv12
    port map (
            O => \N__33004\,
            I => buf_dds0_5
        );

    \I__6126\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32992\
        );

    \I__6125\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32989\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32995\,
            I => \N__32986\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__32992\,
            I => \N__32983\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__32989\,
            I => buf_dds0_3
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__32986\,
            I => buf_dds0_3
        );

    \I__6120\ : Odrv4
    port map (
            O => \N__32983\,
            I => buf_dds0_3
        );

    \I__6119\ : InMux
    port map (
            O => \N__32976\,
            I => \N__32972\
        );

    \I__6118\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32968\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__32972\,
            I => \N__32965\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32962\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__32968\,
            I => \acadc_skipCount_5\
        );

    \I__6114\ : Odrv12
    port map (
            O => \N__32965\,
            I => \acadc_skipCount_5\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32962\,
            I => \acadc_skipCount_5\
        );

    \I__6112\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32952\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__32952\,
            I => n20_adj_1670
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__32949\,
            I => \n8_adj_1560_cascade_\
        );

    \I__6109\ : CascadeMux
    port map (
            O => \N__32946\,
            I => \N__32943\
        );

    \I__6108\ : CascadeBuf
    port map (
            O => \N__32943\,
            I => \N__32940\
        );

    \I__6107\ : CascadeMux
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__6106\ : CascadeBuf
    port map (
            O => \N__32937\,
            I => \N__32934\
        );

    \I__6105\ : CascadeMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__6104\ : CascadeBuf
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__6103\ : CascadeMux
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__6102\ : CascadeBuf
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__6101\ : CascadeMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__6100\ : CascadeBuf
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__32916\,
            I => \N__32913\
        );

    \I__6098\ : CascadeBuf
    port map (
            O => \N__32913\,
            I => \N__32910\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__6096\ : CascadeBuf
    port map (
            O => \N__32907\,
            I => \N__32904\
        );

    \I__6095\ : CascadeMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__6094\ : CascadeBuf
    port map (
            O => \N__32901\,
            I => \N__32897\
        );

    \I__6093\ : CascadeMux
    port map (
            O => \N__32900\,
            I => \N__32894\
        );

    \I__6092\ : CascadeMux
    port map (
            O => \N__32897\,
            I => \N__32891\
        );

    \I__6091\ : CascadeBuf
    port map (
            O => \N__32894\,
            I => \N__32888\
        );

    \I__6090\ : CascadeBuf
    port map (
            O => \N__32891\,
            I => \N__32885\
        );

    \I__6089\ : CascadeMux
    port map (
            O => \N__32888\,
            I => \N__32882\
        );

    \I__6088\ : CascadeMux
    port map (
            O => \N__32885\,
            I => \N__32879\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32876\
        );

    \I__6086\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32873\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32870\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__32873\,
            I => \N__32867\
        );

    \I__6083\ : Span4Mux_h
    port map (
            O => \N__32870\,
            I => \N__32864\
        );

    \I__6082\ : Span4Mux_h
    port map (
            O => \N__32867\,
            I => \N__32861\
        );

    \I__6081\ : Span4Mux_v
    port map (
            O => \N__32864\,
            I => \N__32858\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__32861\,
            I => \N__32855\
        );

    \I__6079\ : Span4Mux_h
    port map (
            O => \N__32858\,
            I => \N__32852\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__32855\,
            I => \N__32849\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__32852\,
            I => \data_index_9_N_212_7\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__32849\,
            I => \data_index_9_N_212_7\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32841\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32841\,
            I => n24_adj_1593
        );

    \I__6073\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32835\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32832\
        );

    \I__6071\ : Odrv12
    port map (
            O => \N__32832\,
            I => n23_adj_1591
        );

    \I__6070\ : CascadeMux
    port map (
            O => \N__32829\,
            I => \n22_adj_1590_cascade_\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32826\,
            I => \N__32823\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__32823\,
            I => n18
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__32820\,
            I => \n30_adj_1543_cascade_\
        );

    \I__6066\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32810\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32810\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32807\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__32810\,
            I => \N__32804\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32801\
        );

    \I__6061\ : Odrv4
    port map (
            O => \N__32804\,
            I => n31_adj_1537
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__32801\,
            I => n31_adj_1537
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__32796\,
            I => \N__32793\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32790\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32787\
        );

    \I__6056\ : Span4Mux_v
    port map (
            O => \N__32787\,
            I => \N__32783\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__32786\,
            I => \N__32780\
        );

    \I__6054\ : Span4Mux_h
    port map (
            O => \N__32783\,
            I => \N__32776\
        );

    \I__6053\ : InMux
    port map (
            O => \N__32780\,
            I => \N__32773\
        );

    \I__6052\ : InMux
    port map (
            O => \N__32779\,
            I => \N__32770\
        );

    \I__6051\ : Odrv4
    port map (
            O => \N__32776\,
            I => cmd_rdadctmp_26
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32773\,
            I => cmd_rdadctmp_26
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__32770\,
            I => cmd_rdadctmp_26
        );

    \I__6048\ : InMux
    port map (
            O => \N__32763\,
            I => \N__32760\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__32760\,
            I => \N__32757\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__32757\,
            I => \N__32753\
        );

    \I__6045\ : InMux
    port map (
            O => \N__32756\,
            I => \N__32750\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__32753\,
            I => \N__32746\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__32750\,
            I => \N__32743\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32740\
        );

    \I__6041\ : Span4Mux_h
    port map (
            O => \N__32746\,
            I => \N__32737\
        );

    \I__6040\ : Span4Mux_v
    port map (
            O => \N__32743\,
            I => \N__32734\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__32740\,
            I => buf_adcdata_iac_18
        );

    \I__6038\ : Odrv4
    port map (
            O => \N__32737\,
            I => buf_adcdata_iac_18
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__32734\,
            I => buf_adcdata_iac_18
        );

    \I__6036\ : InMux
    port map (
            O => \N__32727\,
            I => \N__32723\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32726\,
            I => \N__32720\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__32723\,
            I => \N__32716\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__32720\,
            I => \N__32713\
        );

    \I__6032\ : InMux
    port map (
            O => \N__32719\,
            I => \N__32710\
        );

    \I__6031\ : Span4Mux_v
    port map (
            O => \N__32716\,
            I => \N__32707\
        );

    \I__6030\ : Span4Mux_h
    port map (
            O => \N__32713\,
            I => \N__32704\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__32710\,
            I => \acadc_skipCount_8\
        );

    \I__6028\ : Odrv4
    port map (
            O => \N__32707\,
            I => \acadc_skipCount_8\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__32704\,
            I => \acadc_skipCount_8\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__32697\,
            I => \n14_adj_1538_cascade_\
        );

    \I__6025\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32691\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32691\,
            I => n26_adj_1525
        );

    \I__6023\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32684\
        );

    \I__6022\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32680\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__32684\,
            I => \N__32677\
        );

    \I__6020\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32674\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__32680\,
            I => buf_dds1_3
        );

    \I__6018\ : Odrv12
    port map (
            O => \N__32677\,
            I => buf_dds1_3
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__32674\,
            I => buf_dds1_3
        );

    \I__6016\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32664\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__32664\,
            I => \N__32661\
        );

    \I__6014\ : Span4Mux_h
    port map (
            O => \N__32661\,
            I => \N__32656\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32660\,
            I => \N__32651\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32651\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__32656\,
            I => \acadc_skipCount_4\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__32651\,
            I => \acadc_skipCount_4\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32643\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__32643\,
            I => n8_adj_1560
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__32640\,
            I => \n30_adj_1631_cascade_\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32634\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__32634\,
            I => \N__32631\
        );

    \I__6004\ : Sp12to4
    port map (
            O => \N__32631\,
            I => \N__32628\
        );

    \I__6003\ : Odrv12
    port map (
            O => \N__32628\,
            I => n9
        );

    \I__6002\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__32622\,
            I => \N__32619\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__32619\,
            I => \N__32616\
        );

    \I__5999\ : Span4Mux_h
    port map (
            O => \N__32616\,
            I => \N__32613\
        );

    \I__5998\ : Span4Mux_h
    port map (
            O => \N__32613\,
            I => \N__32610\
        );

    \I__5997\ : Span4Mux_v
    port map (
            O => \N__32610\,
            I => \N__32607\
        );

    \I__5996\ : Odrv4
    port map (
            O => \N__32607\,
            I => buf_data_iac_22
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__32604\,
            I => \N__32601\
        );

    \I__5994\ : InMux
    port map (
            O => \N__32601\,
            I => \N__32597\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__32600\,
            I => \N__32594\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__32597\,
            I => \N__32591\
        );

    \I__5991\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32588\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__32591\,
            I => \N__32585\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__32588\,
            I => data_idxvec_14
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__32585\,
            I => data_idxvec_14
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__32580\,
            I => \N__32577\
        );

    \I__5986\ : InMux
    port map (
            O => \N__32577\,
            I => \N__32574\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__32574\,
            I => \N__32571\
        );

    \I__5984\ : Span4Mux_v
    port map (
            O => \N__32571\,
            I => \N__32568\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__32568\,
            I => \N__32565\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__32565\,
            I => n21330
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__32562\,
            I => \N__32558\
        );

    \I__5980\ : InMux
    port map (
            O => \N__32561\,
            I => \N__32555\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32551\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__32555\,
            I => \N__32548\
        );

    \I__5977\ : InMux
    port map (
            O => \N__32554\,
            I => \N__32545\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__32551\,
            I => \acadc_skipCount_11\
        );

    \I__5975\ : Odrv4
    port map (
            O => \N__32548\,
            I => \acadc_skipCount_11\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__32545\,
            I => \acadc_skipCount_11\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__32538\,
            I => \N__32535\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32532\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32529\
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__32529\,
            I => n23_adj_1677
        );

    \I__5969\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32522\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32525\,
            I => \N__32519\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__32522\,
            I => \N__32513\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__32519\,
            I => \N__32513\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32518\,
            I => \N__32510\
        );

    \I__5964\ : Span4Mux_v
    port map (
            O => \N__32513\,
            I => \N__32507\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__32510\,
            I => \N__32502\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__32507\,
            I => \N__32502\
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__32502\,
            I => buf_dds1_9
        );

    \I__5960\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32496\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__32496\,
            I => \N__32493\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__32493\,
            I => \N__32490\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__32490\,
            I => \N__32486\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__32489\,
            I => \N__32483\
        );

    \I__5955\ : Span4Mux_h
    port map (
            O => \N__32486\,
            I => \N__32480\
        );

    \I__5954\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32477\
        );

    \I__5953\ : Odrv4
    port map (
            O => \N__32480\,
            I => buf_adcdata_vdc_14
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__32477\,
            I => buf_adcdata_vdc_14
        );

    \I__5951\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32469\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__32469\,
            I => \N__32465\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32462\
        );

    \I__5948\ : Span12Mux_v
    port map (
            O => \N__32465\,
            I => \N__32458\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__32462\,
            I => \N__32455\
        );

    \I__5946\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32452\
        );

    \I__5945\ : Span12Mux_h
    port map (
            O => \N__32458\,
            I => \N__32449\
        );

    \I__5944\ : Span4Mux_h
    port map (
            O => \N__32455\,
            I => \N__32446\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32452\,
            I => buf_adcdata_vac_14
        );

    \I__5942\ : Odrv12
    port map (
            O => \N__32449\,
            I => buf_adcdata_vac_14
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__32446\,
            I => buf_adcdata_vac_14
        );

    \I__5940\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32436\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__32433\,
            I => n20
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__32430\,
            I => \n17_cascade_\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__32424\,
            I => n19_adj_1526
        );

    \I__5934\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32415\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32420\,
            I => \N__32415\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__32415\,
            I => n29
        );

    \I__5931\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32408\
        );

    \I__5930\ : CascadeMux
    port map (
            O => \N__32411\,
            I => \N__32405\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32408\,
            I => \N__32402\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32405\,
            I => \N__32399\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__32402\,
            I => \N__32396\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32399\,
            I => data_idxvec_13
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__32396\,
            I => data_idxvec_13
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__32391\,
            I => \N__32387\
        );

    \I__5923\ : InMux
    port map (
            O => \N__32390\,
            I => \N__32384\
        );

    \I__5922\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32381\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32384\,
            I => \N__32378\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32372\
        );

    \I__5919\ : Span4Mux_h
    port map (
            O => \N__32378\,
            I => \N__32372\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32369\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__32372\,
            I => comm_cmd_4
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__32369\,
            I => comm_cmd_4
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__32364\,
            I => \n16818_cascade_\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32358\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__32358\,
            I => \N__32355\
        );

    \I__5912\ : Span4Mux_v
    port map (
            O => \N__32355\,
            I => \N__32352\
        );

    \I__5911\ : Span4Mux_h
    port map (
            O => \N__32352\,
            I => \N__32349\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__32349\,
            I => n16_adj_1628
        );

    \I__5909\ : InMux
    port map (
            O => \N__32346\,
            I => \N__32343\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__32343\,
            I => \N__32340\
        );

    \I__5907\ : Span4Mux_h
    port map (
            O => \N__32340\,
            I => \N__32337\
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__32337\,
            I => n22365
        );

    \I__5905\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32331\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__32331\,
            I => \N__32328\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__32328\,
            I => \N__32324\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32327\,
            I => \N__32321\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__32324\,
            I => \N__32318\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__32321\,
            I => data_idxvec_5
        );

    \I__5899\ : Odrv4
    port map (
            O => \N__32318\,
            I => data_idxvec_5
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__32313\,
            I => \n26_adj_1630_cascade_\
        );

    \I__5897\ : CascadeMux
    port map (
            O => \N__32310\,
            I => \n22449_cascade_\
        );

    \I__5896\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32302\
        );

    \I__5895\ : CascadeMux
    port map (
            O => \N__32306\,
            I => \N__32299\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32305\,
            I => \N__32296\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__32302\,
            I => \N__32293\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32299\,
            I => \N__32290\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__32296\,
            I => req_data_cnt_5
        );

    \I__5890\ : Odrv4
    port map (
            O => \N__32293\,
            I => req_data_cnt_5
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__32290\,
            I => req_data_cnt_5
        );

    \I__5888\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32280\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__32280\,
            I => n22368
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__32277\,
            I => \n22452_cascade_\
        );

    \I__5885\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__32271\,
            I => \N__32267\
        );

    \I__5883\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32264\
        );

    \I__5882\ : Span4Mux_h
    port map (
            O => \N__32267\,
            I => \N__32261\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__32264\,
            I => n14_adj_1551
        );

    \I__5880\ : Odrv4
    port map (
            O => \N__32261\,
            I => n14_adj_1551
        );

    \I__5879\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32252\
        );

    \I__5878\ : InMux
    port map (
            O => \N__32255\,
            I => \N__32249\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__32252\,
            I => \N__32246\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__32249\,
            I => \N__32242\
        );

    \I__5875\ : Span12Mux_v
    port map (
            O => \N__32246\,
            I => \N__32239\
        );

    \I__5874\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32236\
        );

    \I__5873\ : Span4Mux_v
    port map (
            O => \N__32242\,
            I => \N__32233\
        );

    \I__5872\ : Odrv12
    port map (
            O => \N__32239\,
            I => buf_dds0_4
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__32236\,
            I => buf_dds0_4
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__32233\,
            I => buf_dds0_4
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__5868\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32220\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__32220\,
            I => n23_adj_1661
        );

    \I__5866\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32212\
        );

    \I__5865\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32207\
        );

    \I__5864\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32207\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__32212\,
            I => \acadc_skipCount_14\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__32207\,
            I => \acadc_skipCount_14\
        );

    \I__5861\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32199\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__32199\,
            I => \N__32196\
        );

    \I__5859\ : Span4Mux_v
    port map (
            O => \N__32196\,
            I => \N__32192\
        );

    \I__5858\ : InMux
    port map (
            O => \N__32195\,
            I => \N__32189\
        );

    \I__5857\ : Odrv4
    port map (
            O => \N__32192\,
            I => buf_adcdata_vdc_1
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__32189\,
            I => buf_adcdata_vdc_1
        );

    \I__5855\ : InMux
    port map (
            O => \N__32184\,
            I => \N__32181\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__5853\ : Span4Mux_h
    port map (
            O => \N__32178\,
            I => \N__32175\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__32175\,
            I => \N__32171\
        );

    \I__5851\ : InMux
    port map (
            O => \N__32174\,
            I => \N__32168\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__32171\,
            I => \N__32163\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__32168\,
            I => \N__32163\
        );

    \I__5848\ : Span4Mux_h
    port map (
            O => \N__32163\,
            I => \N__32159\
        );

    \I__5847\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32156\
        );

    \I__5846\ : Span4Mux_h
    port map (
            O => \N__32159\,
            I => \N__32153\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__32156\,
            I => buf_adcdata_vac_1
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__32153\,
            I => buf_adcdata_vac_1
        );

    \I__5843\ : InMux
    port map (
            O => \N__32148\,
            I => \N__32145\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__32145\,
            I => \N__32142\
        );

    \I__5841\ : Span4Mux_v
    port map (
            O => \N__32142\,
            I => \N__32138\
        );

    \I__5840\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32135\
        );

    \I__5839\ : Sp12to4
    port map (
            O => \N__32138\,
            I => \N__32132\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__32135\,
            I => \N__32129\
        );

    \I__5837\ : Span12Mux_h
    port map (
            O => \N__32132\,
            I => \N__32125\
        );

    \I__5836\ : Span4Mux_v
    port map (
            O => \N__32129\,
            I => \N__32122\
        );

    \I__5835\ : InMux
    port map (
            O => \N__32128\,
            I => \N__32119\
        );

    \I__5834\ : Span12Mux_v
    port map (
            O => \N__32125\,
            I => \N__32116\
        );

    \I__5833\ : Span4Mux_v
    port map (
            O => \N__32122\,
            I => \N__32113\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__32119\,
            I => buf_adcdata_iac_20
        );

    \I__5831\ : Odrv12
    port map (
            O => \N__32116\,
            I => buf_adcdata_iac_20
        );

    \I__5830\ : Odrv4
    port map (
            O => \N__32113\,
            I => buf_adcdata_iac_20
        );

    \I__5829\ : IoInMux
    port map (
            O => \N__32106\,
            I => \N__32103\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32100\
        );

    \I__5827\ : Span4Mux_s1_h
    port map (
            O => \N__32100\,
            I => \N__32097\
        );

    \I__5826\ : Sp12to4
    port map (
            O => \N__32097\,
            I => \N__32094\
        );

    \I__5825\ : Span12Mux_v
    port map (
            O => \N__32094\,
            I => \N__32091\
        );

    \I__5824\ : Span12Mux_h
    port map (
            O => \N__32091\,
            I => \N__32086\
        );

    \I__5823\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32083\
        );

    \I__5822\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32080\
        );

    \I__5821\ : Odrv12
    port map (
            O => \N__32086\,
            I => \VAC_OSR0\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__32083\,
            I => \VAC_OSR0\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__32080\,
            I => \VAC_OSR0\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__32073\,
            I => \N__32070\
        );

    \I__5817\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32066\
        );

    \I__5816\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32063\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__32060\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__32063\,
            I => \N__32057\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__32060\,
            I => \N__32054\
        );

    \I__5812\ : Span4Mux_v
    port map (
            O => \N__32057\,
            I => \N__32049\
        );

    \I__5811\ : Span4Mux_h
    port map (
            O => \N__32054\,
            I => \N__32049\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__32049\,
            I => n30
        );

    \I__5809\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32043\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32039\
        );

    \I__5807\ : InMux
    port map (
            O => \N__32042\,
            I => \N__32036\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__32039\,
            I => \N__32033\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__32030\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__32033\,
            I => \N__32025\
        );

    \I__5803\ : Span4Mux_v
    port map (
            O => \N__32030\,
            I => \N__32025\
        );

    \I__5802\ : Span4Mux_v
    port map (
            O => \N__32025\,
            I => \N__32022\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__32022\,
            I => n14_adj_1574
        );

    \I__5800\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__5798\ : Span4Mux_h
    port map (
            O => \N__32013\,
            I => \N__32010\
        );

    \I__5797\ : Span4Mux_h
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__5796\ : Span4Mux_v
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__5795\ : Odrv4
    port map (
            O => \N__32004\,
            I => buf_data_iac_3
        );

    \I__5794\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31998\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31995\
        );

    \I__5792\ : Odrv12
    port map (
            O => \N__31995\,
            I => n22_adj_1610
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__31992\,
            I => \N__31987\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31991\,
            I => \N__31982\
        );

    \I__5789\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31982\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31979\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__31982\,
            I => req_data_cnt_14
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__31979\,
            I => req_data_cnt_14
        );

    \I__5785\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31971\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__31971\,
            I => \N__31968\
        );

    \I__5783\ : Span12Mux_v
    port map (
            O => \N__31968\,
            I => \N__31963\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31958\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31958\
        );

    \I__5780\ : Odrv12
    port map (
            O => \N__31963\,
            I => req_data_cnt_11
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31958\,
            I => req_data_cnt_11
        );

    \I__5778\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31950\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__31950\,
            I => n23
        );

    \I__5776\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31944\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31944\,
            I => \ADC_VDC.n21211\
        );

    \I__5774\ : CEMux
    port map (
            O => \N__31941\,
            I => \N__31938\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31938\,
            I => \N__31935\
        );

    \I__5772\ : Odrv4
    port map (
            O => \N__31935\,
            I => \ADC_VDC.n13368\
        );

    \I__5771\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31925\
        );

    \I__5769\ : InMux
    port map (
            O => \N__31928\,
            I => \N__31922\
        );

    \I__5768\ : Span4Mux_h
    port map (
            O => \N__31925\,
            I => \N__31919\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__31922\,
            I => secclk_cnt_20
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__31919\,
            I => secclk_cnt_20
        );

    \I__5765\ : CascadeMux
    port map (
            O => \N__31914\,
            I => \n20048_cascade_\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31908\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31905\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__31905\,
            I => n14
        );

    \I__5761\ : InMux
    port map (
            O => \N__31902\,
            I => \N__31899\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__5759\ : Span4Mux_h
    port map (
            O => \N__31896\,
            I => \N__31892\
        );

    \I__5758\ : InMux
    port map (
            O => \N__31895\,
            I => \N__31889\
        );

    \I__5757\ : Odrv4
    port map (
            O => \N__31892\,
            I => buf_adcdata_vdc_20
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__31889\,
            I => buf_adcdata_vdc_20
        );

    \I__5755\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31881\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__31881\,
            I => \N__31878\
        );

    \I__5753\ : Span4Mux_h
    port map (
            O => \N__31878\,
            I => \N__31875\
        );

    \I__5752\ : Span4Mux_v
    port map (
            O => \N__31875\,
            I => \N__31872\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__31872\,
            I => \N__31868\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31871\,
            I => \N__31865\
        );

    \I__5749\ : Span4Mux_h
    port map (
            O => \N__31868\,
            I => \N__31860\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31860\
        );

    \I__5747\ : Span4Mux_h
    port map (
            O => \N__31860\,
            I => \N__31856\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31853\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__31856\,
            I => \N__31850\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__31853\,
            I => buf_adcdata_vac_20
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__31850\,
            I => buf_adcdata_vac_20
        );

    \I__5742\ : InMux
    port map (
            O => \N__31845\,
            I => \N__31841\
        );

    \I__5741\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31838\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__31841\,
            I => secclk_cnt_6
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__31838\,
            I => secclk_cnt_6
        );

    \I__5738\ : InMux
    port map (
            O => \N__31833\,
            I => \N__31829\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31832\,
            I => \N__31826\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__31829\,
            I => secclk_cnt_14
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31826\,
            I => secclk_cnt_14
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__31821\,
            I => \N__31818\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31818\,
            I => \N__31814\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31811\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__31814\,
            I => \N__31808\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31811\,
            I => secclk_cnt_10
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__31808\,
            I => secclk_cnt_10
        );

    \I__5728\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31799\
        );

    \I__5727\ : InMux
    port map (
            O => \N__31802\,
            I => \N__31796\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__31799\,
            I => secclk_cnt_3
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31796\,
            I => secclk_cnt_3
        );

    \I__5724\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__31788\,
            I => n27
        );

    \I__5722\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31781\
        );

    \I__5721\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31778\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__31781\,
            I => secclk_cnt_2
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__31778\,
            I => secclk_cnt_2
        );

    \I__5718\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31769\
        );

    \I__5717\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31766\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__31769\,
            I => secclk_cnt_13
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__31766\,
            I => secclk_cnt_13
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__31761\,
            I => \N__31757\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31754\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31757\,
            I => \N__31751\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__31754\,
            I => secclk_cnt_7
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__31751\,
            I => secclk_cnt_7
        );

    \I__5709\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31742\
        );

    \I__5708\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31739\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__31742\,
            I => secclk_cnt_16
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__31739\,
            I => secclk_cnt_16
        );

    \I__5705\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__31731\,
            I => n26_adj_1656
        );

    \I__5703\ : InMux
    port map (
            O => \N__31728\,
            I => \N__31724\
        );

    \I__5702\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31721\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__31724\,
            I => \N__31718\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__31721\,
            I => \N__31715\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__31718\,
            I => \N__31710\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__31715\,
            I => \N__31710\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__31710\,
            I => n14_adj_1552
        );

    \I__5696\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31704\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__31704\,
            I => \ADC_VDC.n11\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31698\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__31698\,
            I => \ADC_VDC.n65\
        );

    \I__5692\ : CascadeMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31692\,
            I => \N__31689\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__31689\,
            I => \ADC_VDC.n21133\
        );

    \I__5689\ : CEMux
    port map (
            O => \N__31686\,
            I => \N__31683\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__31683\,
            I => \ADC_VDC.n42_adj_1452\
        );

    \I__5687\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__31674\,
            I => \ADC_VDC.n20998\
        );

    \I__5684\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31668\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__31668\,
            I => \ADC_VDC.n11494\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__31665\,
            I => \ADC_VDC.n11494_cascade_\
        );

    \I__5681\ : CascadeMux
    port map (
            O => \N__31662\,
            I => \N__31658\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31655\
        );

    \I__5679\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31652\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31649\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__31652\,
            I => \N__31646\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__31649\,
            I => \N__31643\
        );

    \I__5675\ : Span4Mux_v
    port map (
            O => \N__31646\,
            I => \N__31640\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__31643\,
            I => \ADC_VDC.n15\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__31640\,
            I => \ADC_VDC.n15\
        );

    \I__5672\ : CascadeMux
    port map (
            O => \N__31635\,
            I => \ADC_VDC.n15_cascade_\
        );

    \I__5671\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31629\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__31629\,
            I => \ADC_VDC.n21185\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31621\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31614\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__31624\,
            I => \N__31611\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31621\,
            I => \N__31605\
        );

    \I__5665\ : InMux
    port map (
            O => \N__31620\,
            I => \N__31602\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__31619\,
            I => \N__31597\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__31618\,
            I => \N__31594\
        );

    \I__5662\ : CascadeMux
    port map (
            O => \N__31617\,
            I => \N__31591\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__31614\,
            I => \N__31577\
        );

    \I__5660\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31570\
        );

    \I__5659\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31570\
        );

    \I__5658\ : InMux
    port map (
            O => \N__31609\,
            I => \N__31570\
        );

    \I__5657\ : InMux
    port map (
            O => \N__31608\,
            I => \N__31567\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__31605\,
            I => \N__31562\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__31602\,
            I => \N__31562\
        );

    \I__5654\ : InMux
    port map (
            O => \N__31601\,
            I => \N__31549\
        );

    \I__5653\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31549\
        );

    \I__5652\ : InMux
    port map (
            O => \N__31597\,
            I => \N__31549\
        );

    \I__5651\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31549\
        );

    \I__5650\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31549\
        );

    \I__5649\ : InMux
    port map (
            O => \N__31590\,
            I => \N__31549\
        );

    \I__5648\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31540\
        );

    \I__5647\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31540\
        );

    \I__5646\ : InMux
    port map (
            O => \N__31587\,
            I => \N__31540\
        );

    \I__5645\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31540\
        );

    \I__5644\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31537\
        );

    \I__5643\ : InMux
    port map (
            O => \N__31584\,
            I => \N__31526\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31583\,
            I => \N__31526\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31526\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31581\,
            I => \N__31526\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31580\,
            I => \N__31526\
        );

    \I__5638\ : Span4Mux_v
    port map (
            O => \N__31577\,
            I => \N__31521\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__31570\,
            I => \N__31521\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__31567\,
            I => \N__31518\
        );

    \I__5635\ : Span4Mux_h
    port map (
            O => \N__31562\,
            I => \N__31513\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__31549\,
            I => \N__31513\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__31540\,
            I => \N__31502\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__31537\,
            I => \N__31502\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__31526\,
            I => \N__31502\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__31521\,
            I => \N__31502\
        );

    \I__5629\ : Span4Mux_v
    port map (
            O => \N__31518\,
            I => \N__31502\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__31513\,
            I => n11891
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__31502\,
            I => n11891
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__31497\,
            I => \N__31494\
        );

    \I__5625\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31490\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__31493\,
            I => \N__31487\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__31490\,
            I => \N__31484\
        );

    \I__5622\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31481\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__31484\,
            I => \N__31478\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__31481\,
            I => \N__31475\
        );

    \I__5619\ : Odrv4
    port map (
            O => \N__31478\,
            I => cmd_rdadcbuf_12
        );

    \I__5618\ : Odrv4
    port map (
            O => \N__31475\,
            I => cmd_rdadcbuf_12
        );

    \I__5617\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31467\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__31467\,
            I => \ADC_VDC.n21203\
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__31464\,
            I => \N__31461\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31458\
        );

    \I__5613\ : LocalMux
    port map (
            O => \N__31458\,
            I => \SIG_DDS.tmp_buf_1\
        );

    \I__5612\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31452\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N__31449\
        );

    \I__5610\ : Span4Mux_v
    port map (
            O => \N__31449\,
            I => \N__31444\
        );

    \I__5609\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31439\
        );

    \I__5608\ : InMux
    port map (
            O => \N__31447\,
            I => \N__31439\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__31444\,
            I => buf_dds0_2
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__31439\,
            I => buf_dds0_2
        );

    \I__5605\ : CascadeMux
    port map (
            O => \N__31434\,
            I => \N__31431\
        );

    \I__5604\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31428\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31428\,
            I => \SIG_DDS.tmp_buf_2\
        );

    \I__5602\ : CascadeMux
    port map (
            O => \N__31425\,
            I => \N__31422\
        );

    \I__5601\ : InMux
    port map (
            O => \N__31422\,
            I => \N__31419\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__31419\,
            I => \SIG_DDS.tmp_buf_3\
        );

    \I__5599\ : CascadeMux
    port map (
            O => \N__31416\,
            I => \N__31413\
        );

    \I__5598\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__31410\,
            I => \SIG_DDS.tmp_buf_4\
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__31401\,
            I => \SIG_DDS.tmp_buf_5\
        );

    \I__5593\ : CascadeMux
    port map (
            O => \N__31398\,
            I => \N__31395\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31395\,
            I => \N__31392\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__31392\,
            I => \N__31389\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__31389\,
            I => \ADC_VDC.n21007\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__31386\,
            I => \ADC_VDC.n21007_cascade_\
        );

    \I__5588\ : SRMux
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__31380\,
            I => \ADC_VDC.n4\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__31377\,
            I => \N__31374\
        );

    \I__5585\ : InMux
    port map (
            O => \N__31374\,
            I => \N__31371\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31371\,
            I => \SIG_DDS.tmp_buf_10\
        );

    \I__5583\ : InMux
    port map (
            O => \N__31368\,
            I => \N__31363\
        );

    \I__5582\ : InMux
    port map (
            O => \N__31367\,
            I => \N__31360\
        );

    \I__5581\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31357\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__31363\,
            I => buf_dds0_11
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__31360\,
            I => buf_dds0_11
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__31357\,
            I => buf_dds0_11
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__31350\,
            I => \N__31347\
        );

    \I__5576\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31344\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__31344\,
            I => \SIG_DDS.tmp_buf_11\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__31341\,
            I => \N__31338\
        );

    \I__5573\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31335\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__31335\,
            I => \SIG_DDS.tmp_buf_12\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__31332\,
            I => \N__31329\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31329\,
            I => \N__31326\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__31326\,
            I => \SIG_DDS.tmp_buf_13\
        );

    \I__5568\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31315\
        );

    \I__5566\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31312\
        );

    \I__5565\ : InMux
    port map (
            O => \N__31318\,
            I => \N__31309\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__31315\,
            I => \N__31306\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__31312\,
            I => buf_dds0_14
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__31309\,
            I => buf_dds0_14
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__31306\,
            I => buf_dds0_14
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__31299\,
            I => \N__31295\
        );

    \I__5559\ : CascadeMux
    port map (
            O => \N__31298\,
            I => \N__31291\
        );

    \I__5558\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31288\
        );

    \I__5557\ : CascadeMux
    port map (
            O => \N__31294\,
            I => \N__31285\
        );

    \I__5556\ : InMux
    port map (
            O => \N__31291\,
            I => \N__31282\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__31288\,
            I => \N__31279\
        );

    \I__5554\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31276\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__31282\,
            I => \N__31273\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__31279\,
            I => \N__31270\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__31276\,
            I => buf_dds0_15
        );

    \I__5550\ : Odrv12
    port map (
            O => \N__31273\,
            I => buf_dds0_15
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__31270\,
            I => buf_dds0_15
        );

    \I__5548\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31260\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__31260\,
            I => \SIG_DDS.tmp_buf_14\
        );

    \I__5546\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31254\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__31254\,
            I => \N__31249\
        );

    \I__5544\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31246\
        );

    \I__5543\ : InMux
    port map (
            O => \N__31252\,
            I => \N__31243\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__31249\,
            I => \N__31238\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31238\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__31243\,
            I => buf_dds0_9
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__31238\,
            I => buf_dds0_9
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__31233\,
            I => \N__31230\
        );

    \I__5537\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__31227\,
            I => \SIG_DDS.tmp_buf_9\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__31224\,
            I => \N__31221\
        );

    \I__5534\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__31218\,
            I => \N__31215\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__31215\,
            I => \SIG_DDS.tmp_buf_8\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__5530\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31206\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__31206\,
            I => \SIG_DDS.tmp_buf_0\
        );

    \I__5528\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31200\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__31200\,
            I => \N__31195\
        );

    \I__5526\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31190\
        );

    \I__5525\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31190\
        );

    \I__5524\ : Odrv4
    port map (
            O => \N__31195\,
            I => buf_dds0_1
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__31190\,
            I => buf_dds0_1
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__31185\,
            I => \N__31181\
        );

    \I__5521\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31178\
        );

    \I__5520\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31175\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N__31172\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__31175\,
            I => \N__31166\
        );

    \I__5517\ : Sp12to4
    port map (
            O => \N__31172\,
            I => \N__31166\
        );

    \I__5516\ : InMux
    port map (
            O => \N__31171\,
            I => \N__31163\
        );

    \I__5515\ : Odrv12
    port map (
            O => \N__31166\,
            I => \acadc_skipCount_15\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__31163\,
            I => \acadc_skipCount_15\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__31158\,
            I => \N__31155\
        );

    \I__5512\ : InMux
    port map (
            O => \N__31155\,
            I => \N__31151\
        );

    \I__5511\ : InMux
    port map (
            O => \N__31154\,
            I => \N__31148\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__31151\,
            I => \N__31145\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__31148\,
            I => n11570
        );

    \I__5508\ : Odrv12
    port map (
            O => \N__31145\,
            I => n11570
        );

    \I__5507\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31137\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__5505\ : Sp12to4
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__5504\ : Span12Mux_v
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__5503\ : Odrv12
    port map (
            O => \N__31128\,
            I => \EIS_SYNCCLK\
        );

    \I__5502\ : IoInMux
    port map (
            O => \N__31125\,
            I => \N__31122\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__31122\,
            I => \N__31118\
        );

    \I__5500\ : IoInMux
    port map (
            O => \N__31121\,
            I => \N__31115\
        );

    \I__5499\ : Span4Mux_s2_v
    port map (
            O => \N__31118\,
            I => \N__31112\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__31115\,
            I => \N__31109\
        );

    \I__5497\ : Span4Mux_v
    port map (
            O => \N__31112\,
            I => \N__31106\
        );

    \I__5496\ : IoSpan4Mux
    port map (
            O => \N__31109\,
            I => \N__31103\
        );

    \I__5495\ : Span4Mux_v
    port map (
            O => \N__31106\,
            I => \N__31098\
        );

    \I__5494\ : Span4Mux_s3_h
    port map (
            O => \N__31103\,
            I => \N__31098\
        );

    \I__5493\ : Sp12to4
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__5492\ : Odrv12
    port map (
            O => \N__31095\,
            I => \IAC_CLK\
        );

    \I__5491\ : InMux
    port map (
            O => \N__31092\,
            I => \N__31088\
        );

    \I__5490\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31085\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__31088\,
            I => \N__31082\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__31085\,
            I => \N__31078\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__31082\,
            I => \N__31075\
        );

    \I__5486\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31072\
        );

    \I__5485\ : Span4Mux_h
    port map (
            O => \N__31078\,
            I => \N__31069\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__31075\,
            I => buf_dds0_10
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__31072\,
            I => buf_dds0_10
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__31069\,
            I => buf_dds0_10
        );

    \I__5481\ : CascadeMux
    port map (
            O => \N__31062\,
            I => \n21501_cascade_\
        );

    \I__5480\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31056\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__31056\,
            I => \eis_state_2_N_392_0\
        );

    \I__5478\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31050\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__31050\,
            I => n22479
        );

    \I__5476\ : InMux
    port map (
            O => \N__31047\,
            I => \N__31040\
        );

    \I__5475\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31040\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__31045\,
            I => \N__31037\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__31040\,
            I => \N__31034\
        );

    \I__5472\ : InMux
    port map (
            O => \N__31037\,
            I => \N__31031\
        );

    \I__5471\ : Span4Mux_v
    port map (
            O => \N__31034\,
            I => \N__31025\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__31031\,
            I => \N__31022\
        );

    \I__5469\ : InMux
    port map (
            O => \N__31030\,
            I => \N__31017\
        );

    \I__5468\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31017\
        );

    \I__5467\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31014\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__31025\,
            I => \N__31011\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__31022\,
            I => \N__31006\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__31017\,
            I => \N__31006\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__31014\,
            I => eis_start
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__31011\,
            I => eis_start
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__31006\,
            I => eis_start
        );

    \I__5460\ : CascadeMux
    port map (
            O => \N__30999\,
            I => \n11_adj_1632_cascade_\
        );

    \I__5459\ : CEMux
    port map (
            O => \N__30996\,
            I => \N__30992\
        );

    \I__5458\ : CEMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30992\,
            I => n11908
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30989\,
            I => n11908
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__30984\,
            I => \N__30976\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__30983\,
            I => \N__30973\
        );

    \I__5453\ : CascadeMux
    port map (
            O => \N__30982\,
            I => \N__30970\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__30981\,
            I => \N__30959\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__30980\,
            I => \N__30956\
        );

    \I__5450\ : InMux
    port map (
            O => \N__30979\,
            I => \N__30944\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30976\,
            I => \N__30944\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30944\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30944\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30944\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30968\,
            I => \N__30937\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30967\,
            I => \N__30937\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30937\
        );

    \I__5442\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30932\
        );

    \I__5441\ : InMux
    port map (
            O => \N__30964\,
            I => \N__30932\
        );

    \I__5440\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30929\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30920\
        );

    \I__5438\ : InMux
    port map (
            O => \N__30959\,
            I => \N__30920\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30956\,
            I => \N__30920\
        );

    \I__5436\ : InMux
    port map (
            O => \N__30955\,
            I => \N__30920\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__30944\,
            I => eis_state_0
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__30937\,
            I => eis_state_0
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30932\,
            I => eis_state_0
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__30929\,
            I => eis_state_0
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30920\,
            I => eis_state_0
        );

    \I__5430\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30905\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30908\,
            I => \N__30902\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30905\,
            I => n21041
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__30902\,
            I => n21041
        );

    \I__5426\ : InMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__30894\,
            I => \N__30890\
        );

    \I__5424\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30886\
        );

    \I__5423\ : Span4Mux_h
    port map (
            O => \N__30890\,
            I => \N__30883\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30880\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30886\,
            I => buf_dds1_15
        );

    \I__5420\ : Odrv4
    port map (
            O => \N__30883\,
            I => buf_dds1_15
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30880\,
            I => buf_dds1_15
        );

    \I__5418\ : InMux
    port map (
            O => \N__30873\,
            I => \N__30869\
        );

    \I__5417\ : InMux
    port map (
            O => \N__30872\,
            I => \N__30866\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__30869\,
            I => \N__30863\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30857\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__30863\,
            I => \N__30857\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30862\,
            I => \N__30854\
        );

    \I__5412\ : Odrv4
    port map (
            O => \N__30857\,
            I => buf_dds1_10
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__30854\,
            I => buf_dds1_10
        );

    \I__5410\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \n22395_cascade_\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__30846\,
            I => \N__30842\
        );

    \I__5408\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30838\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30835\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30841\,
            I => \N__30832\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30827\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30827\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__30832\,
            I => req_data_cnt_8
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__30827\,
            I => req_data_cnt_8
        );

    \I__5401\ : IoInMux
    port map (
            O => \N__30822\,
            I => \N__30819\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__5399\ : Span4Mux_s3_h
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__5398\ : Span4Mux_h
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__5397\ : Span4Mux_h
    port map (
            O => \N__30810\,
            I => \N__30807\
        );

    \I__5396\ : Sp12to4
    port map (
            O => \N__30807\,
            I => \N__30802\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30799\
        );

    \I__5394\ : InMux
    port map (
            O => \N__30805\,
            I => \N__30796\
        );

    \I__5393\ : Span12Mux_v
    port map (
            O => \N__30802\,
            I => \N__30793\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__30799\,
            I => \N__30790\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__30796\,
            I => \N__30787\
        );

    \I__5390\ : Odrv12
    port map (
            O => \N__30793\,
            I => \VAC_FLT0\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__30790\,
            I => \VAC_FLT0\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__30787\,
            I => \VAC_FLT0\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__30780\,
            I => \N__30775\
        );

    \I__5386\ : InMux
    port map (
            O => \N__30779\,
            I => \N__30772\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__30778\,
            I => \N__30769\
        );

    \I__5384\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30766\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__30772\,
            I => \N__30763\
        );

    \I__5382\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30760\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__30766\,
            I => \N__30757\
        );

    \I__5380\ : Span4Mux_h
    port map (
            O => \N__30763\,
            I => \N__30754\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__30760\,
            I => \N__30749\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__30757\,
            I => \N__30749\
        );

    \I__5377\ : Sp12to4
    port map (
            O => \N__30754\,
            I => \N__30746\
        );

    \I__5376\ : Sp12to4
    port map (
            O => \N__30749\,
            I => \N__30741\
        );

    \I__5375\ : Span12Mux_v
    port map (
            O => \N__30746\,
            I => \N__30741\
        );

    \I__5374\ : Odrv12
    port map (
            O => \N__30741\,
            I => buf_adcdata_iac_22
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__30738\,
            I => \n22635_cascade_\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__5369\ : Odrv4
    port map (
            O => \N__30726\,
            I => n21236
        );

    \I__5368\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30718\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__30722\,
            I => \N__30715\
        );

    \I__5366\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30712\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__30718\,
            I => \N__30709\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30715\,
            I => \N__30706\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__30712\,
            I => \N__30703\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__30709\,
            I => \N__30700\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__30706\,
            I => \N__30697\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__30703\,
            I => \N__30694\
        );

    \I__5359\ : Sp12to4
    port map (
            O => \N__30700\,
            I => \N__30689\
        );

    \I__5358\ : Span12Mux_v
    port map (
            O => \N__30697\,
            I => \N__30689\
        );

    \I__5357\ : Span4Mux_h
    port map (
            O => \N__30694\,
            I => \N__30686\
        );

    \I__5356\ : Odrv12
    port map (
            O => \N__30689\,
            I => n14_adj_1578
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__30686\,
            I => n14_adj_1578
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__30681\,
            I => \n2_cascade_\
        );

    \I__5353\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30674\
        );

    \I__5352\ : CascadeMux
    port map (
            O => \N__30677\,
            I => \N__30671\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__30674\,
            I => \N__30668\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30671\,
            I => \N__30665\
        );

    \I__5349\ : Span4Mux_v
    port map (
            O => \N__30668\,
            I => \N__30662\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30657\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__30662\,
            I => \N__30657\
        );

    \I__5346\ : Sp12to4
    port map (
            O => \N__30657\,
            I => \N__30654\
        );

    \I__5345\ : Odrv12
    port map (
            O => \N__30654\,
            I => data_idxvec_4
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__30651\,
            I => \n26_adj_1635_cascade_\
        );

    \I__5343\ : CascadeMux
    port map (
            O => \N__30648\,
            I => \n22443_cascade_\
        );

    \I__5342\ : CascadeMux
    port map (
            O => \N__30645\,
            I => \n22446_cascade_\
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__30642\,
            I => \n30_adj_1636_cascade_\
        );

    \I__5340\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__30636\,
            I => n19_adj_1634
        );

    \I__5338\ : CascadeMux
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__5337\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__30624\,
            I => \N__30621\
        );

    \I__5334\ : Span4Mux_h
    port map (
            O => \N__30621\,
            I => \N__30617\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30614\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__30617\,
            I => \buf_readRTD_4\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__30614\,
            I => \buf_readRTD_4\
        );

    \I__5330\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30605\
        );

    \I__5329\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30602\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__30605\,
            I => \N__30598\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30602\,
            I => \N__30595\
        );

    \I__5326\ : InMux
    port map (
            O => \N__30601\,
            I => \N__30592\
        );

    \I__5325\ : Span12Mux_h
    port map (
            O => \N__30598\,
            I => \N__30589\
        );

    \I__5324\ : Span4Mux_v
    port map (
            O => \N__30595\,
            I => \N__30586\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__30592\,
            I => buf_adcdata_iac_12
        );

    \I__5322\ : Odrv12
    port map (
            O => \N__30589\,
            I => buf_adcdata_iac_12
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__30586\,
            I => buf_adcdata_iac_12
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__30579\,
            I => \n22467_cascade_\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30573\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__30570\,
            I => \N__30567\
        );

    \I__5316\ : Odrv4
    port map (
            O => \N__30567\,
            I => n16_adj_1633
        );

    \I__5315\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30561\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__30561\,
            I => n22470
        );

    \I__5313\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30555\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__30555\,
            I => \N__30552\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__30549\,
            I => n21329
        );

    \I__5309\ : IoInMux
    port map (
            O => \N__30546\,
            I => \N__30543\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__30543\,
            I => \N__30539\
        );

    \I__5307\ : InMux
    port map (
            O => \N__30542\,
            I => \N__30536\
        );

    \I__5306\ : IoSpan4Mux
    port map (
            O => \N__30539\,
            I => \N__30533\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__30536\,
            I => \N__30530\
        );

    \I__5304\ : Span4Mux_s2_v
    port map (
            O => \N__30533\,
            I => \N__30527\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__30530\,
            I => \N__30523\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__30527\,
            I => \N__30520\
        );

    \I__5301\ : InMux
    port map (
            O => \N__30526\,
            I => \N__30517\
        );

    \I__5300\ : Span4Mux_v
    port map (
            O => \N__30523\,
            I => \N__30514\
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__30520\,
            I => \IAC_FLT0\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__30517\,
            I => \IAC_FLT0\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__30514\,
            I => \IAC_FLT0\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30507\,
            I => \N__30504\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30504\,
            I => \N__30501\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__30501\,
            I => n22374
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__30498\,
            I => \N__30495\
        );

    \I__5292\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__30489\,
            I => n21240
        );

    \I__5289\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__5287\ : Odrv4
    port map (
            O => \N__30480\,
            I => n22401
        );

    \I__5286\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30474\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__5284\ : Span4Mux_h
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__30468\,
            I => n21122
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__30465\,
            I => \n21122_cascade_\
        );

    \I__5281\ : CascadeMux
    port map (
            O => \N__30462\,
            I => \n12610_cascade_\
        );

    \I__5280\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__5278\ : Span4Mux_v
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5277\ : Span4Mux_h
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__30447\,
            I => buf_data_iac_5
        );

    \I__5275\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30441\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__5273\ : Odrv12
    port map (
            O => \N__30438\,
            I => n22_adj_1604
        );

    \I__5272\ : InMux
    port map (
            O => \N__30435\,
            I => n19974
        );

    \I__5271\ : InMux
    port map (
            O => \N__30432\,
            I => n19975
        );

    \I__5270\ : InMux
    port map (
            O => \N__30429\,
            I => n19976
        );

    \I__5269\ : InMux
    port map (
            O => \N__30426\,
            I => n19977
        );

    \I__5268\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30419\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30416\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__30419\,
            I => \N__30413\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__30416\,
            I => secclk_cnt_21
        );

    \I__5264\ : Odrv4
    port map (
            O => \N__30413\,
            I => secclk_cnt_21
        );

    \I__5263\ : InMux
    port map (
            O => \N__30408\,
            I => \N__30404\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30407\,
            I => \N__30401\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__30404\,
            I => secclk_cnt_19
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__30401\,
            I => secclk_cnt_19
        );

    \I__5259\ : CascadeMux
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__5258\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30389\
        );

    \I__5257\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30386\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__30389\,
            I => \N__30383\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__30386\,
            I => secclk_cnt_12
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__30383\,
            I => secclk_cnt_12
        );

    \I__5253\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30374\
        );

    \I__5252\ : InMux
    port map (
            O => \N__30377\,
            I => \N__30371\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__30374\,
            I => secclk_cnt_22
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__30371\,
            I => secclk_cnt_22
        );

    \I__5249\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__30360\,
            I => \N__30356\
        );

    \I__5246\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30353\
        );

    \I__5245\ : Span4Mux_h
    port map (
            O => \N__30356\,
            I => \N__30348\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30348\
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__30348\,
            I => n14_adj_1571
        );

    \I__5242\ : InMux
    port map (
            O => \N__30345\,
            I => n19965
        );

    \I__5241\ : InMux
    port map (
            O => \N__30342\,
            I => n19966
        );

    \I__5240\ : InMux
    port map (
            O => \N__30339\,
            I => n19967
        );

    \I__5239\ : InMux
    port map (
            O => \N__30336\,
            I => n19968
        );

    \I__5238\ : InMux
    port map (
            O => \N__30333\,
            I => n19969
        );

    \I__5237\ : InMux
    port map (
            O => \N__30330\,
            I => n19970
        );

    \I__5236\ : InMux
    port map (
            O => \N__30327\,
            I => \bfn_11_9_0_\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30324\,
            I => n19972
        );

    \I__5234\ : InMux
    port map (
            O => \N__30321\,
            I => n19973
        );

    \I__5233\ : InMux
    port map (
            O => \N__30318\,
            I => n19956
        );

    \I__5232\ : InMux
    port map (
            O => \N__30315\,
            I => n19957
        );

    \I__5231\ : InMux
    port map (
            O => \N__30312\,
            I => n19958
        );

    \I__5230\ : InMux
    port map (
            O => \N__30309\,
            I => n19959
        );

    \I__5229\ : InMux
    port map (
            O => \N__30306\,
            I => n19960
        );

    \I__5228\ : InMux
    port map (
            O => \N__30303\,
            I => n19961
        );

    \I__5227\ : InMux
    port map (
            O => \N__30300\,
            I => n19962
        );

    \I__5226\ : InMux
    port map (
            O => \N__30297\,
            I => \bfn_11_8_0_\
        );

    \I__5225\ : InMux
    port map (
            O => \N__30294\,
            I => n19964
        );

    \I__5224\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30288\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__30288\,
            I => \ADC_VDC.n22587\
        );

    \I__5222\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30282\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__30282\,
            I => \ADC_VDC.n10708\
        );

    \I__5220\ : CascadeMux
    port map (
            O => \N__30279\,
            I => \N__30275\
        );

    \I__5219\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30271\
        );

    \I__5218\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30268\
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30265\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__30271\,
            I => \N__30262\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__30268\,
            I => \N__30259\
        );

    \I__5214\ : InMux
    port map (
            O => \N__30265\,
            I => \N__30256\
        );

    \I__5213\ : Span4Mux_v
    port map (
            O => \N__30262\,
            I => \N__30251\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__30259\,
            I => \N__30251\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__30256\,
            I => cmd_rdadctmp_22_adj_1501
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__30251\,
            I => cmd_rdadctmp_22_adj_1501
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__30246\,
            I => \ADC_VDC.n10708_cascade_\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__5207\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30237\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__30237\,
            I => \N__30233\
        );

    \I__5205\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30230\
        );

    \I__5204\ : Span4Mux_v
    port map (
            O => \N__30233\,
            I => \N__30227\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__30230\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__30227\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__5201\ : SRMux
    port map (
            O => \N__30222\,
            I => \N__30219\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__30216\,
            I => \N__30213\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__30213\,
            I => \ADC_VDC.n5\
        );

    \I__5197\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30206\
        );

    \I__5196\ : InMux
    port map (
            O => \N__30209\,
            I => \N__30203\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__30206\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__30203\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__5193\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30194\
        );

    \I__5192\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30191\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__30194\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__30191\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__30186\,
            I => \N__30182\
        );

    \I__5188\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30179\
        );

    \I__5187\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30176\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__30179\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__30176\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__5184\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30167\
        );

    \I__5183\ : InMux
    port map (
            O => \N__30170\,
            I => \N__30164\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__30167\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__30164\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__5180\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__5178\ : Span4Mux_h
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__30150\,
            I => \ADC_VDC.n20\
        );

    \I__5176\ : CEMux
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__30144\,
            I => \N__30140\
        );

    \I__5174\ : CEMux
    port map (
            O => \N__30143\,
            I => \N__30137\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__30140\,
            I => \N__30132\
        );

    \I__5172\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30132\
        );

    \I__5171\ : Span4Mux_v
    port map (
            O => \N__30132\,
            I => \N__30129\
        );

    \I__5170\ : Span4Mux_v
    port map (
            O => \N__30129\,
            I => \N__30126\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__30126\,
            I => \CLK_DDS.n13005\
        );

    \I__5168\ : CEMux
    port map (
            O => \N__30123\,
            I => \N__30120\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__30120\,
            I => \N__30117\
        );

    \I__5166\ : Odrv12
    port map (
            O => \N__30117\,
            I => \CLK_DDS.n9_adj_1433\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__30114\,
            I => \N__30111\
        );

    \I__5164\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30090\
        );

    \I__5163\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30075\
        );

    \I__5162\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30075\
        );

    \I__5161\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30075\
        );

    \I__5160\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30075\
        );

    \I__5159\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30075\
        );

    \I__5158\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30075\
        );

    \I__5157\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30075\
        );

    \I__5156\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30069\
        );

    \I__5155\ : InMux
    port map (
            O => \N__30102\,
            I => \N__30066\
        );

    \I__5154\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30049\
        );

    \I__5153\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30049\
        );

    \I__5152\ : InMux
    port map (
            O => \N__30099\,
            I => \N__30049\
        );

    \I__5151\ : InMux
    port map (
            O => \N__30098\,
            I => \N__30049\
        );

    \I__5150\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30049\
        );

    \I__5149\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30049\
        );

    \I__5148\ : InMux
    port map (
            O => \N__30095\,
            I => \N__30049\
        );

    \I__5147\ : InMux
    port map (
            O => \N__30094\,
            I => \N__30049\
        );

    \I__5146\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30046\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__30090\,
            I => \N__30042\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__30075\,
            I => \N__30039\
        );

    \I__5143\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30032\
        );

    \I__5142\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30032\
        );

    \I__5141\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30032\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__30069\,
            I => \N__30026\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__30066\,
            I => \N__30026\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__30049\,
            I => \N__30023\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__30046\,
            I => \N__30020\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__30045\,
            I => \N__30017\
        );

    \I__5135\ : Span4Mux_v
    port map (
            O => \N__30042\,
            I => \N__30011\
        );

    \I__5134\ : Span4Mux_v
    port map (
            O => \N__30039\,
            I => \N__30011\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30008\
        );

    \I__5132\ : CascadeMux
    port map (
            O => \N__30031\,
            I => \N__30004\
        );

    \I__5131\ : Span4Mux_v
    port map (
            O => \N__30026\,
            I => \N__30001\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__30023\,
            I => \N__29998\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__30020\,
            I => \N__29995\
        );

    \I__5128\ : InMux
    port map (
            O => \N__30017\,
            I => \N__29990\
        );

    \I__5127\ : InMux
    port map (
            O => \N__30016\,
            I => \N__29990\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__30011\,
            I => \N__29987\
        );

    \I__5125\ : Sp12to4
    port map (
            O => \N__30008\,
            I => \N__29984\
        );

    \I__5124\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29981\
        );

    \I__5123\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29978\
        );

    \I__5122\ : Span4Mux_h
    port map (
            O => \N__30001\,
            I => \N__29973\
        );

    \I__5121\ : Span4Mux_h
    port map (
            O => \N__29998\,
            I => \N__29973\
        );

    \I__5120\ : Span4Mux_h
    port map (
            O => \N__29995\,
            I => \N__29968\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29968\
        );

    \I__5118\ : Sp12to4
    port map (
            O => \N__29987\,
            I => \N__29963\
        );

    \I__5117\ : Span12Mux_v
    port map (
            O => \N__29984\,
            I => \N__29963\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__29981\,
            I => dds_state_2_adj_1494
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29978\,
            I => dds_state_2_adj_1494
        );

    \I__5114\ : Odrv4
    port map (
            O => \N__29973\,
            I => dds_state_2_adj_1494
        );

    \I__5113\ : Odrv4
    port map (
            O => \N__29968\,
            I => dds_state_2_adj_1494
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__29963\,
            I => dds_state_2_adj_1494
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__29952\,
            I => \N__29948\
        );

    \I__5110\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29943\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29934\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29947\,
            I => \N__29934\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29934\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29931\
        );

    \I__5105\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29928\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29925\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29934\,
            I => \N__29922\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__29931\,
            I => \N__29919\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__29928\,
            I => \N__29914\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__29925\,
            I => \N__29914\
        );

    \I__5099\ : Span4Mux_v
    port map (
            O => \N__29922\,
            I => \N__29911\
        );

    \I__5098\ : Span4Mux_h
    port map (
            O => \N__29919\,
            I => \N__29904\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__29914\,
            I => \N__29899\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__29911\,
            I => \N__29899\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29894\
        );

    \I__5094\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29894\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29908\,
            I => \N__29889\
        );

    \I__5092\ : InMux
    port map (
            O => \N__29907\,
            I => \N__29889\
        );

    \I__5091\ : Odrv4
    port map (
            O => \N__29904\,
            I => dds_state_0_adj_1496
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__29899\,
            I => dds_state_0_adj_1496
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__29894\,
            I => dds_state_0_adj_1496
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__29889\,
            I => dds_state_0_adj_1496
        );

    \I__5087\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29855\
        );

    \I__5086\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29855\
        );

    \I__5085\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29855\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29855\
        );

    \I__5083\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29855\
        );

    \I__5082\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29855\
        );

    \I__5081\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29855\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29855\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__29872\,
            I => \N__29848\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29841\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29854\,
            I => \N__29823\
        );

    \I__5076\ : InMux
    port map (
            O => \N__29853\,
            I => \N__29823\
        );

    \I__5075\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29823\
        );

    \I__5074\ : InMux
    port map (
            O => \N__29851\,
            I => \N__29823\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29823\
        );

    \I__5072\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29823\
        );

    \I__5071\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29823\
        );

    \I__5070\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29823\
        );

    \I__5069\ : SRMux
    port map (
            O => \N__29844\,
            I => \N__29816\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__29841\,
            I => \N__29813\
        );

    \I__5067\ : InMux
    port map (
            O => \N__29840\,
            I => \N__29810\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__29823\,
            I => \N__29807\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29804\
        );

    \I__5064\ : CEMux
    port map (
            O => \N__29821\,
            I => \N__29801\
        );

    \I__5063\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29798\
        );

    \I__5062\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29795\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__29816\,
            I => \N__29787\
        );

    \I__5060\ : Span4Mux_v
    port map (
            O => \N__29813\,
            I => \N__29782\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__29810\,
            I => \N__29782\
        );

    \I__5058\ : Span4Mux_v
    port map (
            O => \N__29807\,
            I => \N__29777\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__29804\,
            I => \N__29777\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29801\,
            I => \N__29774\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29798\,
            I => \N__29771\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__29795\,
            I => \N__29768\
        );

    \I__5053\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29760\
        );

    \I__5052\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29760\
        );

    \I__5051\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29760\
        );

    \I__5050\ : InMux
    port map (
            O => \N__29791\,
            I => \N__29755\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29790\,
            I => \N__29755\
        );

    \I__5048\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29750\
        );

    \I__5047\ : Span4Mux_v
    port map (
            O => \N__29782\,
            I => \N__29750\
        );

    \I__5046\ : Span4Mux_v
    port map (
            O => \N__29777\,
            I => \N__29747\
        );

    \I__5045\ : Span4Mux_h
    port map (
            O => \N__29774\,
            I => \N__29742\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__29771\,
            I => \N__29742\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__29768\,
            I => \N__29739\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29736\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__29760\,
            I => \N__29731\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29731\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__29750\,
            I => dds_state_1_adj_1495
        );

    \I__5038\ : Odrv4
    port map (
            O => \N__29747\,
            I => dds_state_1_adj_1495
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__29742\,
            I => dds_state_1_adj_1495
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__29739\,
            I => dds_state_1_adj_1495
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__29736\,
            I => dds_state_1_adj_1495
        );

    \I__5034\ : Odrv12
    port map (
            O => \N__29731\,
            I => dds_state_1_adj_1495
        );

    \I__5033\ : CEMux
    port map (
            O => \N__29718\,
            I => \N__29715\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__29712\,
            I => \N__29708\
        );

    \I__5030\ : CEMux
    port map (
            O => \N__29711\,
            I => \N__29705\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__29708\,
            I => \N__29702\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29699\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__29702\,
            I => \CLK_DDS.n9\
        );

    \I__5026\ : Odrv12
    port map (
            O => \N__29699\,
            I => \CLK_DDS.n9\
        );

    \I__5025\ : InMux
    port map (
            O => \N__29694\,
            I => \bfn_11_7_0_\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__29691\,
            I => \ADC_VDC.n7_cascade_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29688\,
            I => \N__29683\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29687\,
            I => \N__29680\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29686\,
            I => \N__29677\
        );

    \I__5020\ : LocalMux
    port map (
            O => \N__29683\,
            I => \ADC_VDC.n21193\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__29680\,
            I => \ADC_VDC.n21193\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29677\,
            I => \ADC_VDC.n21193\
        );

    \I__5017\ : InMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29667\,
            I => \N__29663\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__29666\,
            I => \N__29660\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__29663\,
            I => \N__29657\
        );

    \I__5013\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29654\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__29657\,
            I => cmd_rdadcbuf_19
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__29654\,
            I => cmd_rdadcbuf_19
        );

    \I__5010\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29646\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__29646\,
            I => \N__29643\
        );

    \I__5008\ : Span4Mux_h
    port map (
            O => \N__29643\,
            I => \N__29639\
        );

    \I__5007\ : InMux
    port map (
            O => \N__29642\,
            I => \N__29636\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__29639\,
            I => cmd_rdadcbuf_24
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__29636\,
            I => cmd_rdadcbuf_24
        );

    \I__5004\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29628\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__29628\,
            I => \N__29625\
        );

    \I__5002\ : Span4Mux_v
    port map (
            O => \N__29625\,
            I => \N__29622\
        );

    \I__5001\ : Span4Mux_v
    port map (
            O => \N__29622\,
            I => \N__29618\
        );

    \I__5000\ : InMux
    port map (
            O => \N__29621\,
            I => \N__29615\
        );

    \I__4999\ : Odrv4
    port map (
            O => \N__29618\,
            I => buf_adcdata_vdc_13
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__29615\,
            I => buf_adcdata_vdc_13
        );

    \I__4997\ : InMux
    port map (
            O => \N__29610\,
            I => \N__29607\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29607\,
            I => \N__29604\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__29604\,
            I => \N__29601\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__29601\,
            I => \N__29597\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29594\
        );

    \I__4992\ : Odrv4
    port map (
            O => \N__29597\,
            I => cmd_rdadcbuf_30
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__29594\,
            I => cmd_rdadcbuf_30
        );

    \I__4990\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29586\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29586\,
            I => \N__29583\
        );

    \I__4988\ : Span12Mux_h
    port map (
            O => \N__29583\,
            I => \N__29579\
        );

    \I__4987\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29576\
        );

    \I__4986\ : Odrv12
    port map (
            O => \N__29579\,
            I => buf_adcdata_vdc_19
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__29576\,
            I => buf_adcdata_vdc_19
        );

    \I__4984\ : InMux
    port map (
            O => \N__29571\,
            I => \N__29568\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__29565\,
            I => \N__29561\
        );

    \I__4981\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29558\
        );

    \I__4980\ : Odrv4
    port map (
            O => \N__29561\,
            I => cmd_rdadcbuf_28
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__29558\,
            I => cmd_rdadcbuf_28
        );

    \I__4978\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29550\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__4976\ : Span4Mux_h
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__4975\ : Span4Mux_v
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4974\ : Sp12to4
    port map (
            O => \N__29541\,
            I => \N__29537\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29534\
        );

    \I__4972\ : Odrv12
    port map (
            O => \N__29537\,
            I => buf_adcdata_vdc_17
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__29534\,
            I => buf_adcdata_vdc_17
        );

    \I__4970\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__29520\,
            I => \N__29516\
        );

    \I__4966\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29513\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__29516\,
            I => cmd_rdadcbuf_32
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__29513\,
            I => cmd_rdadcbuf_32
        );

    \I__4963\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__29502\,
            I => \N__29498\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__29501\,
            I => \N__29495\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__29498\,
            I => \N__29492\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29489\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__29492\,
            I => buf_adcdata_vdc_21
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__29489\,
            I => buf_adcdata_vdc_21
        );

    \I__4955\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__4953\ : Span4Mux_h
    port map (
            O => \N__29478\,
            I => \N__29475\
        );

    \I__4952\ : Span4Mux_v
    port map (
            O => \N__29475\,
            I => \N__29471\
        );

    \I__4951\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29468\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__29471\,
            I => cmd_rdadcbuf_31
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29468\,
            I => cmd_rdadcbuf_31
        );

    \I__4948\ : InMux
    port map (
            O => \N__29463\,
            I => \N__29460\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__29457\,
            I => \N__29453\
        );

    \I__4945\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29449\
        );

    \I__4944\ : Span4Mux_h
    port map (
            O => \N__29453\,
            I => \N__29446\
        );

    \I__4943\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29443\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__29449\,
            I => \N__29440\
        );

    \I__4941\ : Span4Mux_v
    port map (
            O => \N__29446\,
            I => \N__29437\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__29443\,
            I => buf_dds1_4
        );

    \I__4939\ : Odrv4
    port map (
            O => \N__29440\,
            I => buf_dds1_4
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__29437\,
            I => buf_dds1_4
        );

    \I__4937\ : CascadeMux
    port map (
            O => \N__29430\,
            I => \N__29425\
        );

    \I__4936\ : CascadeMux
    port map (
            O => \N__29429\,
            I => \N__29422\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__29428\,
            I => \N__29419\
        );

    \I__4934\ : InMux
    port map (
            O => \N__29425\,
            I => \N__29416\
        );

    \I__4933\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29413\
        );

    \I__4932\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29410\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__29416\,
            I => \N__29407\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__29413\,
            I => \N__29402\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__29410\,
            I => \N__29402\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__29407\,
            I => \N__29399\
        );

    \I__4927\ : Odrv4
    port map (
            O => \N__29402\,
            I => cmd_rdadctmp_20
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__29399\,
            I => cmd_rdadctmp_20
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__29394\,
            I => \N__29387\
        );

    \I__4924\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29375\
        );

    \I__4923\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29375\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__29391\,
            I => \N__29369\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__29390\,
            I => \N__29366\
        );

    \I__4920\ : InMux
    port map (
            O => \N__29387\,
            I => \N__29357\
        );

    \I__4919\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29357\
        );

    \I__4918\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29354\
        );

    \I__4917\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29349\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29349\
        );

    \I__4915\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29344\
        );

    \I__4914\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29344\
        );

    \I__4913\ : InMux
    port map (
            O => \N__29380\,
            I => \N__29341\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__29375\,
            I => \N__29338\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__29374\,
            I => \N__29329\
        );

    \I__4910\ : InMux
    port map (
            O => \N__29373\,
            I => \N__29320\
        );

    \I__4909\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29313\
        );

    \I__4908\ : InMux
    port map (
            O => \N__29369\,
            I => \N__29313\
        );

    \I__4907\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29313\
        );

    \I__4906\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29308\
        );

    \I__4905\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29308\
        );

    \I__4904\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29303\
        );

    \I__4903\ : InMux
    port map (
            O => \N__29362\,
            I => \N__29303\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__29357\,
            I => \N__29298\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__29354\,
            I => \N__29298\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__29349\,
            I => \N__29295\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29292\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__29341\,
            I => \N__29287\
        );

    \I__4897\ : Span4Mux_v
    port map (
            O => \N__29338\,
            I => \N__29287\
        );

    \I__4896\ : InMux
    port map (
            O => \N__29337\,
            I => \N__29284\
        );

    \I__4895\ : InMux
    port map (
            O => \N__29336\,
            I => \N__29277\
        );

    \I__4894\ : InMux
    port map (
            O => \N__29335\,
            I => \N__29277\
        );

    \I__4893\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29277\
        );

    \I__4892\ : InMux
    port map (
            O => \N__29333\,
            I => \N__29272\
        );

    \I__4891\ : InMux
    port map (
            O => \N__29332\,
            I => \N__29272\
        );

    \I__4890\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29263\
        );

    \I__4889\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29263\
        );

    \I__4888\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29263\
        );

    \I__4887\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29263\
        );

    \I__4886\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29256\
        );

    \I__4885\ : InMux
    port map (
            O => \N__29324\,
            I => \N__29256\
        );

    \I__4884\ : InMux
    port map (
            O => \N__29323\,
            I => \N__29256\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__29320\,
            I => \N__29249\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__29313\,
            I => \N__29249\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29249\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__29303\,
            I => \N__29246\
        );

    \I__4879\ : Span4Mux_h
    port map (
            O => \N__29298\,
            I => \N__29241\
        );

    \I__4878\ : Span4Mux_v
    port map (
            O => \N__29295\,
            I => \N__29241\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__29292\,
            I => \N__29236\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__29287\,
            I => \N__29236\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__29284\,
            I => n12771
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__29277\,
            I => n12771
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__29272\,
            I => n12771
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__29263\,
            I => n12771
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__29256\,
            I => n12771
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__29249\,
            I => n12771
        );

    \I__4869\ : Odrv12
    port map (
            O => \N__29246\,
            I => n12771
        );

    \I__4868\ : Odrv4
    port map (
            O => \N__29241\,
            I => n12771
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__29236\,
            I => n12771
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__29217\,
            I => \N__29214\
        );

    \I__4865\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29210\
        );

    \I__4864\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__29210\,
            I => cmd_rdadctmp_31
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__29207\,
            I => cmd_rdadctmp_31
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__29202\,
            I => \N__29198\
        );

    \I__4860\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29195\
        );

    \I__4859\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29192\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29189\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__29192\,
            I => \N__29185\
        );

    \I__4856\ : Span12Mux_h
    port map (
            O => \N__29189\,
            I => \N__29182\
        );

    \I__4855\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29179\
        );

    \I__4854\ : Span4Mux_v
    port map (
            O => \N__29185\,
            I => \N__29176\
        );

    \I__4853\ : Span12Mux_v
    port map (
            O => \N__29182\,
            I => \N__29173\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__29179\,
            I => buf_adcdata_iac_23
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__29176\,
            I => buf_adcdata_iac_23
        );

    \I__4850\ : Odrv12
    port map (
            O => \N__29173\,
            I => buf_adcdata_iac_23
        );

    \I__4849\ : CEMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29160\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__29160\,
            I => \N__29157\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__29157\,
            I => \ADC_VDC.n16\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__29154\,
            I => \ADC_VDC.n21593_cascade_\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__29151\,
            I => \ADC_VDC.n21590_cascade_\
        );

    \I__4843\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__29145\,
            I => \ADC_VDC.n22590\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__29142\,
            I => \N__29131\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__29141\,
            I => \N__29128\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__29140\,
            I => \N__29125\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__29139\,
            I => \N__29122\
        );

    \I__4837\ : CascadeMux
    port map (
            O => \N__29138\,
            I => \N__29119\
        );

    \I__4836\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29097\
        );

    \I__4835\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29097\
        );

    \I__4834\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29097\
        );

    \I__4833\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29097\
        );

    \I__4832\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29097\
        );

    \I__4831\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29097\
        );

    \I__4830\ : InMux
    port map (
            O => \N__29125\,
            I => \N__29097\
        );

    \I__4829\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29097\
        );

    \I__4828\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29094\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__29118\,
            I => \N__29088\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__29117\,
            I => \N__29085\
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__29116\,
            I => \N__29077\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__29115\,
            I => \N__29074\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__29114\,
            I => \N__29071\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__29097\,
            I => \N__29067\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__29094\,
            I => \N__29064\
        );

    \I__4820\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29047\
        );

    \I__4819\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29047\
        );

    \I__4818\ : InMux
    port map (
            O => \N__29091\,
            I => \N__29047\
        );

    \I__4817\ : InMux
    port map (
            O => \N__29088\,
            I => \N__29047\
        );

    \I__4816\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29047\
        );

    \I__4815\ : InMux
    port map (
            O => \N__29084\,
            I => \N__29047\
        );

    \I__4814\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29047\
        );

    \I__4813\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29047\
        );

    \I__4812\ : InMux
    port map (
            O => \N__29081\,
            I => \N__29034\
        );

    \I__4811\ : InMux
    port map (
            O => \N__29080\,
            I => \N__29034\
        );

    \I__4810\ : InMux
    port map (
            O => \N__29077\,
            I => \N__29034\
        );

    \I__4809\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29034\
        );

    \I__4808\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29034\
        );

    \I__4807\ : InMux
    port map (
            O => \N__29070\,
            I => \N__29034\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__29067\,
            I => \N__29031\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__29064\,
            I => \N__29028\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__29047\,
            I => \N__29023\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__29034\,
            I => \N__29023\
        );

    \I__4802\ : Sp12to4
    port map (
            O => \N__29031\,
            I => \N__29020\
        );

    \I__4801\ : Span4Mux_v
    port map (
            O => \N__29028\,
            I => \N__29017\
        );

    \I__4800\ : Span4Mux_h
    port map (
            O => \N__29023\,
            I => \N__29014\
        );

    \I__4799\ : Odrv12
    port map (
            O => \N__29020\,
            I => n13324
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__29017\,
            I => n13324
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__29014\,
            I => n13324
        );

    \I__4796\ : IoInMux
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__29004\,
            I => \N__29001\
        );

    \I__4794\ : Span4Mux_s1_h
    port map (
            O => \N__29001\,
            I => \N__28998\
        );

    \I__4793\ : Sp12to4
    port map (
            O => \N__28998\,
            I => \N__28995\
        );

    \I__4792\ : Span12Mux_s5_v
    port map (
            O => \N__28995\,
            I => \N__28991\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28987\
        );

    \I__4790\ : Span12Mux_h
    port map (
            O => \N__28991\,
            I => \N__28984\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28981\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28987\,
            I => \N__28978\
        );

    \I__4787\ : Odrv12
    port map (
            O => \N__28984\,
            I => \VAC_FLT1\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__28981\,
            I => \VAC_FLT1\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28978\,
            I => \VAC_FLT1\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__28971\,
            I => \N__28968\
        );

    \I__4783\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28965\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28965\,
            I => \N__28962\
        );

    \I__4781\ : Span4Mux_h
    port map (
            O => \N__28962\,
            I => \N__28957\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28952\
        );

    \I__4779\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28952\
        );

    \I__4778\ : Odrv4
    port map (
            O => \N__28957\,
            I => cmd_rdadctmp_29
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28952\,
            I => cmd_rdadctmp_29
        );

    \I__4776\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28944\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__4774\ : Span4Mux_h
    port map (
            O => \N__28941\,
            I => \N__28937\
        );

    \I__4773\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28934\
        );

    \I__4772\ : Sp12to4
    port map (
            O => \N__28937\,
            I => \N__28930\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__28934\,
            I => \N__28927\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28924\
        );

    \I__4769\ : Span12Mux_v
    port map (
            O => \N__28930\,
            I => \N__28921\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__28927\,
            I => \N__28918\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28924\,
            I => buf_adcdata_iac_21
        );

    \I__4766\ : Odrv12
    port map (
            O => \N__28921\,
            I => buf_adcdata_iac_21
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__28918\,
            I => buf_adcdata_iac_21
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__28911\,
            I => \N__28908\
        );

    \I__4763\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28904\
        );

    \I__4762\ : CascadeMux
    port map (
            O => \N__28907\,
            I => \N__28901\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__28904\,
            I => \N__28897\
        );

    \I__4760\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28892\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28892\
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__28897\,
            I => cmd_rdadctmp_28
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__28892\,
            I => cmd_rdadctmp_28
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__28887\,
            I => \N__28883\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__28886\,
            I => \N__28880\
        );

    \I__4754\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28876\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28873\
        );

    \I__4752\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28870\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28876\,
            I => cmd_rdadctmp_25
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__28873\,
            I => cmd_rdadctmp_25
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__28870\,
            I => cmd_rdadctmp_25
        );

    \I__4748\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28859\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28856\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__28859\,
            I => n17728
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28856\,
            I => n17728
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__28851\,
            I => \n11_cascade_\
        );

    \I__4743\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28843\
        );

    \I__4742\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28840\
        );

    \I__4741\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28836\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28843\,
            I => \N__28833\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__28840\,
            I => \N__28830\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28827\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28823\
        );

    \I__4736\ : Span4Mux_h
    port map (
            O => \N__28833\,
            I => \N__28816\
        );

    \I__4735\ : Span4Mux_v
    port map (
            O => \N__28830\,
            I => \N__28816\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__28827\,
            I => \N__28816\
        );

    \I__4733\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28813\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__28823\,
            I => acadc_dtrig_v
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__28816\,
            I => acadc_dtrig_v
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28813\,
            I => acadc_dtrig_v
        );

    \I__4729\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28803\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28798\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28795\
        );

    \I__4726\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28792\
        );

    \I__4725\ : Span4Mux_v
    port map (
            O => \N__28798\,
            I => \N__28787\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28787\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28782\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__28787\,
            I => \N__28779\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28774\
        );

    \I__4720\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28774\
        );

    \I__4719\ : Span4Mux_v
    port map (
            O => \N__28782\,
            I => \N__28771\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__28779\,
            I => acadc_dtrig_i
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__28774\,
            I => acadc_dtrig_i
        );

    \I__4716\ : Odrv4
    port map (
            O => \N__28771\,
            I => acadc_dtrig_i
        );

    \I__4715\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28761\,
            I => \eis_state_2_N_392_1\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__28758\,
            I => \eis_state_2_N_392_1_cascade_\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__28755\,
            I => \n2_adj_1696_cascade_\
        );

    \I__4711\ : InMux
    port map (
            O => \N__28752\,
            I => \N__28749\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__28749\,
            I => n22437
        );

    \I__4709\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28742\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28745\,
            I => \N__28739\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__28742\,
            I => \N__28735\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__28739\,
            I => \N__28732\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28729\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__28735\,
            I => cmd_rdadctmp_23
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__28732\,
            I => cmd_rdadctmp_23
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__28729\,
            I => cmd_rdadctmp_23
        );

    \I__4701\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__28719\,
            I => n22371
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__28716\,
            I => \n12_adj_1454_cascade_\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__28710\,
            I => \N__28705\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28709\,
            I => \N__28702\
        );

    \I__4695\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28699\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__28705\,
            I => \N__28692\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__28702\,
            I => \N__28692\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__28699\,
            I => \N__28689\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28686\
        );

    \I__4690\ : InMux
    port map (
            O => \N__28697\,
            I => \N__28683\
        );

    \I__4689\ : Span4Mux_h
    port map (
            O => \N__28692\,
            I => \N__28680\
        );

    \I__4688\ : Span4Mux_v
    port map (
            O => \N__28689\,
            I => \N__28677\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__28686\,
            I => \N__28674\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__28683\,
            I => acadc_trig
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__28680\,
            I => acadc_trig
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__28677\,
            I => acadc_trig
        );

    \I__4683\ : Odrv12
    port map (
            O => \N__28674\,
            I => acadc_trig
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__28665\,
            I => \N__28661\
        );

    \I__4681\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28658\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28655\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__28658\,
            I => n21053
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__28655\,
            I => n21053
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__28650\,
            I => \n21042_cascade_\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__28647\,
            I => \n21030_cascade_\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28640\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28637\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28640\,
            I => eis_end
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__28637\,
            I => eis_end
        );

    \I__4671\ : SRMux
    port map (
            O => \N__28632\,
            I => \N__28628\
        );

    \I__4670\ : SRMux
    port map (
            O => \N__28631\,
            I => \N__28623\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28618\
        );

    \I__4668\ : SRMux
    port map (
            O => \N__28627\,
            I => \N__28615\
        );

    \I__4667\ : SRMux
    port map (
            O => \N__28626\,
            I => \N__28611\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28607\
        );

    \I__4665\ : SRMux
    port map (
            O => \N__28622\,
            I => \N__28604\
        );

    \I__4664\ : SRMux
    port map (
            O => \N__28621\,
            I => \N__28599\
        );

    \I__4663\ : Span4Mux_h
    port map (
            O => \N__28618\,
            I => \N__28596\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__28615\,
            I => \N__28593\
        );

    \I__4661\ : SRMux
    port map (
            O => \N__28614\,
            I => \N__28590\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__28611\,
            I => \N__28587\
        );

    \I__4659\ : SRMux
    port map (
            O => \N__28610\,
            I => \N__28584\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__28607\,
            I => \N__28579\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__28604\,
            I => \N__28579\
        );

    \I__4656\ : SRMux
    port map (
            O => \N__28603\,
            I => \N__28576\
        );

    \I__4655\ : SRMux
    port map (
            O => \N__28602\,
            I => \N__28572\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28568\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__28596\,
            I => \N__28563\
        );

    \I__4652\ : Span4Mux_h
    port map (
            O => \N__28593\,
            I => \N__28563\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__28590\,
            I => \N__28560\
        );

    \I__4650\ : Span4Mux_v
    port map (
            O => \N__28587\,
            I => \N__28555\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__28584\,
            I => \N__28555\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__28579\,
            I => \N__28550\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__28576\,
            I => \N__28550\
        );

    \I__4646\ : SRMux
    port map (
            O => \N__28575\,
            I => \N__28547\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28544\
        );

    \I__4644\ : SRMux
    port map (
            O => \N__28571\,
            I => \N__28541\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__28568\,
            I => \N__28538\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__28563\,
            I => \N__28533\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__28560\,
            I => \N__28533\
        );

    \I__4640\ : Span4Mux_v
    port map (
            O => \N__28555\,
            I => \N__28528\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__28550\,
            I => \N__28528\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__28547\,
            I => \N__28525\
        );

    \I__4637\ : Span4Mux_v
    port map (
            O => \N__28544\,
            I => \N__28520\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28541\,
            I => \N__28520\
        );

    \I__4635\ : Span4Mux_v
    port map (
            O => \N__28538\,
            I => \N__28511\
        );

    \I__4634\ : Span4Mux_v
    port map (
            O => \N__28533\,
            I => \N__28511\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__28528\,
            I => \N__28511\
        );

    \I__4632\ : Span4Mux_h
    port map (
            O => \N__28525\,
            I => \N__28511\
        );

    \I__4631\ : Sp12to4
    port map (
            O => \N__28520\,
            I => \N__28508\
        );

    \I__4630\ : Span4Mux_h
    port map (
            O => \N__28511\,
            I => \N__28505\
        );

    \I__4629\ : Span12Mux_v
    port map (
            O => \N__28508\,
            I => \N__28502\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__28505\,
            I => \N__28499\
        );

    \I__4627\ : Odrv12
    port map (
            O => \N__28502\,
            I => \iac_raw_buf_N_774\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__28499\,
            I => \iac_raw_buf_N_774\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28494\,
            I => \N__28491\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__28491\,
            I => n21334
        );

    \I__4623\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__28485\,
            I => n22512
        );

    \I__4621\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28478\
        );

    \I__4620\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28475\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__28478\,
            I => \N__28472\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__28475\,
            I => data_idxvec_15
        );

    \I__4617\ : Odrv4
    port map (
            O => \N__28472\,
            I => data_idxvec_15
        );

    \I__4616\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__28464\,
            I => \N__28461\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__4613\ : Span4Mux_h
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__4612\ : Sp12to4
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__4611\ : Span12Mux_v
    port map (
            O => \N__28452\,
            I => \N__28449\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__28449\,
            I => buf_data_iac_23
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__28446\,
            I => \n26_adj_1659_cascade_\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__28443\,
            I => \n21324_cascade_\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28437\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__4605\ : Span4Mux_h
    port map (
            O => \N__28434\,
            I => \N__28429\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28426\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__28432\,
            I => \N__28423\
        );

    \I__4602\ : Span4Mux_h
    port map (
            O => \N__28429\,
            I => \N__28418\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__28426\,
            I => \N__28418\
        );

    \I__4600\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28415\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__28418\,
            I => \N__28412\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__28415\,
            I => buf_adcdata_vac_15
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__28412\,
            I => buf_adcdata_vac_15
        );

    \I__4596\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__28404\,
            I => \N__28400\
        );

    \I__4594\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28397\
        );

    \I__4593\ : Span4Mux_v
    port map (
            O => \N__28400\,
            I => \N__28392\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__28397\,
            I => \N__28392\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__28392\,
            I => buf_adcdata_vdc_15
        );

    \I__4590\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28386\,
            I => \N__28383\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__4587\ : Odrv4
    port map (
            O => \N__28380\,
            I => n19_adj_1621
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__28377\,
            I => \N__28374\
        );

    \I__4585\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28371\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__4583\ : Odrv12
    port map (
            O => \N__28368\,
            I => n23_adj_1658
        );

    \I__4582\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28362\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__28362\,
            I => n21323
        );

    \I__4580\ : InMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__4578\ : Span4Mux_h
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__28350\,
            I => n19_adj_1652
        );

    \I__4576\ : CascadeMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28338\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__28338\,
            I => \N__28334\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__28337\,
            I => \N__28331\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__28334\,
            I => \N__28328\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28331\,
            I => \N__28325\
        );

    \I__4569\ : Odrv4
    port map (
            O => \N__28328\,
            I => \buf_readRTD_1\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__28325\,
            I => \buf_readRTD_1\
        );

    \I__4567\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28317\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__28317\,
            I => \N__28314\
        );

    \I__4565\ : Sp12to4
    port map (
            O => \N__28314\,
            I => \N__28309\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__28313\,
            I => \N__28306\
        );

    \I__4563\ : InMux
    port map (
            O => \N__28312\,
            I => \N__28303\
        );

    \I__4562\ : Span12Mux_v
    port map (
            O => \N__28309\,
            I => \N__28300\
        );

    \I__4561\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28297\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__28303\,
            I => \N__28292\
        );

    \I__4559\ : Span12Mux_h
    port map (
            O => \N__28300\,
            I => \N__28292\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__28297\,
            I => buf_adcdata_vac_13
        );

    \I__4557\ : Odrv12
    port map (
            O => \N__28292\,
            I => buf_adcdata_vac_13
        );

    \I__4556\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28284\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__28284\,
            I => \N__28280\
        );

    \I__4554\ : InMux
    port map (
            O => \N__28283\,
            I => \N__28277\
        );

    \I__4553\ : Odrv12
    port map (
            O => \N__28280\,
            I => \buf_readRTD_5\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__28277\,
            I => \buf_readRTD_5\
        );

    \I__4551\ : CascadeMux
    port map (
            O => \N__28272\,
            I => \n19_adj_1629_cascade_\
        );

    \I__4550\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28262\
        );

    \I__4549\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28257\
        );

    \I__4548\ : InMux
    port map (
            O => \N__28267\,
            I => \N__28257\
        );

    \I__4547\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28251\
        );

    \I__4546\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28248\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__28262\,
            I => \N__28241\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28234\
        );

    \I__4543\ : InMux
    port map (
            O => \N__28256\,
            I => \N__28227\
        );

    \I__4542\ : InMux
    port map (
            O => \N__28255\,
            I => \N__28227\
        );

    \I__4541\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28227\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28224\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__28248\,
            I => \N__28221\
        );

    \I__4538\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28216\
        );

    \I__4537\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28216\
        );

    \I__4536\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28205\
        );

    \I__4535\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28205\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__28241\,
            I => \N__28202\
        );

    \I__4533\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28195\
        );

    \I__4532\ : InMux
    port map (
            O => \N__28239\,
            I => \N__28195\
        );

    \I__4531\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28195\
        );

    \I__4530\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28192\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__28234\,
            I => \N__28180\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28180\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__28224\,
            I => \N__28173\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__28221\,
            I => \N__28173\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28173\
        );

    \I__4524\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28160\
        );

    \I__4523\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28160\
        );

    \I__4522\ : InMux
    port map (
            O => \N__28213\,
            I => \N__28160\
        );

    \I__4521\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28160\
        );

    \I__4520\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28160\
        );

    \I__4519\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28160\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__28205\,
            I => \N__28157\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__28202\,
            I => \N__28150\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__28195\,
            I => \N__28150\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__28192\,
            I => \N__28150\
        );

    \I__4514\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28145\
        );

    \I__4513\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28145\
        );

    \I__4512\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28138\
        );

    \I__4511\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28138\
        );

    \I__4510\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28138\
        );

    \I__4509\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28133\
        );

    \I__4508\ : InMux
    port map (
            O => \N__28185\,
            I => \N__28133\
        );

    \I__4507\ : Span4Mux_v
    port map (
            O => \N__28180\,
            I => \N__28127\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__28173\,
            I => \N__28122\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__28160\,
            I => \N__28122\
        );

    \I__4504\ : Span4Mux_v
    port map (
            O => \N__28157\,
            I => \N__28117\
        );

    \I__4503\ : Span4Mux_h
    port map (
            O => \N__28150\,
            I => \N__28117\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__28145\,
            I => \N__28112\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__28138\,
            I => \N__28112\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28109\
        );

    \I__4499\ : InMux
    port map (
            O => \N__28132\,
            I => \N__28102\
        );

    \I__4498\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28102\
        );

    \I__4497\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28102\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__28127\,
            I => n12850
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__28122\,
            I => n12850
        );

    \I__4494\ : Odrv4
    port map (
            O => \N__28117\,
            I => n12850
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__28112\,
            I => n12850
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__28109\,
            I => n12850
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__28102\,
            I => n12850
        );

    \I__4490\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28085\
        );

    \I__4489\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28082\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__28085\,
            I => \N__28079\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__28082\,
            I => \N__28075\
        );

    \I__4486\ : Span4Mux_v
    port map (
            O => \N__28079\,
            I => \N__28072\
        );

    \I__4485\ : InMux
    port map (
            O => \N__28078\,
            I => \N__28069\
        );

    \I__4484\ : Odrv12
    port map (
            O => \N__28075\,
            I => cmd_rdadctmp_21_adj_1471
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__28072\,
            I => cmd_rdadctmp_21_adj_1471
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__28069\,
            I => cmd_rdadctmp_21_adj_1471
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__4480\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28056\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__28053\,
            I => n8
        );

    \I__4477\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__28047\,
            I => \N__28043\
        );

    \I__4475\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28040\
        );

    \I__4474\ : Span4Mux_v
    port map (
            O => \N__28043\,
            I => \N__28035\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__28040\,
            I => \N__28035\
        );

    \I__4472\ : Span4Mux_v
    port map (
            O => \N__28035\,
            I => \N__28031\
        );

    \I__4471\ : InMux
    port map (
            O => \N__28034\,
            I => \N__28028\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__28031\,
            I => n10695
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__28028\,
            I => n10695
        );

    \I__4468\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__28020\,
            I => \N__28016\
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__28019\,
            I => \N__28013\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__28010\
        );

    \I__4464\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28007\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__28010\,
            I => buf_adcdata_vdc_12
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__28007\,
            I => buf_adcdata_vdc_12
        );

    \I__4461\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27992\
        );

    \I__4460\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27992\
        );

    \I__4459\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27985\
        );

    \I__4458\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27982\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27998\,
            I => \N__27968\
        );

    \I__4456\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27968\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27992\,
            I => \N__27961\
        );

    \I__4454\ : InMux
    port map (
            O => \N__27991\,
            I => \N__27952\
        );

    \I__4453\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27952\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27952\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27952\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__27985\,
            I => \N__27947\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27982\,
            I => \N__27947\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27940\
        );

    \I__4447\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27940\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27940\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27937\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27928\
        );

    \I__4443\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27928\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27928\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27974\,
            I => \N__27928\
        );

    \I__4440\ : InMux
    port map (
            O => \N__27973\,
            I => \N__27925\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27922\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27917\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27917\
        );

    \I__4436\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27914\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__27964\,
            I => \N__27911\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__27961\,
            I => \N__27906\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__27952\,
            I => \N__27906\
        );

    \I__4432\ : Span4Mux_v
    port map (
            O => \N__27947\,
            I => \N__27899\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27899\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27937\,
            I => \N__27899\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__27928\,
            I => \N__27894\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27925\,
            I => \N__27894\
        );

    \I__4427\ : Span4Mux_v
    port map (
            O => \N__27922\,
            I => \N__27887\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27917\,
            I => \N__27887\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__27914\,
            I => \N__27887\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27884\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__27906\,
            I => \N__27880\
        );

    \I__4422\ : Span4Mux_h
    port map (
            O => \N__27899\,
            I => \N__27877\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__27894\,
            I => \N__27870\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__27887\,
            I => \N__27870\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27884\,
            I => \N__27870\
        );

    \I__4418\ : InMux
    port map (
            O => \N__27883\,
            I => \N__27867\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__27880\,
            I => n21076
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__27877\,
            I => n21076
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__27870\,
            I => n21076
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__27867\,
            I => n21076
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__27858\,
            I => \N__27852\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__27857\,
            I => \N__27844\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__27856\,
            I => \N__27836\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__27855\,
            I => \N__27828\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27852\,
            I => \N__27817\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27812\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27812\
        );

    \I__4406\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27807\
        );

    \I__4405\ : InMux
    port map (
            O => \N__27848\,
            I => \N__27807\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__27847\,
            I => \N__27797\
        );

    \I__4403\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27787\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27784\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27842\,
            I => \N__27779\
        );

    \I__4400\ : InMux
    port map (
            O => \N__27841\,
            I => \N__27779\
        );

    \I__4399\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27773\
        );

    \I__4398\ : InMux
    port map (
            O => \N__27839\,
            I => \N__27773\
        );

    \I__4397\ : InMux
    port map (
            O => \N__27836\,
            I => \N__27760\
        );

    \I__4396\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27760\
        );

    \I__4395\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27760\
        );

    \I__4394\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27760\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27760\
        );

    \I__4392\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27760\
        );

    \I__4391\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27752\
        );

    \I__4390\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27747\
        );

    \I__4389\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27747\
        );

    \I__4388\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27742\
        );

    \I__4387\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27742\
        );

    \I__4386\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27733\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27733\
        );

    \I__4384\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27733\
        );

    \I__4383\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27733\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__27817\,
            I => \N__27726\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__27812\,
            I => \N__27726\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__27807\,
            I => \N__27726\
        );

    \I__4379\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27708\
        );

    \I__4378\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27708\
        );

    \I__4377\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27708\
        );

    \I__4376\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27708\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27708\
        );

    \I__4374\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27708\
        );

    \I__4373\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27705\
        );

    \I__4372\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27700\
        );

    \I__4371\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27700\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27687\
        );

    \I__4369\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27687\
        );

    \I__4368\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27687\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27792\,
            I => \N__27687\
        );

    \I__4366\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27687\
        );

    \I__4365\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27687\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__27787\,
            I => \N__27684\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27679\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27679\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27676\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__27773\,
            I => \N__27671\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__27760\,
            I => \N__27671\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__27759\,
            I => \N__27665\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__27758\,
            I => \N__27662\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__27757\,
            I => \N__27659\
        );

    \I__4355\ : CascadeMux
    port map (
            O => \N__27756\,
            I => \N__27652\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__27755\,
            I => \N__27647\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__27752\,
            I => \N__27639\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__27747\,
            I => \N__27639\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27632\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__27733\,
            I => \N__27632\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__27726\,
            I => \N__27632\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27621\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27621\
        );

    \I__4346\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27621\
        );

    \I__4345\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27616\
        );

    \I__4344\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27616\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__27708\,
            I => \N__27613\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__27705\,
            I => \N__27610\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27601\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27687\,
            I => \N__27601\
        );

    \I__4339\ : Span4Mux_h
    port map (
            O => \N__27684\,
            I => \N__27601\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__27679\,
            I => \N__27601\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__27676\,
            I => \N__27596\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__27671\,
            I => \N__27596\
        );

    \I__4335\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27589\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27589\
        );

    \I__4333\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27589\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27574\
        );

    \I__4331\ : InMux
    port map (
            O => \N__27662\,
            I => \N__27574\
        );

    \I__4330\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27574\
        );

    \I__4329\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27574\
        );

    \I__4328\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27574\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27574\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27574\
        );

    \I__4325\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27571\
        );

    \I__4324\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27566\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27566\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27557\
        );

    \I__4321\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27557\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27557\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27557\
        );

    \I__4318\ : Span4Mux_v
    port map (
            O => \N__27639\,
            I => \N__27552\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__27632\,
            I => \N__27552\
        );

    \I__4316\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27543\
        );

    \I__4315\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27543\
        );

    \I__4314\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27543\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27543\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27526\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__27616\,
            I => \N__27526\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__27613\,
            I => \N__27526\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__27610\,
            I => \N__27526\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__27601\,
            I => \N__27526\
        );

    \I__4307\ : Span4Mux_h
    port map (
            O => \N__27596\,
            I => \N__27526\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__27589\,
            I => \N__27526\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27526\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__27571\,
            I => adc_state_0_adj_1460
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__27566\,
            I => adc_state_0_adj_1460
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__27557\,
            I => adc_state_0_adj_1460
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__27552\,
            I => adc_state_0_adj_1460
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__27543\,
            I => adc_state_0_adj_1460
        );

    \I__4299\ : Odrv4
    port map (
            O => \N__27526\,
            I => adc_state_0_adj_1460
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__27513\,
            I => \N__27509\
        );

    \I__4297\ : InMux
    port map (
            O => \N__27512\,
            I => \N__27504\
        );

    \I__4296\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27504\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__27501\,
            I => \N__27497\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27500\,
            I => \N__27494\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__27497\,
            I => \N__27489\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__27494\,
            I => \N__27489\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__27489\,
            I => cmd_rdadctmp_20_adj_1472
        );

    \I__4289\ : InMux
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27483\,
            I => \N__27478\
        );

    \I__4287\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27473\
        );

    \I__4286\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27473\
        );

    \I__4285\ : Span12Mux_v
    port map (
            O => \N__27478\,
            I => \N__27470\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__27473\,
            I => buf_adcdata_vac_12
        );

    \I__4283\ : Odrv12
    port map (
            O => \N__27470\,
            I => buf_adcdata_vac_12
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__27465\,
            I => \N__27462\
        );

    \I__4281\ : InMux
    port map (
            O => \N__27462\,
            I => \N__27459\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27459\,
            I => \N__27455\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27458\,
            I => \N__27452\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__27455\,
            I => \N__27449\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__27452\,
            I => \N__27446\
        );

    \I__4276\ : Span4Mux_v
    port map (
            O => \N__27449\,
            I => \N__27442\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__27446\,
            I => \N__27439\
        );

    \I__4274\ : InMux
    port map (
            O => \N__27445\,
            I => \N__27436\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__27442\,
            I => cmd_rdadctmp_19_adj_1473
        );

    \I__4272\ : Odrv4
    port map (
            O => \N__27439\,
            I => cmd_rdadctmp_19_adj_1473
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__27436\,
            I => cmd_rdadctmp_19_adj_1473
        );

    \I__4270\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27426\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27426\,
            I => \N__27422\
        );

    \I__4268\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27418\
        );

    \I__4267\ : Span4Mux_v
    port map (
            O => \N__27422\,
            I => \N__27415\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__27421\,
            I => \N__27412\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27409\
        );

    \I__4264\ : Sp12to4
    port map (
            O => \N__27415\,
            I => \N__27406\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27403\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__27409\,
            I => \N__27400\
        );

    \I__4261\ : Span12Mux_h
    port map (
            O => \N__27406\,
            I => \N__27397\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27403\,
            I => buf_adcdata_vac_21
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__27400\,
            I => buf_adcdata_vac_21
        );

    \I__4258\ : Odrv12
    port map (
            O => \N__27397\,
            I => buf_adcdata_vac_21
        );

    \I__4257\ : IoInMux
    port map (
            O => \N__27390\,
            I => \N__27387\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27384\
        );

    \I__4255\ : IoSpan4Mux
    port map (
            O => \N__27384\,
            I => \N__27380\
        );

    \I__4254\ : InMux
    port map (
            O => \N__27383\,
            I => \N__27377\
        );

    \I__4253\ : Sp12to4
    port map (
            O => \N__27380\,
            I => \N__27374\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__27377\,
            I => \N__27370\
        );

    \I__4251\ : Span12Mux_h
    port map (
            O => \N__27374\,
            I => \N__27367\
        );

    \I__4250\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27364\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__27370\,
            I => \N__27361\
        );

    \I__4248\ : Odrv12
    port map (
            O => \N__27367\,
            I => \VAC_OSR1\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__27364\,
            I => \VAC_OSR1\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__27361\,
            I => \VAC_OSR1\
        );

    \I__4245\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27351\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__27351\,
            I => \N__27347\
        );

    \I__4243\ : CascadeMux
    port map (
            O => \N__27350\,
            I => \N__27344\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__27347\,
            I => \N__27341\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27338\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__27341\,
            I => buf_adcdata_vdc_10
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__27338\,
            I => buf_adcdata_vdc_10
        );

    \I__4238\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27326\
        );

    \I__4236\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27322\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__27326\,
            I => \N__27319\
        );

    \I__4234\ : CascadeMux
    port map (
            O => \N__27325\,
            I => \N__27316\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__27322\,
            I => \N__27313\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__27319\,
            I => \N__27310\
        );

    \I__4231\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27307\
        );

    \I__4230\ : Span4Mux_h
    port map (
            O => \N__27313\,
            I => \N__27304\
        );

    \I__4229\ : Sp12to4
    port map (
            O => \N__27310\,
            I => \N__27301\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__27307\,
            I => buf_adcdata_vac_10
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__27304\,
            I => buf_adcdata_vac_10
        );

    \I__4226\ : Odrv12
    port map (
            O => \N__27301\,
            I => buf_adcdata_vac_10
        );

    \I__4225\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27290\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__27293\,
            I => \N__27287\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27290\,
            I => \N__27284\
        );

    \I__4222\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27281\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__27284\,
            I => \N__27276\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27276\
        );

    \I__4219\ : Odrv4
    port map (
            O => \N__27276\,
            I => buf_adcdata_vdc_0
        );

    \I__4218\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27269\
        );

    \I__4217\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27266\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__27269\,
            I => \N__27263\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27260\
        );

    \I__4214\ : Span12Mux_s11_h
    port map (
            O => \N__27263\,
            I => \N__27256\
        );

    \I__4213\ : Span4Mux_v
    port map (
            O => \N__27260\,
            I => \N__27253\
        );

    \I__4212\ : InMux
    port map (
            O => \N__27259\,
            I => \N__27250\
        );

    \I__4211\ : Span12Mux_h
    port map (
            O => \N__27256\,
            I => \N__27247\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__27253\,
            I => \N__27244\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__27250\,
            I => buf_adcdata_vac_0
        );

    \I__4208\ : Odrv12
    port map (
            O => \N__27247\,
            I => buf_adcdata_vac_0
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__27244\,
            I => buf_adcdata_vac_0
        );

    \I__4206\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4204\ : Span4Mux_v
    port map (
            O => \N__27231\,
            I => \N__27227\
        );

    \I__4203\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27224\
        );

    \I__4202\ : Sp12to4
    port map (
            O => \N__27227\,
            I => \N__27220\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__27224\,
            I => \N__27217\
        );

    \I__4200\ : InMux
    port map (
            O => \N__27223\,
            I => \N__27214\
        );

    \I__4199\ : Span12Mux_h
    port map (
            O => \N__27220\,
            I => \N__27211\
        );

    \I__4198\ : Span4Mux_h
    port map (
            O => \N__27217\,
            I => \N__27208\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__27214\,
            I => buf_adcdata_iac_0
        );

    \I__4196\ : Odrv12
    port map (
            O => \N__27211\,
            I => buf_adcdata_iac_0
        );

    \I__4195\ : Odrv4
    port map (
            O => \N__27208\,
            I => buf_adcdata_iac_0
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__27201\,
            I => \n19_adj_1534_cascade_\
        );

    \I__4193\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27195\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__4191\ : Odrv12
    port map (
            O => \N__27192\,
            I => buf_control_7
        );

    \I__4190\ : IoInMux
    port map (
            O => \N__27189\,
            I => \N__27186\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4188\ : Span4Mux_s3_v
    port map (
            O => \N__27183\,
            I => \N__27180\
        );

    \I__4187\ : Sp12to4
    port map (
            O => \N__27180\,
            I => \N__27176\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__27179\,
            I => \N__27173\
        );

    \I__4185\ : Span12Mux_h
    port map (
            O => \N__27176\,
            I => \N__27170\
        );

    \I__4184\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27167\
        );

    \I__4183\ : Odrv12
    port map (
            O => \N__27170\,
            I => \DDS_SCK1\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__27167\,
            I => \DDS_SCK1\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__27162\,
            I => \N__27159\
        );

    \I__4180\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__27156\,
            I => \N__27153\
        );

    \I__4178\ : Span4Mux_h
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__27150\,
            I => \N__27146\
        );

    \I__4176\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27143\
        );

    \I__4175\ : Odrv4
    port map (
            O => \N__27146\,
            I => \buf_readRTD_15\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__27143\,
            I => \buf_readRTD_15\
        );

    \I__4173\ : CascadeMux
    port map (
            O => \N__27138\,
            I => \N__27134\
        );

    \I__4172\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27131\
        );

    \I__4171\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27128\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__27131\,
            I => buf_adcdata_vdc_23
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__27128\,
            I => buf_adcdata_vdc_23
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__27123\,
            I => \n22593_cascade_\
        );

    \I__4167\ : InMux
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27114\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__27114\,
            I => \N__27110\
        );

    \I__4164\ : InMux
    port map (
            O => \N__27113\,
            I => \N__27107\
        );

    \I__4163\ : Sp12to4
    port map (
            O => \N__27110\,
            I => \N__27104\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27101\
        );

    \I__4161\ : Span12Mux_v
    port map (
            O => \N__27104\,
            I => \N__27097\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__27101\,
            I => \N__27094\
        );

    \I__4159\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27091\
        );

    \I__4158\ : Span12Mux_h
    port map (
            O => \N__27097\,
            I => \N__27088\
        );

    \I__4157\ : Span4Mux_h
    port map (
            O => \N__27094\,
            I => \N__27085\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__27091\,
            I => buf_adcdata_vac_23
        );

    \I__4155\ : Odrv12
    port map (
            O => \N__27088\,
            I => buf_adcdata_vac_23
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__27085\,
            I => buf_adcdata_vac_23
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__27078\,
            I => \N__27074\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__27077\,
            I => \N__27071\
        );

    \I__4151\ : InMux
    port map (
            O => \N__27074\,
            I => \N__27067\
        );

    \I__4150\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27064\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__27070\,
            I => \N__27061\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__27067\,
            I => \N__27057\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__27064\,
            I => \N__27054\
        );

    \I__4146\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27050\
        );

    \I__4145\ : InMux
    port map (
            O => \N__27060\,
            I => \N__27047\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__27057\,
            I => \N__27044\
        );

    \I__4143\ : Span4Mux_v
    port map (
            O => \N__27054\,
            I => \N__27041\
        );

    \I__4142\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27038\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__27050\,
            I => \N__27033\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__27047\,
            I => \N__27033\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__27044\,
            I => \buf_cfgRTD_6\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__27041\,
            I => \buf_cfgRTD_6\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__27038\,
            I => \buf_cfgRTD_6\
        );

    \I__4136\ : Odrv12
    port map (
            O => \N__27033\,
            I => \buf_cfgRTD_6\
        );

    \I__4135\ : CascadeMux
    port map (
            O => \N__27024\,
            I => \N__27021\
        );

    \I__4134\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__27011\
        );

    \I__4132\ : InMux
    port map (
            O => \N__27017\,
            I => \N__27006\
        );

    \I__4131\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27006\
        );

    \I__4130\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27001\
        );

    \I__4129\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27001\
        );

    \I__4128\ : Span4Mux_v
    port map (
            O => \N__27011\,
            I => \N__26998\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__27006\,
            I => \N__26995\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__27001\,
            I => \N__26992\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__26998\,
            I => \buf_cfgRTD_7\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__26995\,
            I => \buf_cfgRTD_7\
        );

    \I__4123\ : Odrv4
    port map (
            O => \N__26992\,
            I => \buf_cfgRTD_7\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__26985\,
            I => \N__26982\
        );

    \I__4121\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26979\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__26979\,
            I => n30_adj_1499
        );

    \I__4119\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26972\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26969\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26972\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__26969\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__4115\ : InMux
    port map (
            O => \N__26964\,
            I => \ADC_VDC.n19886\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26961\,
            I => \ADC_VDC.n19887\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26954\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26951\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26954\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__26951\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__4109\ : CEMux
    port map (
            O => \N__26946\,
            I => \N__26942\
        );

    \I__4108\ : CEMux
    port map (
            O => \N__26945\,
            I => \N__26937\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26942\,
            I => \N__26934\
        );

    \I__4106\ : CEMux
    port map (
            O => \N__26941\,
            I => \N__26931\
        );

    \I__4105\ : CEMux
    port map (
            O => \N__26940\,
            I => \N__26926\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26923\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__26934\,
            I => \N__26918\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26931\,
            I => \N__26918\
        );

    \I__4101\ : CEMux
    port map (
            O => \N__26930\,
            I => \N__26915\
        );

    \I__4100\ : CEMux
    port map (
            O => \N__26929\,
            I => \N__26912\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__26926\,
            I => \N__26909\
        );

    \I__4098\ : Span4Mux_v
    port map (
            O => \N__26923\,
            I => \N__26901\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__26918\,
            I => \N__26901\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__26915\,
            I => \N__26901\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26912\,
            I => \N__26897\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__26909\,
            I => \N__26894\
        );

    \I__4093\ : CEMux
    port map (
            O => \N__26908\,
            I => \N__26891\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__26901\,
            I => \N__26888\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26885\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__26897\,
            I => \N__26880\
        );

    \I__4089\ : Span4Mux_h
    port map (
            O => \N__26894\,
            I => \N__26880\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26891\,
            I => \N__26873\
        );

    \I__4087\ : Span4Mux_h
    port map (
            O => \N__26888\,
            I => \N__26873\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__26885\,
            I => \N__26873\
        );

    \I__4085\ : Odrv4
    port map (
            O => \N__26880\,
            I => \ADC_VDC.n13463\
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__26873\,
            I => \ADC_VDC.n13463\
        );

    \I__4083\ : SRMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26865\,
            I => \N__26860\
        );

    \I__4081\ : SRMux
    port map (
            O => \N__26864\,
            I => \N__26857\
        );

    \I__4080\ : SRMux
    port map (
            O => \N__26863\,
            I => \N__26850\
        );

    \I__4079\ : Span4Mux_h
    port map (
            O => \N__26860\,
            I => \N__26845\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__26857\,
            I => \N__26845\
        );

    \I__4077\ : SRMux
    port map (
            O => \N__26856\,
            I => \N__26842\
        );

    \I__4076\ : SRMux
    port map (
            O => \N__26855\,
            I => \N__26839\
        );

    \I__4075\ : SRMux
    port map (
            O => \N__26854\,
            I => \N__26836\
        );

    \I__4074\ : SRMux
    port map (
            O => \N__26853\,
            I => \N__26833\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26830\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__26845\,
            I => \N__26827\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__26842\,
            I => \N__26824\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__26839\,
            I => \N__26819\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__26836\,
            I => \N__26819\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__26833\,
            I => \N__26816\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__26830\,
            I => \N__26813\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__26827\,
            I => \N__26810\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__26824\,
            I => \N__26805\
        );

    \I__4064\ : Span4Mux_v
    port map (
            O => \N__26819\,
            I => \N__26805\
        );

    \I__4063\ : Odrv12
    port map (
            O => \N__26816\,
            I => \ADC_VDC.n15175\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__26813\,
            I => \ADC_VDC.n15175\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__26810\,
            I => \ADC_VDC.n15175\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26805\,
            I => \ADC_VDC.n15175\
        );

    \I__4059\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__26793\,
            I => \N__26789\
        );

    \I__4057\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26786\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__26789\,
            I => cmd_rdadcbuf_23
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__26786\,
            I => cmd_rdadcbuf_23
        );

    \I__4054\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26778\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26778\,
            I => \N__26774\
        );

    \I__4052\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26771\
        );

    \I__4051\ : Odrv4
    port map (
            O => \N__26774\,
            I => cmd_rdadcbuf_18
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__26771\,
            I => cmd_rdadcbuf_18
        );

    \I__4049\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26760\
        );

    \I__4047\ : Span12Mux_v
    port map (
            O => \N__26760\,
            I => \N__26756\
        );

    \I__4046\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26753\
        );

    \I__4045\ : Odrv12
    port map (
            O => \N__26756\,
            I => buf_adcdata_vdc_7
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__26753\,
            I => buf_adcdata_vdc_7
        );

    \I__4043\ : CascadeMux
    port map (
            O => \N__26748\,
            I => \n11891_cascade_\
        );

    \I__4042\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26739\
        );

    \I__4040\ : Span4Mux_h
    port map (
            O => \N__26739\,
            I => \N__26735\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26732\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__26735\,
            I => cmd_rdadcbuf_26
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__26732\,
            I => cmd_rdadcbuf_26
        );

    \I__4036\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26724\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26721\
        );

    \I__4034\ : Span4Mux_v
    port map (
            O => \N__26721\,
            I => \N__26717\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26714\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__26717\,
            I => cmd_rdadcbuf_25
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__26714\,
            I => cmd_rdadcbuf_25
        );

    \I__4030\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26706\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__26706\,
            I => \N__26702\
        );

    \I__4028\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26699\
        );

    \I__4027\ : Odrv12
    port map (
            O => \N__26702\,
            I => cmd_rdadcbuf_22
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__26699\,
            I => cmd_rdadcbuf_22
        );

    \I__4025\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26691\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__26691\,
            I => \N__26687\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26684\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__26687\,
            I => \N__26681\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__26684\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__26681\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__4019\ : InMux
    port map (
            O => \N__26676\,
            I => \ADC_VDC.n19877\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__26673\,
            I => \N__26670\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26666\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26663\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__26666\,
            I => \N__26660\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__26663\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__26660\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__4012\ : InMux
    port map (
            O => \N__26655\,
            I => \ADC_VDC.n19878\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26652\,
            I => \ADC_VDC.n19879\
        );

    \I__4010\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26645\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26642\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__26645\,
            I => \N__26639\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__26642\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__26639\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26634\,
            I => \ADC_VDC.n19880\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__26631\,
            I => \N__26627\
        );

    \I__4003\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26624\
        );

    \I__4002\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26621\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__26624\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__26621\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26616\,
            I => \ADC_VDC.n19881\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26613\,
            I => \ADC_VDC.n19882\
        );

    \I__3997\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26606\
        );

    \I__3996\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26603\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__26606\,
            I => \N__26600\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26603\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__26600\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26595\,
            I => \ADC_VDC.n19883\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26592\,
            I => \bfn_10_7_0_\
        );

    \I__3990\ : InMux
    port map (
            O => \N__26589\,
            I => \ADC_VDC.n19885\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__26586\,
            I => \N__26581\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26578\
        );

    \I__3987\ : InMux
    port map (
            O => \N__26584\,
            I => \N__26575\
        );

    \I__3986\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26572\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26578\,
            I => cmd_rdadctmp_30
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__26575\,
            I => cmd_rdadctmp_30
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__26572\,
            I => cmd_rdadctmp_30
        );

    \I__3982\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26562\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__26562\,
            I => \N__26559\
        );

    \I__3980\ : Span4Mux_v
    port map (
            O => \N__26559\,
            I => \N__26556\
        );

    \I__3979\ : Odrv4
    port map (
            O => \N__26556\,
            I => \ADC_VDC.n18780\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__26553\,
            I => \ADC_VDC.n18783_cascade_\
        );

    \I__3977\ : CEMux
    port map (
            O => \N__26550\,
            I => \N__26547\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__26547\,
            I => \ADC_VDC.n16_adj_1450\
        );

    \I__3975\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26541\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__26541\,
            I => \ADC_VDC.n18\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__26538\,
            I => \ADC_VDC.n18_cascade_\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26532\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26529\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__26529\,
            I => \N__26526\
        );

    \I__3969\ : Sp12to4
    port map (
            O => \N__26526\,
            I => \N__26523\
        );

    \I__3968\ : Span12Mux_v
    port map (
            O => \N__26523\,
            I => \N__26520\
        );

    \I__3967\ : Odrv12
    port map (
            O => \N__26520\,
            I => \THERMOSTAT\
        );

    \I__3966\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26513\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26510\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__26513\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__26510\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__3962\ : InMux
    port map (
            O => \N__26505\,
            I => \bfn_10_6_0_\
        );

    \I__3961\ : IoInMux
    port map (
            O => \N__26502\,
            I => \N__26499\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26499\,
            I => \N__26496\
        );

    \I__3959\ : IoSpan4Mux
    port map (
            O => \N__26496\,
            I => \N__26493\
        );

    \I__3958\ : Span4Mux_s1_v
    port map (
            O => \N__26493\,
            I => \N__26490\
        );

    \I__3957\ : Span4Mux_v
    port map (
            O => \N__26490\,
            I => \N__26487\
        );

    \I__3956\ : Span4Mux_v
    port map (
            O => \N__26487\,
            I => \N__26482\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26477\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26477\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__26482\,
            I => \IAC_FLT1\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26477\,
            I => \IAC_FLT1\
        );

    \I__3951\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26469\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__3949\ : Span12Mux_v
    port map (
            O => \N__26466\,
            I => \N__26462\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__26465\,
            I => \N__26458\
        );

    \I__3947\ : Span12Mux_h
    port map (
            O => \N__26462\,
            I => \N__26455\
        );

    \I__3946\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26450\
        );

    \I__3945\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26450\
        );

    \I__3944\ : Odrv12
    port map (
            O => \N__26455\,
            I => buf_adcdata_iac_19
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__26450\,
            I => buf_adcdata_iac_19
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__26445\,
            I => \n22605_cascade_\
        );

    \I__3941\ : InMux
    port map (
            O => \N__26442\,
            I => \N__26438\
        );

    \I__3940\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26435\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__26438\,
            I => \N__26432\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__26435\,
            I => \N__26426\
        );

    \I__3937\ : Span4Mux_v
    port map (
            O => \N__26432\,
            I => \N__26426\
        );

    \I__3936\ : InMux
    port map (
            O => \N__26431\,
            I => \N__26423\
        );

    \I__3935\ : Odrv4
    port map (
            O => \N__26426\,
            I => buf_dds1_11
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__26423\,
            I => buf_dds1_11
        );

    \I__3933\ : InMux
    port map (
            O => \N__26418\,
            I => \N__26415\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26412\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__26412\,
            I => n22608
        );

    \I__3930\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26405\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__26408\,
            I => \N__26402\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__26405\,
            I => \N__26398\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26395\
        );

    \I__3926\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26392\
        );

    \I__3925\ : Odrv4
    port map (
            O => \N__26398\,
            I => cmd_rdadctmp_27
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__26395\,
            I => cmd_rdadctmp_27
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__26392\,
            I => cmd_rdadctmp_27
        );

    \I__3922\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26380\
        );

    \I__3921\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26375\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26375\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__26380\,
            I => cmd_rdadctmp_19
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__26375\,
            I => cmd_rdadctmp_19
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__26370\,
            I => \N__26366\
        );

    \I__3916\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26358\
        );

    \I__3915\ : InMux
    port map (
            O => \N__26366\,
            I => \N__26358\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26358\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__26358\,
            I => cmd_rdadctmp_24
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__26355\,
            I => \N__26351\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__26354\,
            I => \N__26348\
        );

    \I__3910\ : InMux
    port map (
            O => \N__26351\,
            I => \N__26342\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26342\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__26347\,
            I => \N__26339\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__26342\,
            I => \N__26336\
        );

    \I__3906\ : InMux
    port map (
            O => \N__26339\,
            I => \N__26333\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__26336\,
            I => cmd_rdadctmp_22_adj_1470
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26333\,
            I => cmd_rdadctmp_22_adj_1470
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__26328\,
            I => \N__26324\
        );

    \I__3902\ : InMux
    port map (
            O => \N__26327\,
            I => \N__26316\
        );

    \I__3901\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26316\
        );

    \I__3900\ : InMux
    port map (
            O => \N__26323\,
            I => \N__26316\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__26316\,
            I => cmd_rdadctmp_23_adj_1469
        );

    \I__3898\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26310\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26307\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__26307\,
            I => \N__26304\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__26304\,
            I => n69
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__26301\,
            I => \N__26297\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__26300\,
            I => \N__26294\
        );

    \I__3892\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26291\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26288\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__26291\,
            I => \N__26285\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26282\
        );

    \I__3888\ : Span4Mux_v
    port map (
            O => \N__26285\,
            I => \N__26278\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__26282\,
            I => \N__26275\
        );

    \I__3886\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26272\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__26278\,
            I => cmd_rdadctmp_15
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__26275\,
            I => cmd_rdadctmp_15
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__26272\,
            I => cmd_rdadctmp_15
        );

    \I__3882\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26260\
        );

    \I__3881\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26255\
        );

    \I__3880\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26255\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__26260\,
            I => buf_dds1_2
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__26255\,
            I => buf_dds1_2
        );

    \I__3877\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26247\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26244\
        );

    \I__3875\ : Span4Mux_v
    port map (
            O => \N__26244\,
            I => \N__26241\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__26241\,
            I => n22476
        );

    \I__3873\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26235\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__26235\,
            I => \N__26231\
        );

    \I__3871\ : CascadeMux
    port map (
            O => \N__26234\,
            I => \N__26228\
        );

    \I__3870\ : Span4Mux_h
    port map (
            O => \N__26231\,
            I => \N__26225\
        );

    \I__3869\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26222\
        );

    \I__3868\ : Sp12to4
    port map (
            O => \N__26225\,
            I => \N__26216\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__26222\,
            I => \N__26216\
        );

    \I__3866\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26213\
        );

    \I__3865\ : Odrv12
    port map (
            O => \N__26216\,
            I => cmd_rdadctmp_16_adj_1476
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__26213\,
            I => cmd_rdadctmp_16_adj_1476
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__26208\,
            I => \N__26204\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__26207\,
            I => \N__26201\
        );

    \I__3861\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26198\
        );

    \I__3860\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26195\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__26198\,
            I => \N__26189\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__26195\,
            I => \N__26189\
        );

    \I__3857\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26186\
        );

    \I__3856\ : Odrv12
    port map (
            O => \N__26189\,
            I => cmd_rdadctmp_25_adj_1467
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__26186\,
            I => cmd_rdadctmp_25_adj_1467
        );

    \I__3854\ : InMux
    port map (
            O => \N__26181\,
            I => \N__26178\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__26178\,
            I => \N__26175\
        );

    \I__3852\ : Span4Mux_h
    port map (
            O => \N__26175\,
            I => \N__26170\
        );

    \I__3851\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26165\
        );

    \I__3850\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26165\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__26170\,
            I => cmd_rdadctmp_24_adj_1468
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__26165\,
            I => cmd_rdadctmp_24_adj_1468
        );

    \I__3847\ : CEMux
    port map (
            O => \N__26160\,
            I => \N__26157\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26153\
        );

    \I__3845\ : CEMux
    port map (
            O => \N__26156\,
            I => \N__26150\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__26153\,
            I => \N__26147\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__26150\,
            I => \N__26142\
        );

    \I__3842\ : Span4Mux_v
    port map (
            O => \N__26147\,
            I => \N__26142\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__26142\,
            I => n12493
        );

    \I__3840\ : InMux
    port map (
            O => \N__26139\,
            I => \N__26136\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__26136\,
            I => \N__26133\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__26133\,
            I => \N__26130\
        );

    \I__3837\ : Odrv4
    port map (
            O => \N__26130\,
            I => n21705
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__26127\,
            I => \N__26123\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__26126\,
            I => \N__26119\
        );

    \I__3834\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26116\
        );

    \I__3833\ : InMux
    port map (
            O => \N__26122\,
            I => \N__26113\
        );

    \I__3832\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26110\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__26116\,
            I => \N__26107\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__26113\,
            I => cmd_rdadctmp_18_adj_1474
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__26110\,
            I => cmd_rdadctmp_18_adj_1474
        );

    \I__3828\ : Odrv12
    port map (
            O => \N__26107\,
            I => cmd_rdadctmp_18_adj_1474
        );

    \I__3827\ : IoInMux
    port map (
            O => \N__26100\,
            I => \N__26097\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__26097\,
            I => \N__26094\
        );

    \I__3825\ : IoSpan4Mux
    port map (
            O => \N__26094\,
            I => \N__26091\
        );

    \I__3824\ : IoSpan4Mux
    port map (
            O => \N__26091\,
            I => \N__26087\
        );

    \I__3823\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26084\
        );

    \I__3822\ : Sp12to4
    port map (
            O => \N__26087\,
            I => \N__26081\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__26084\,
            I => \N__26077\
        );

    \I__3820\ : Span12Mux_s6_v
    port map (
            O => \N__26081\,
            I => \N__26074\
        );

    \I__3819\ : InMux
    port map (
            O => \N__26080\,
            I => \N__26071\
        );

    \I__3818\ : Span4Mux_v
    port map (
            O => \N__26077\,
            I => \N__26068\
        );

    \I__3817\ : Odrv12
    port map (
            O => \N__26074\,
            I => \IAC_OSR1\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__26071\,
            I => \IAC_OSR1\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__26068\,
            I => \IAC_OSR1\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__26061\,
            I => \N__26057\
        );

    \I__3813\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26054\
        );

    \I__3812\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26051\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__26054\,
            I => \N__26048\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__26051\,
            I => data_idxvec_11
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__26048\,
            I => data_idxvec_11
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__26043\,
            I => \n26_adj_1678_cascade_\
        );

    \I__3807\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26037\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__26037\,
            I => n22509
        );

    \I__3805\ : InMux
    port map (
            O => \N__26034\,
            I => \bfn_9_12_0_\
        );

    \I__3804\ : InMux
    port map (
            O => \N__26031\,
            I => n19821
        );

    \I__3803\ : InMux
    port map (
            O => \N__26028\,
            I => n19822
        );

    \I__3802\ : InMux
    port map (
            O => \N__26025\,
            I => n19823
        );

    \I__3801\ : InMux
    port map (
            O => \N__26022\,
            I => n19824
        );

    \I__3800\ : InMux
    port map (
            O => \N__26019\,
            I => n19825
        );

    \I__3799\ : InMux
    port map (
            O => \N__26016\,
            I => n19826
        );

    \I__3798\ : InMux
    port map (
            O => \N__26013\,
            I => n19827
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__26010\,
            I => \N__26007\
        );

    \I__3796\ : InMux
    port map (
            O => \N__26007\,
            I => \N__26004\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__26004\,
            I => \N__26000\
        );

    \I__3794\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25997\
        );

    \I__3793\ : Span4Mux_v
    port map (
            O => \N__26000\,
            I => \N__25993\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25997\,
            I => \N__25990\
        );

    \I__3791\ : InMux
    port map (
            O => \N__25996\,
            I => \N__25987\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__25993\,
            I => cmd_rdadctmp_27_adj_1465
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__25990\,
            I => cmd_rdadctmp_27_adj_1465
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25987\,
            I => cmd_rdadctmp_27_adj_1465
        );

    \I__3787\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25977\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25977\,
            I => \N__25974\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__25974\,
            I => \N__25971\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__25971\,
            I => \N__25966\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25963\
        );

    \I__3782\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25960\
        );

    \I__3781\ : Sp12to4
    port map (
            O => \N__25966\,
            I => \N__25957\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__25963\,
            I => \N__25954\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25960\,
            I => buf_adcdata_vac_19
        );

    \I__3778\ : Odrv12
    port map (
            O => \N__25957\,
            I => buf_adcdata_vac_19
        );

    \I__3777\ : Odrv12
    port map (
            O => \N__25954\,
            I => buf_adcdata_vac_19
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__25947\,
            I => \N__25943\
        );

    \I__3775\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25939\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25934\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25942\,
            I => \N__25934\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25939\,
            I => \N__25929\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__25934\,
            I => \N__25929\
        );

    \I__3770\ : Span4Mux_v
    port map (
            O => \N__25929\,
            I => \N__25924\
        );

    \I__3769\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25919\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25919\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__25924\,
            I => \buf_cfgRTD_3\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__25919\,
            I => \buf_cfgRTD_3\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__25914\,
            I => \N__25911\
        );

    \I__3764\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25908\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__25908\,
            I => \N__25904\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25901\
        );

    \I__3761\ : Odrv12
    port map (
            O => \N__25904\,
            I => \buf_readRTD_11\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__25901\,
            I => \buf_readRTD_11\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25896\,
            I => \N__25893\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__25893\,
            I => \N__25890\
        );

    \I__3757\ : Odrv12
    port map (
            O => \N__25890\,
            I => n22473
        );

    \I__3756\ : InMux
    port map (
            O => \N__25887\,
            I => \bfn_9_11_0_\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25884\,
            I => n19813
        );

    \I__3754\ : InMux
    port map (
            O => \N__25881\,
            I => n19814
        );

    \I__3753\ : InMux
    port map (
            O => \N__25878\,
            I => n19815
        );

    \I__3752\ : InMux
    port map (
            O => \N__25875\,
            I => n19816
        );

    \I__3751\ : InMux
    port map (
            O => \N__25872\,
            I => n19817
        );

    \I__3750\ : InMux
    port map (
            O => \N__25869\,
            I => n19818
        );

    \I__3749\ : InMux
    port map (
            O => \N__25866\,
            I => n19819
        );

    \I__3748\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25858\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25855\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25852\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__25858\,
            I => cmd_rdadcbuf_34
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25855\,
            I => cmd_rdadcbuf_34
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__25852\,
            I => cmd_rdadcbuf_34
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__25845\,
            I => \ADC_VDC.n18780_cascade_\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__25842\,
            I => \N__25839\
        );

    \I__3740\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25836\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__25836\,
            I => \ADC_VDC.n4_adj_1451\
        );

    \I__3738\ : CEMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__25827\,
            I => \ADC_VDC.n13503\
        );

    \I__3735\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__3733\ : Span4Mux_h
    port map (
            O => \N__25818\,
            I => \N__25814\
        );

    \I__3732\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25811\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__25814\,
            I => \buf_readRTD_8\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__25811\,
            I => \buf_readRTD_8\
        );

    \I__3729\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25803\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__3727\ : Span4Mux_v
    port map (
            O => \N__25800\,
            I => \N__25796\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__25799\,
            I => \N__25793\
        );

    \I__3725\ : Span4Mux_v
    port map (
            O => \N__25796\,
            I => \N__25790\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25787\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__25790\,
            I => buf_adcdata_vdc_16
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__25787\,
            I => buf_adcdata_vdc_16
        );

    \I__3721\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25779\,
            I => \N__25775\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25772\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__25775\,
            I => \N__25769\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__25772\,
            I => \N__25766\
        );

    \I__3716\ : Span4Mux_h
    port map (
            O => \N__25769\,
            I => \N__25763\
        );

    \I__3715\ : Span4Mux_h
    port map (
            O => \N__25766\,
            I => \N__25759\
        );

    \I__3714\ : Span4Mux_h
    port map (
            O => \N__25763\,
            I => \N__25756\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25753\
        );

    \I__3712\ : Span4Mux_v
    port map (
            O => \N__25759\,
            I => \N__25748\
        );

    \I__3711\ : Span4Mux_h
    port map (
            O => \N__25756\,
            I => \N__25748\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__25753\,
            I => buf_adcdata_vac_16
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__25748\,
            I => buf_adcdata_vac_16
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__25743\,
            I => \n22575_cascade_\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__25740\,
            I => \N__25736\
        );

    \I__3706\ : InMux
    port map (
            O => \N__25739\,
            I => \N__25732\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25729\
        );

    \I__3704\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25726\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25723\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25729\,
            I => \N__25720\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__25726\,
            I => \N__25717\
        );

    \I__3700\ : Span12Mux_h
    port map (
            O => \N__25723\,
            I => \N__25712\
        );

    \I__3699\ : Span4Mux_h
    port map (
            O => \N__25720\,
            I => \N__25709\
        );

    \I__3698\ : Span4Mux_h
    port map (
            O => \N__25717\,
            I => \N__25706\
        );

    \I__3697\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25701\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25715\,
            I => \N__25701\
        );

    \I__3695\ : Odrv12
    port map (
            O => \N__25712\,
            I => \buf_cfgRTD_0\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__25709\,
            I => \buf_cfgRTD_0\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__25706\,
            I => \buf_cfgRTD_0\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__25701\,
            I => \buf_cfgRTD_0\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__25692\,
            I => \n10902_cascade_\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__25689\,
            I => \n12624_cascade_\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__25686\,
            I => \N__25683\
        );

    \I__3688\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25680\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__3686\ : Span4Mux_v
    port map (
            O => \N__25677\,
            I => \N__25673\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__25676\,
            I => \N__25670\
        );

    \I__3684\ : Span4Mux_h
    port map (
            O => \N__25673\,
            I => \N__25667\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25664\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__25667\,
            I => buf_adcdata_vdc_22
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__25664\,
            I => buf_adcdata_vdc_22
        );

    \I__3680\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25655\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25652\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__25655\,
            I => cmd_rdadcbuf_13
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__25652\,
            I => cmd_rdadcbuf_13
        );

    \I__3676\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__25644\,
            I => \N__25640\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__3673\ : Span4Mux_h
    port map (
            O => \N__25640\,
            I => \N__25634\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25637\,
            I => \N__25631\
        );

    \I__3671\ : Sp12to4
    port map (
            O => \N__25634\,
            I => \N__25628\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__25631\,
            I => \N__25625\
        );

    \I__3669\ : Odrv12
    port map (
            O => \N__25628\,
            I => buf_adcdata_vdc_2
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__25625\,
            I => buf_adcdata_vdc_2
        );

    \I__3667\ : InMux
    port map (
            O => \N__25620\,
            I => \N__25616\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25613\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25616\,
            I => cmd_rdadcbuf_15
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__25613\,
            I => cmd_rdadcbuf_15
        );

    \I__3663\ : InMux
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__25605\,
            I => \N__25601\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__25604\,
            I => \N__25598\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__25601\,
            I => \N__25595\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25592\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__25595\,
            I => buf_adcdata_vdc_4
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__25592\,
            I => buf_adcdata_vdc_4
        );

    \I__3656\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25583\
        );

    \I__3655\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25580\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__25583\,
            I => cmd_rdadcbuf_16
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25580\,
            I => cmd_rdadcbuf_16
        );

    \I__3652\ : InMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__25572\,
            I => \N__25568\
        );

    \I__3650\ : CascadeMux
    port map (
            O => \N__25571\,
            I => \N__25565\
        );

    \I__3649\ : Span4Mux_v
    port map (
            O => \N__25568\,
            I => \N__25562\
        );

    \I__3648\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25559\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__25562\,
            I => buf_adcdata_vdc_5
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__25559\,
            I => buf_adcdata_vdc_5
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__25554\,
            I => \N__25550\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25546\
        );

    \I__3643\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25543\
        );

    \I__3642\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25540\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__25546\,
            I => \N__25535\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25543\,
            I => \N__25535\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__25540\,
            I => cmd_rdadctmp_20_adj_1503
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__25535\,
            I => cmd_rdadctmp_20_adj_1503
        );

    \I__3637\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25526\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__25529\,
            I => \N__25522\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__25526\,
            I => \N__25519\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25525\,
            I => \N__25516\
        );

    \I__3633\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25513\
        );

    \I__3632\ : Odrv12
    port map (
            O => \N__25519\,
            I => cmd_rdadctmp_21_adj_1502
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__25516\,
            I => cmd_rdadctmp_21_adj_1502
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25513\,
            I => cmd_rdadctmp_21_adj_1502
        );

    \I__3629\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__25503\,
            I => \ADC_VDC.cmd_rdadcbuf_35_N_1296_34\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__25497\,
            I => \N__25494\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__25494\,
            I => \ADC_VDC.n19\
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__25491\,
            I => \ADC_VDC.n21_cascade_\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__25488\,
            I => \N__25483\
        );

    \I__3622\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25478\
        );

    \I__3621\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25478\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25475\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25478\,
            I => cmd_rdadctmp_14_adj_1509
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25475\,
            I => cmd_rdadctmp_14_adj_1509
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__25470\,
            I => \N__25465\
        );

    \I__3616\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25462\
        );

    \I__3615\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25459\
        );

    \I__3614\ : InMux
    port map (
            O => \N__25465\,
            I => \N__25456\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25462\,
            I => cmd_rdadctmp_15_adj_1508
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__25459\,
            I => cmd_rdadctmp_15_adj_1508
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__25456\,
            I => cmd_rdadctmp_15_adj_1508
        );

    \I__3610\ : InMux
    port map (
            O => \N__25449\,
            I => \N__25445\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25448\,
            I => \N__25442\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__25445\,
            I => cmd_rdadcbuf_20
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__25442\,
            I => cmd_rdadcbuf_20
        );

    \I__3606\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25434\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__3604\ : Span4Mux_v
    port map (
            O => \N__25431\,
            I => \N__25427\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25430\,
            I => \N__25424\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__25427\,
            I => buf_adcdata_vdc_9
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__25424\,
            I => buf_adcdata_vdc_9
        );

    \I__3600\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25415\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25412\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__25415\,
            I => \N__25409\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__25412\,
            I => cmd_rdadcbuf_17
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__25409\,
            I => cmd_rdadcbuf_17
        );

    \I__3595\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__25398\,
            I => \N__25394\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__25397\,
            I => \N__25391\
        );

    \I__3591\ : Span4Mux_v
    port map (
            O => \N__25394\,
            I => \N__25388\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25385\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__25388\,
            I => buf_adcdata_vdc_6
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__25385\,
            I => buf_adcdata_vdc_6
        );

    \I__3587\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25376\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25373\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__25376\,
            I => cmd_rdadcbuf_11
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25373\,
            I => cmd_rdadcbuf_11
        );

    \I__3583\ : InMux
    port map (
            O => \N__25368\,
            I => \N__25365\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__25365\,
            I => \N__25360\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25357\
        );

    \I__3580\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25354\
        );

    \I__3579\ : Span4Mux_v
    port map (
            O => \N__25360\,
            I => \N__25351\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__25357\,
            I => buf_dds1_5
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__25354\,
            I => buf_dds1_5
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__25351\,
            I => buf_dds1_5
        );

    \I__3575\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25340\
        );

    \I__3574\ : InMux
    port map (
            O => \N__25343\,
            I => \N__25337\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25340\,
            I => cmd_rdadcbuf_21
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25337\,
            I => cmd_rdadcbuf_21
        );

    \I__3571\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25329\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__25329\,
            I => \N__25325\
        );

    \I__3569\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25322\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__25325\,
            I => cmd_rdadcbuf_33
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25322\,
            I => cmd_rdadcbuf_33
        );

    \I__3566\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25310\
        );

    \I__3565\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25310\
        );

    \I__3564\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25307\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__25310\,
            I => cmd_rdadctmp_4_adj_1519
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__25307\,
            I => cmd_rdadctmp_4_adj_1519
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__25302\,
            I => \N__25297\
        );

    \I__3560\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25294\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25291\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25288\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__25294\,
            I => cmd_rdadctmp_5_adj_1518
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__25291\,
            I => cmd_rdadctmp_5_adj_1518
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__25288\,
            I => cmd_rdadctmp_5_adj_1518
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__25281\,
            I => \N__25278\
        );

    \I__3553\ : InMux
    port map (
            O => \N__25278\,
            I => \N__25273\
        );

    \I__3552\ : InMux
    port map (
            O => \N__25277\,
            I => \N__25270\
        );

    \I__3551\ : InMux
    port map (
            O => \N__25276\,
            I => \N__25267\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__25273\,
            I => cmd_rdadctmp_7_adj_1516
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__25270\,
            I => cmd_rdadctmp_7_adj_1516
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__25267\,
            I => cmd_rdadctmp_7_adj_1516
        );

    \I__3547\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25255\
        );

    \I__3546\ : InMux
    port map (
            O => \N__25259\,
            I => \N__25252\
        );

    \I__3545\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25249\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__25255\,
            I => \N__25246\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__25252\,
            I => cmd_rdadctmp_19_adj_1504
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__25249\,
            I => cmd_rdadctmp_19_adj_1504
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__25246\,
            I => cmd_rdadctmp_19_adj_1504
        );

    \I__3540\ : CascadeMux
    port map (
            O => \N__25239\,
            I => \N__25235\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__25238\,
            I => \N__25231\
        );

    \I__3538\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25228\
        );

    \I__3537\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25225\
        );

    \I__3536\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25222\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__25228\,
            I => cmd_rdadctmp_8_adj_1515
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__25225\,
            I => cmd_rdadctmp_8_adj_1515
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__25222\,
            I => cmd_rdadctmp_8_adj_1515
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__25215\,
            I => \N__25210\
        );

    \I__3531\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25207\
        );

    \I__3530\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25204\
        );

    \I__3529\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25201\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__25207\,
            I => cmd_rdadctmp_9_adj_1514
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__25204\,
            I => cmd_rdadctmp_9_adj_1514
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__25201\,
            I => cmd_rdadctmp_9_adj_1514
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__25194\,
            I => \N__25190\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__25193\,
            I => \N__25186\
        );

    \I__3523\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25183\
        );

    \I__3522\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25180\
        );

    \I__3521\ : InMux
    port map (
            O => \N__25186\,
            I => \N__25177\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__25183\,
            I => \N__25174\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__25180\,
            I => cmd_rdadctmp_10_adj_1513
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__25177\,
            I => cmd_rdadctmp_10_adj_1513
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__25174\,
            I => cmd_rdadctmp_10_adj_1513
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__25167\,
            I => \N__25162\
        );

    \I__3515\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25157\
        );

    \I__3514\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25157\
        );

    \I__3513\ : InMux
    port map (
            O => \N__25162\,
            I => \N__25154\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__25157\,
            I => cmd_rdadctmp_11_adj_1512
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__25154\,
            I => cmd_rdadctmp_11_adj_1512
        );

    \I__3510\ : InMux
    port map (
            O => \N__25149\,
            I => \N__25142\
        );

    \I__3509\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25142\
        );

    \I__3508\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25139\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__25142\,
            I => cmd_rdadctmp_12_adj_1511
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__25139\,
            I => cmd_rdadctmp_12_adj_1511
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__25134\,
            I => \N__25130\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__25133\,
            I => \N__25127\
        );

    \I__3503\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25121\
        );

    \I__3502\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25121\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__25126\,
            I => \N__25118\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__25121\,
            I => \N__25115\
        );

    \I__3499\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25112\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__25115\,
            I => cmd_rdadctmp_13_adj_1510
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__25112\,
            I => cmd_rdadctmp_13_adj_1510
        );

    \I__3496\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25104\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__25104\,
            I => \N__25101\
        );

    \I__3494\ : Span4Mux_v
    port map (
            O => \N__25101\,
            I => \N__25097\
        );

    \I__3493\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25094\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__25097\,
            I => cmd_rdadcbuf_27
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__25094\,
            I => cmd_rdadcbuf_27
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__25089\,
            I => \ADC_VDC.n10309_cascade_\
        );

    \I__3489\ : CEMux
    port map (
            O => \N__25086\,
            I => \N__25083\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__25083\,
            I => \N__25080\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__25080\,
            I => \N__25077\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__25077\,
            I => \ADC_VDC.n13276\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__25074\,
            I => \N__25069\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__25073\,
            I => \N__25066\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__25072\,
            I => \N__25063\
        );

    \I__3482\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25060\
        );

    \I__3481\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25057\
        );

    \I__3480\ : InMux
    port map (
            O => \N__25063\,
            I => \N__25054\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__25060\,
            I => cmd_rdadctmp_1_adj_1522
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__25057\,
            I => cmd_rdadctmp_1_adj_1522
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__25054\,
            I => cmd_rdadctmp_1_adj_1522
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__25047\,
            I => \N__25042\
        );

    \I__3475\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25037\
        );

    \I__3474\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25037\
        );

    \I__3473\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25034\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__25037\,
            I => cmd_rdadctmp_2_adj_1521
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__25034\,
            I => cmd_rdadctmp_2_adj_1521
        );

    \I__3470\ : CascadeMux
    port map (
            O => \N__25029\,
            I => \N__25024\
        );

    \I__3469\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25019\
        );

    \I__3468\ : InMux
    port map (
            O => \N__25027\,
            I => \N__25019\
        );

    \I__3467\ : InMux
    port map (
            O => \N__25024\,
            I => \N__25016\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__25019\,
            I => cmd_rdadctmp_3_adj_1520
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__25016\,
            I => cmd_rdadctmp_3_adj_1520
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__25011\,
            I => \ADC_IAC.n21159_cascade_\
        );

    \I__3463\ : CEMux
    port map (
            O => \N__25008\,
            I => \N__25005\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__25002\
        );

    \I__3461\ : Odrv12
    port map (
            O => \N__25002\,
            I => \ADC_IAC.n21160\
        );

    \I__3460\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24993\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24993\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24993\,
            I => cmd_rdadctmp_1
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__24990\,
            I => \N__24986\
        );

    \I__3456\ : InMux
    port map (
            O => \N__24989\,
            I => \N__24983\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24980\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24983\,
            I => cmd_rdadctmp_2
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__24980\,
            I => cmd_rdadctmp_2
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__24975\,
            I => \N__24972\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24969\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__3449\ : Span4Mux_v
    port map (
            O => \N__24966\,
            I => \N__24963\
        );

    \I__3448\ : Sp12to4
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__3447\ : Span12Mux_h
    port map (
            O => \N__24960\,
            I => \N__24957\
        );

    \I__3446\ : Odrv12
    port map (
            O => \N__24957\,
            I => \IAC_MISO\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__24954\,
            I => \N__24951\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24951\,
            I => \N__24945\
        );

    \I__3443\ : InMux
    port map (
            O => \N__24950\,
            I => \N__24945\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__24945\,
            I => cmd_rdadctmp_0
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__24942\,
            I => \N__24936\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24941\,
            I => \N__24932\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__24940\,
            I => \N__24929\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24919\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24919\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24919\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__24932\,
            I => \N__24915\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24912\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__24928\,
            I => \N__24909\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__24927\,
            I => \N__24905\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24926\,
            I => \N__24900\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24897\
        );

    \I__3429\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24894\
        );

    \I__3428\ : Span4Mux_v
    port map (
            O => \N__24915\,
            I => \N__24891\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__24912\,
            I => \N__24888\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24885\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24908\,
            I => \N__24878\
        );

    \I__3424\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24878\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24878\
        );

    \I__3422\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24875\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__24900\,
            I => \N__24868\
        );

    \I__3420\ : Span4Mux_v
    port map (
            O => \N__24897\,
            I => \N__24868\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__24894\,
            I => \N__24868\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__24891\,
            I => \DTRIG_N_958\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__24888\,
            I => \DTRIG_N_958\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__24885\,
            I => \DTRIG_N_958\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__24878\,
            I => \DTRIG_N_958\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24875\,
            I => \DTRIG_N_958\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__24868\,
            I => \DTRIG_N_958\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24847\
        );

    \I__3411\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24843\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24853\,
            I => \N__24834\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24834\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24851\,
            I => \N__24829\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24850\,
            I => \N__24829\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24847\,
            I => \N__24825\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24822\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__24843\,
            I => \N__24819\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24816\
        );

    \I__3402\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24809\
        );

    \I__3401\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24809\
        );

    \I__3400\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24809\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24804\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24804\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24801\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__24825\,
            I => adc_state_1
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__24822\,
            I => adc_state_1
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__24819\,
            I => adc_state_1
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__24816\,
            I => adc_state_1
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__24809\,
            I => adc_state_1
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__24804\,
            I => adc_state_1
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__24801\,
            I => adc_state_1
        );

    \I__3389\ : IoInMux
    port map (
            O => \N__24786\,
            I => \N__24783\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__24783\,
            I => \N__24780\
        );

    \I__3387\ : IoSpan4Mux
    port map (
            O => \N__24780\,
            I => \N__24777\
        );

    \I__3386\ : Span4Mux_s3_v
    port map (
            O => \N__24777\,
            I => \N__24773\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__24776\,
            I => \N__24770\
        );

    \I__3384\ : Span4Mux_v
    port map (
            O => \N__24773\,
            I => \N__24767\
        );

    \I__3383\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24764\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__24767\,
            I => \IAC_SCLK\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24764\,
            I => \IAC_SCLK\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24756\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24753\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__24753\,
            I => \N__24750\
        );

    \I__3377\ : Span4Mux_v
    port map (
            O => \N__24750\,
            I => \N__24746\
        );

    \I__3376\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24743\
        );

    \I__3375\ : Span4Mux_v
    port map (
            O => \N__24746\,
            I => \N__24739\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__24743\,
            I => \N__24736\
        );

    \I__3373\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24733\
        );

    \I__3372\ : Sp12to4
    port map (
            O => \N__24739\,
            I => \N__24730\
        );

    \I__3371\ : Span4Mux_h
    port map (
            O => \N__24736\,
            I => \N__24727\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__24733\,
            I => buf_adcdata_iac_17
        );

    \I__3369\ : Odrv12
    port map (
            O => \N__24730\,
            I => buf_adcdata_iac_17
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__24727\,
            I => buf_adcdata_iac_17
        );

    \I__3367\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24717\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__24717\,
            I => \N__24714\
        );

    \I__3365\ : Span4Mux_v
    port map (
            O => \N__24714\,
            I => \N__24710\
        );

    \I__3364\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24707\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__24710\,
            I => cmd_rdadctmp_4_adj_1488
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__24707\,
            I => cmd_rdadctmp_4_adj_1488
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__3360\ : InMux
    port map (
            O => \N__24699\,
            I => \N__24693\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24693\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24693\,
            I => cmd_rdadctmp_5_adj_1487
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__3356\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__3354\ : Span4Mux_h
    port map (
            O => \N__24681\,
            I => \N__24677\
        );

    \I__3353\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__24677\,
            I => cmd_rdadctmp_6_adj_1486
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__24674\,
            I => cmd_rdadctmp_6_adj_1486
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__3349\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__24663\,
            I => \N__24660\
        );

    \I__3347\ : Span4Mux_v
    port map (
            O => \N__24660\,
            I => \N__24655\
        );

    \I__3346\ : InMux
    port map (
            O => \N__24659\,
            I => \N__24650\
        );

    \I__3345\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24650\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__24655\,
            I => cmd_rdadctmp_22
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__24650\,
            I => cmd_rdadctmp_22
        );

    \I__3342\ : SRMux
    port map (
            O => \N__24645\,
            I => \N__24642\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__24642\,
            I => \N__24638\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__24641\,
            I => \N__24635\
        );

    \I__3339\ : Span4Mux_h
    port map (
            O => \N__24638\,
            I => \N__24632\
        );

    \I__3338\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24629\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__24632\,
            I => n15092
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__24629\,
            I => n15092
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__24624\,
            I => \N__24620\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__24623\,
            I => \N__24617\
        );

    \I__3333\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24612\
        );

    \I__3332\ : InMux
    port map (
            O => \N__24617\,
            I => \N__24607\
        );

    \I__3331\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24607\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__24615\,
            I => \N__24603\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24612\,
            I => \N__24598\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24607\,
            I => \N__24598\
        );

    \I__3327\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24595\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24603\,
            I => \N__24592\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__24598\,
            I => \N__24587\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__24595\,
            I => \N__24587\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__24592\,
            I => \N__24582\
        );

    \I__3322\ : Sp12to4
    port map (
            O => \N__24587\,
            I => \N__24582\
        );

    \I__3321\ : Span12Mux_h
    port map (
            O => \N__24582\,
            I => \N__24579\
        );

    \I__3320\ : Odrv12
    port map (
            O => \N__24579\,
            I => \IAC_DRDY\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__24576\,
            I => \N__24573\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__24570\,
            I => \CLK_DDS.tmp_buf_3\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__24561\,
            I => \CLK_DDS.tmp_buf_4\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24552\,
            I => \CLK_DDS.tmp_buf_5\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__24549\,
            I => \N__24546\
        );

    \I__3309\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24543\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__24543\,
            I => \CLK_DDS.tmp_buf_6\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24534\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24534\,
            I => \N__24531\
        );

    \I__3304\ : Odrv12
    port map (
            O => \N__24531\,
            I => \CLK_DDS.tmp_buf_7\
        );

    \I__3303\ : InMux
    port map (
            O => \N__24528\,
            I => \N__24525\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__24525\,
            I => \N__24522\
        );

    \I__3301\ : Span12Mux_s8_h
    port map (
            O => \N__24522\,
            I => \N__24517\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24514\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24520\,
            I => \N__24511\
        );

    \I__3298\ : Span12Mux_h
    port map (
            O => \N__24517\,
            I => \N__24508\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24514\,
            I => \N__24505\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__24511\,
            I => buf_adcdata_vac_17
        );

    \I__3295\ : Odrv12
    port map (
            O => \N__24508\,
            I => buf_adcdata_vac_17
        );

    \I__3294\ : Odrv12
    port map (
            O => \N__24505\,
            I => buf_adcdata_vac_17
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__24498\,
            I => \N__24494\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24497\,
            I => \N__24487\
        );

    \I__3291\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24487\
        );

    \I__3290\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24484\
        );

    \I__3289\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24481\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__24487\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__24484\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__24481\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__3285\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24467\
        );

    \I__3284\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24467\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__24472\,
            I => \N__24464\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__24467\,
            I => \N__24461\
        );

    \I__3281\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24458\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__24461\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__24458\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__24453\,
            I => \N__24450\
        );

    \I__3277\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24447\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__24447\,
            I => \N__24444\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__24444\,
            I => \SIG_DDS.n10\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24430\
        );

    \I__3273\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24430\
        );

    \I__3272\ : InMux
    port map (
            O => \N__24439\,
            I => \N__24430\
        );

    \I__3271\ : InMux
    port map (
            O => \N__24438\,
            I => \N__24427\
        );

    \I__3270\ : InMux
    port map (
            O => \N__24437\,
            I => \N__24424\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__24430\,
            I => bit_cnt_0
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__24427\,
            I => bit_cnt_0
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__24424\,
            I => bit_cnt_0
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__24417\,
            I => \N__24413\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__24416\,
            I => \N__24409\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24406\
        );

    \I__3263\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24401\
        );

    \I__3262\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24401\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__24406\,
            I => cmd_rdadctmp_28_adj_1464
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24401\,
            I => cmd_rdadctmp_28_adj_1464
        );

    \I__3259\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24393\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__24393\,
            I => \N__24389\
        );

    \I__3257\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24386\
        );

    \I__3256\ : Odrv12
    port map (
            O => \N__24389\,
            I => tmp_buf_15_adj_1497
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__24386\,
            I => tmp_buf_15_adj_1497
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__3253\ : InMux
    port map (
            O => \N__24378\,
            I => \N__24375\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__24375\,
            I => \CLK_DDS.tmp_buf_0\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24369\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__24369\,
            I => \CLK_DDS.tmp_buf_1\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__24366\,
            I => \N__24363\
        );

    \I__3248\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24360\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__24360\,
            I => \CLK_DDS.tmp_buf_2\
        );

    \I__3246\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24354\,
            I => \N__24350\
        );

    \I__3244\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24347\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__24350\,
            I => \N__24343\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24340\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24337\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__24343\,
            I => cmd_rdadctmp_13
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__24340\,
            I => cmd_rdadctmp_13
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__24337\,
            I => cmd_rdadctmp_13
        );

    \I__3237\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24327\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__24327\,
            I => \N__24323\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__24326\,
            I => \N__24320\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__24323\,
            I => \N__24317\
        );

    \I__3233\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24314\
        );

    \I__3232\ : Sp12to4
    port map (
            O => \N__24317\,
            I => \N__24308\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24308\
        );

    \I__3230\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24305\
        );

    \I__3229\ : Odrv12
    port map (
            O => \N__24308\,
            I => cmd_rdadctmp_10
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__24305\,
            I => cmd_rdadctmp_10
        );

    \I__3227\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__24294\,
            I => \N__24291\
        );

    \I__3224\ : Span4Mux_h
    port map (
            O => \N__24291\,
            I => \N__24287\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__24290\,
            I => \N__24284\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__24287\,
            I => \N__24280\
        );

    \I__3221\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24277\
        );

    \I__3220\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24274\
        );

    \I__3219\ : Span4Mux_h
    port map (
            O => \N__24280\,
            I => \N__24271\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__24277\,
            I => buf_adcdata_iac_2
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__24274\,
            I => buf_adcdata_iac_2
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__24271\,
            I => buf_adcdata_iac_2
        );

    \I__3215\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24261\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__24261\,
            I => \N__24258\
        );

    \I__3213\ : Span4Mux_h
    port map (
            O => \N__24258\,
            I => \N__24254\
        );

    \I__3212\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24250\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__24254\,
            I => \N__24247\
        );

    \I__3210\ : InMux
    port map (
            O => \N__24253\,
            I => \N__24244\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__24250\,
            I => buf_adcdata_vac_5
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__24247\,
            I => buf_adcdata_vac_5
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__24244\,
            I => buf_adcdata_vac_5
        );

    \I__3206\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24234\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__24234\,
            I => \N__24231\
        );

    \I__3204\ : Span4Mux_h
    port map (
            O => \N__24231\,
            I => \N__24228\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__24228\,
            I => \N__24223\
        );

    \I__3202\ : InMux
    port map (
            O => \N__24227\,
            I => \N__24218\
        );

    \I__3201\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24218\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__24223\,
            I => buf_adcdata_iac_5
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__24218\,
            I => buf_adcdata_iac_5
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__24213\,
            I => \n19_adj_1603_cascade_\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__24210\,
            I => \n22377_cascade_\
        );

    \I__3196\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24204\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__24204\,
            I => n21237
        );

    \I__3194\ : InMux
    port map (
            O => \N__24201\,
            I => \ADC_VDC.n19869\
        );

    \I__3193\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24195\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__24195\,
            I => \N__24192\
        );

    \I__3191\ : Span4Mux_v
    port map (
            O => \N__24192\,
            I => \N__24188\
        );

    \I__3190\ : InMux
    port map (
            O => \N__24191\,
            I => \N__24185\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__24188\,
            I => cmd_rdadcbuf_29
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__24185\,
            I => cmd_rdadcbuf_29
        );

    \I__3187\ : InMux
    port map (
            O => \N__24180\,
            I => \ADC_VDC.n19870\
        );

    \I__3186\ : InMux
    port map (
            O => \N__24177\,
            I => \ADC_VDC.n19871\
        );

    \I__3185\ : InMux
    port map (
            O => \N__24174\,
            I => \ADC_VDC.n19872\
        );

    \I__3184\ : InMux
    port map (
            O => \N__24171\,
            I => \bfn_8_10_0_\
        );

    \I__3183\ : InMux
    port map (
            O => \N__24168\,
            I => \ADC_VDC.n19874\
        );

    \I__3182\ : InMux
    port map (
            O => \N__24165\,
            I => \ADC_VDC.n19875\
        );

    \I__3181\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24159\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24156\
        );

    \I__3179\ : Sp12to4
    port map (
            O => \N__24156\,
            I => \N__24152\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__24155\,
            I => \N__24149\
        );

    \I__3177\ : Span12Mux_v
    port map (
            O => \N__24152\,
            I => \N__24146\
        );

    \I__3176\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24143\
        );

    \I__3175\ : Odrv12
    port map (
            O => \N__24146\,
            I => buf_adcdata_vdc_18
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__24143\,
            I => buf_adcdata_vdc_18
        );

    \I__3173\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24135\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__3171\ : Sp12to4
    port map (
            O => \N__24132\,
            I => \N__24127\
        );

    \I__3170\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24124\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__24130\,
            I => \N__24121\
        );

    \I__3168\ : Span12Mux_v
    port map (
            O => \N__24127\,
            I => \N__24118\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__24124\,
            I => \N__24115\
        );

    \I__3166\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24112\
        );

    \I__3165\ : Span12Mux_h
    port map (
            O => \N__24118\,
            I => \N__24109\
        );

    \I__3164\ : Span4Mux_h
    port map (
            O => \N__24115\,
            I => \N__24106\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__24112\,
            I => buf_adcdata_vac_18
        );

    \I__3162\ : Odrv12
    port map (
            O => \N__24109\,
            I => buf_adcdata_vac_18
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__24106\,
            I => buf_adcdata_vac_18
        );

    \I__3160\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24096\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__24096\,
            I => n19_adj_1692
        );

    \I__3158\ : InMux
    port map (
            O => \N__24093\,
            I => \ADC_VDC.n19860\
        );

    \I__3157\ : InMux
    port map (
            O => \N__24090\,
            I => \ADC_VDC.n19861\
        );

    \I__3156\ : InMux
    port map (
            O => \N__24087\,
            I => \ADC_VDC.n19862\
        );

    \I__3155\ : InMux
    port map (
            O => \N__24084\,
            I => \ADC_VDC.n19863\
        );

    \I__3154\ : InMux
    port map (
            O => \N__24081\,
            I => \ADC_VDC.n19864\
        );

    \I__3153\ : InMux
    port map (
            O => \N__24078\,
            I => \bfn_8_9_0_\
        );

    \I__3152\ : InMux
    port map (
            O => \N__24075\,
            I => \ADC_VDC.n19866\
        );

    \I__3151\ : InMux
    port map (
            O => \N__24072\,
            I => \ADC_VDC.n19867\
        );

    \I__3150\ : InMux
    port map (
            O => \N__24069\,
            I => \ADC_VDC.n19868\
        );

    \I__3149\ : InMux
    port map (
            O => \N__24066\,
            I => \ADC_VDC.n19852\
        );

    \I__3148\ : InMux
    port map (
            O => \N__24063\,
            I => \ADC_VDC.n19853\
        );

    \I__3147\ : InMux
    port map (
            O => \N__24060\,
            I => \ADC_VDC.n19854\
        );

    \I__3146\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24054\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24051\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__24051\,
            I => \N__24047\
        );

    \I__3143\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24044\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__24047\,
            I => cmd_rdadcbuf_14
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__24044\,
            I => cmd_rdadcbuf_14
        );

    \I__3140\ : InMux
    port map (
            O => \N__24039\,
            I => \ADC_VDC.n19855\
        );

    \I__3139\ : InMux
    port map (
            O => \N__24036\,
            I => \ADC_VDC.n19856\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__24033\,
            I => \N__24030\
        );

    \I__3137\ : InMux
    port map (
            O => \N__24030\,
            I => \N__24025\
        );

    \I__3136\ : InMux
    port map (
            O => \N__24029\,
            I => \N__24020\
        );

    \I__3135\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24020\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__24025\,
            I => \N__24017\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__24020\,
            I => cmd_rdadctmp_16_adj_1507
        );

    \I__3132\ : Odrv12
    port map (
            O => \N__24017\,
            I => cmd_rdadctmp_16_adj_1507
        );

    \I__3131\ : InMux
    port map (
            O => \N__24012\,
            I => \bfn_8_8_0_\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__24009\,
            I => \N__24006\
        );

    \I__3129\ : InMux
    port map (
            O => \N__24006\,
            I => \N__24001\
        );

    \I__3128\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23996\
        );

    \I__3127\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23996\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__24001\,
            I => \N__23993\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23996\,
            I => cmd_rdadctmp_17_adj_1506
        );

    \I__3124\ : Odrv12
    port map (
            O => \N__23993\,
            I => cmd_rdadctmp_17_adj_1506
        );

    \I__3123\ : InMux
    port map (
            O => \N__23988\,
            I => \ADC_VDC.n19858\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__23985\,
            I => \N__23982\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23978\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__23981\,
            I => \N__23975\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23971\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23968\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23965\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__23971\,
            I => \N__23962\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__23968\,
            I => cmd_rdadctmp_18_adj_1505
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23965\,
            I => cmd_rdadctmp_18_adj_1505
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__23962\,
            I => cmd_rdadctmp_18_adj_1505
        );

    \I__3112\ : InMux
    port map (
            O => \N__23955\,
            I => \ADC_VDC.n19859\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23952\,
            I => \N__23949\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23949\,
            I => \ADC_VDC.cmd_rdadcbuf_2\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23946\,
            I => \ADC_VDC.n19843\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23940\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23940\,
            I => \ADC_VDC.cmd_rdadcbuf_3\
        );

    \I__3106\ : InMux
    port map (
            O => \N__23937\,
            I => \ADC_VDC.n19844\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__23934\,
            I => \N__23931\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23931\,
            I => \N__23928\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__23925\,
            I => \ADC_VDC.cmd_rdadcbuf_4\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23922\,
            I => \ADC_VDC.n19845\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23916\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23916\,
            I => \ADC_VDC.cmd_rdadcbuf_5\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23913\,
            I => \ADC_VDC.n19846\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__23910\,
            I => \N__23906\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__23909\,
            I => \N__23903\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23899\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23896\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23902\,
            I => \N__23893\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__23899\,
            I => \N__23890\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23896\,
            I => cmd_rdadctmp_6_adj_1517
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23893\,
            I => cmd_rdadctmp_6_adj_1517
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__23890\,
            I => cmd_rdadctmp_6_adj_1517
        );

    \I__3088\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23880\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__23880\,
            I => \ADC_VDC.cmd_rdadcbuf_6\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23877\,
            I => \ADC_VDC.n19847\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__23874\,
            I => \N__23871\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__23868\,
            I => \ADC_VDC.cmd_rdadcbuf_7\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23865\,
            I => \ADC_VDC.n19848\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23859\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__23859\,
            I => \ADC_VDC.cmd_rdadcbuf_8\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23856\,
            I => \bfn_8_7_0_\
        );

    \I__3078\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23850\,
            I => \ADC_VDC.cmd_rdadcbuf_9\
        );

    \I__3076\ : InMux
    port map (
            O => \N__23847\,
            I => \ADC_VDC.n19850\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23841\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__23841\,
            I => \ADC_VDC.cmd_rdadcbuf_10\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23838\,
            I => \ADC_VDC.n19851\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__23835\,
            I => \N__23832\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23827\
        );

    \I__3070\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23822\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23830\,
            I => \N__23822\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23819\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__23822\,
            I => cmd_rdadctmp_0_adj_1523
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__23819\,
            I => cmd_rdadctmp_0_adj_1523
        );

    \I__3065\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23811\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__23811\,
            I => \ADC_VDC.cmd_rdadcbuf_0\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23805\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__23805\,
            I => \ADC_VDC.cmd_rdadcbuf_1\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23802\,
            I => \ADC_VDC.n19842\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23796\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__23796\,
            I => n21082
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__23793\,
            I => \n21082_cascade_\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23784\
        );

    \I__3056\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23784\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23784\,
            I => cmd_rdadctmp_3
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__23781\,
            I => \n12771_cascade_\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__23778\,
            I => \N__23775\
        );

    \I__3052\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23769\
        );

    \I__3051\ : InMux
    port map (
            O => \N__23774\,
            I => \N__23769\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__23769\,
            I => cmd_rdadctmp_4
        );

    \I__3049\ : InMux
    port map (
            O => \N__23766\,
            I => \N__23760\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23760\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__23760\,
            I => cmd_rdadctmp_5
        );

    \I__3046\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23754\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23754\,
            I => \ADC_IAC.n17\
        );

    \I__3044\ : IoInMux
    port map (
            O => \N__23751\,
            I => \N__23748\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__23748\,
            I => \N__23745\
        );

    \I__3042\ : Span4Mux_s2_v
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__3041\ : Span4Mux_v
    port map (
            O => \N__23742\,
            I => \N__23739\
        );

    \I__3040\ : Span4Mux_h
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__23736\,
            I => \DDS_MCLK1\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__23727\,
            I => \N__23724\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__23724\,
            I => \N__23720\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__23723\,
            I => \N__23717\
        );

    \I__3033\ : Span4Mux_h
    port map (
            O => \N__23720\,
            I => \N__23714\
        );

    \I__3032\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23711\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__23714\,
            I => \buf_readRTD_7\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__23711\,
            I => \buf_readRTD_7\
        );

    \I__3029\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23703\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__23703\,
            I => \N__23700\
        );

    \I__3027\ : Odrv12
    port map (
            O => \N__23700\,
            I => n16_adj_1690
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__23697\,
            I => \N__23694\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23691\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__23685\,
            I => n17_adj_1691
        );

    \I__3021\ : CEMux
    port map (
            O => \N__23682\,
            I => \N__23679\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__23676\,
            I => \ADC_IAC.n12\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__23670\,
            I => \ADC_IAC.n21457\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__23667\,
            I => \N__23664\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__23661\,
            I => \N__23658\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__23658\,
            I => \N__23654\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23657\,
            I => \N__23651\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__23654\,
            I => cmd_rdadctmp_7
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__23651\,
            I => cmd_rdadctmp_7
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__3008\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23637\
        );

    \I__3007\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23637\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__23637\,
            I => cmd_rdadctmp_6
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__23634\,
            I => \N__23631\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23628\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__23628\,
            I => \CLK_DDS.tmp_buf_10\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23619\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23619\,
            I => \CLK_DDS.tmp_buf_11\
        );

    \I__2999\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__23610\,
            I => \CLK_DDS.tmp_buf_12\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__23607\,
            I => \N__23604\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__23601\,
            I => \N__23598\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__23598\,
            I => \CLK_DDS.tmp_buf_13\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__23595\,
            I => \N__23592\
        );

    \I__2991\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23589\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23589\,
            I => \CLK_DDS.tmp_buf_14\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__23586\,
            I => \N__23583\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23580\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23580\,
            I => \CLK_DDS.tmp_buf_9\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__23577\,
            I => \N__23574\
        );

    \I__2985\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23571\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__23571\,
            I => \CLK_DDS.tmp_buf_8\
        );

    \I__2983\ : InMux
    port map (
            O => \N__23568\,
            I => \N__23565\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__23565\,
            I => \N__23562\
        );

    \I__2981\ : Span12Mux_v
    port map (
            O => \N__23562\,
            I => \N__23557\
        );

    \I__2980\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23554\
        );

    \I__2979\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23551\
        );

    \I__2978\ : Span12Mux_h
    port map (
            O => \N__23557\,
            I => \N__23548\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__23554\,
            I => \N__23545\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__23551\,
            I => buf_adcdata_vac_9
        );

    \I__2975\ : Odrv12
    port map (
            O => \N__23548\,
            I => buf_adcdata_vac_9
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__23545\,
            I => buf_adcdata_vac_9
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__23538\,
            I => \N__23535\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23531\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__23534\,
            I => \N__23528\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23524\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23519\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23519\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__23524\,
            I => cmd_rdadctmp_11
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__23519\,
            I => cmd_rdadctmp_11
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__23514\,
            I => \N__23510\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23504\
        );

    \I__2963\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23504\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23501\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__23504\,
            I => cmd_rdadctmp_12
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__23501\,
            I => cmd_rdadctmp_12
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__23496\,
            I => \N__23493\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23490\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23486\
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__23489\,
            I => \N__23483\
        );

    \I__2955\ : Span4Mux_h
    port map (
            O => \N__23486\,
            I => \N__23479\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23476\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23473\
        );

    \I__2952\ : Odrv4
    port map (
            O => \N__23479\,
            I => cmd_rdadctmp_8
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__23476\,
            I => cmd_rdadctmp_8
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__23473\,
            I => cmd_rdadctmp_8
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__23466\,
            I => \N__23462\
        );

    \I__2948\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23458\
        );

    \I__2947\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23453\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23453\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23458\,
            I => cmd_rdadctmp_17_adj_1475
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__23453\,
            I => cmd_rdadctmp_17_adj_1475
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__23448\,
            I => \N__23444\
        );

    \I__2942\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23438\
        );

    \I__2941\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23438\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__23443\,
            I => \N__23435\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__23438\,
            I => \N__23432\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23429\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__23432\,
            I => cmd_rdadctmp_29_adj_1463
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__23429\,
            I => cmd_rdadctmp_29_adj_1463
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__23424\,
            I => \N__23420\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__23423\,
            I => \N__23417\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23413\
        );

    \I__2932\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23408\
        );

    \I__2931\ : InMux
    port map (
            O => \N__23416\,
            I => \N__23408\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__23413\,
            I => cmd_rdadctmp_9_adj_1483
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23408\,
            I => cmd_rdadctmp_9_adj_1483
        );

    \I__2928\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23400\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__23400\,
            I => \N__23397\
        );

    \I__2926\ : Span4Mux_v
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__23391\,
            I => buf_data_iac_6
        );

    \I__2923\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23385\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__23382\,
            I => n22_adj_1601
        );

    \I__2920\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__2918\ : Span4Mux_v
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__2916\ : Sp12to4
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__2915\ : Span12Mux_h
    port map (
            O => \N__23364\,
            I => \N__23361\
        );

    \I__2914\ : Odrv12
    port map (
            O => \N__23361\,
            I => buf_data_iac_2
        );

    \I__2913\ : InMux
    port map (
            O => \N__23358\,
            I => \N__23355\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__23355\,
            I => n22_adj_1613
        );

    \I__2911\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23349\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23345\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23342\
        );

    \I__2908\ : Span4Mux_h
    port map (
            O => \N__23345\,
            I => \N__23337\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__23342\,
            I => \N__23337\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__23337\,
            I => \buf_readRTD_10\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__23334\,
            I => \N__23331\
        );

    \I__2904\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23327\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__23330\,
            I => \N__23324\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23320\
        );

    \I__2901\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23315\
        );

    \I__2900\ : InMux
    port map (
            O => \N__23323\,
            I => \N__23315\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__23320\,
            I => \N__23308\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23308\
        );

    \I__2897\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23303\
        );

    \I__2896\ : InMux
    port map (
            O => \N__23313\,
            I => \N__23303\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__23308\,
            I => \buf_cfgRTD_2\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__23303\,
            I => \buf_cfgRTD_2\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__23298\,
            I => \N__23294\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__23297\,
            I => \N__23291\
        );

    \I__2891\ : InMux
    port map (
            O => \N__23294\,
            I => \N__23288\
        );

    \I__2890\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23285\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__23288\,
            I => \N__23281\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__23285\,
            I => \N__23278\
        );

    \I__2887\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23275\
        );

    \I__2886\ : Odrv12
    port map (
            O => \N__23281\,
            I => cmd_rdadctmp_11_adj_1481
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__23278\,
            I => cmd_rdadctmp_11_adj_1481
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__23275\,
            I => cmd_rdadctmp_11_adj_1481
        );

    \I__2883\ : InMux
    port map (
            O => \N__23268\,
            I => \N__23265\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__2880\ : Sp12to4
    port map (
            O => \N__23259\,
            I => \N__23254\
        );

    \I__2879\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23251\
        );

    \I__2878\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23248\
        );

    \I__2877\ : Span12Mux_h
    port map (
            O => \N__23254\,
            I => \N__23245\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23242\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__23248\,
            I => buf_adcdata_vac_3
        );

    \I__2874\ : Odrv12
    port map (
            O => \N__23245\,
            I => buf_adcdata_vac_3
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__23242\,
            I => buf_adcdata_vac_3
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__23235\,
            I => \N__23232\
        );

    \I__2871\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23229\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__23229\,
            I => \N__23224\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__23228\,
            I => \N__23221\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__23227\,
            I => \N__23218\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__23224\,
            I => \N__23215\
        );

    \I__2866\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23212\
        );

    \I__2865\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23209\
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__23215\,
            I => cmd_rdadctmp_13_adj_1479
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__23212\,
            I => cmd_rdadctmp_13_adj_1479
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__23209\,
            I => cmd_rdadctmp_13_adj_1479
        );

    \I__2861\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23197\
        );

    \I__2860\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23194\
        );

    \I__2859\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23191\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__23197\,
            I => cmd_rdadctmp_30_adj_1462
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__23194\,
            I => cmd_rdadctmp_30_adj_1462
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__23191\,
            I => cmd_rdadctmp_30_adj_1462
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__23184\,
            I => \N__23181\
        );

    \I__2854\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23178\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__23178\,
            I => n20_adj_1693
        );

    \I__2852\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23172\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__23172\,
            I => n22407
        );

    \I__2850\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23166\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__23163\
        );

    \I__2848\ : Span12Mux_s9_h
    port map (
            O => \N__23163\,
            I => \N__23160\
        );

    \I__2847\ : Span12Mux_h
    port map (
            O => \N__23160\,
            I => \N__23155\
        );

    \I__2846\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23150\
        );

    \I__2845\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23150\
        );

    \I__2844\ : Odrv12
    port map (
            O => \N__23155\,
            I => buf_adcdata_vac_2
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__23150\,
            I => buf_adcdata_vac_2
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__23145\,
            I => \n19_adj_1612_cascade_\
        );

    \I__2841\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23139\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__23139\,
            I => \N__23134\
        );

    \I__2839\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23131\
        );

    \I__2838\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23128\
        );

    \I__2837\ : Span4Mux_h
    port map (
            O => \N__23134\,
            I => \N__23125\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__23131\,
            I => \N__23122\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23117\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__23125\,
            I => \N__23117\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__23122\,
            I => \N__23114\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__23117\,
            I => buf_adcdata_vac_6
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__23114\,
            I => buf_adcdata_vac_6
        );

    \I__2830\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23106\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__23106\,
            I => \N__23103\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__23103\,
            I => \N__23100\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__23100\,
            I => \N__23096\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__23099\,
            I => \N__23093\
        );

    \I__2825\ : Sp12to4
    port map (
            O => \N__23096\,
            I => \N__23089\
        );

    \I__2824\ : InMux
    port map (
            O => \N__23093\,
            I => \N__23086\
        );

    \I__2823\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23083\
        );

    \I__2822\ : Span12Mux_h
    port map (
            O => \N__23089\,
            I => \N__23080\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__23086\,
            I => buf_adcdata_vac_22
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__23083\,
            I => buf_adcdata_vac_22
        );

    \I__2819\ : Odrv12
    port map (
            O => \N__23080\,
            I => buf_adcdata_vac_22
        );

    \I__2818\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23070\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__23070\,
            I => \N__23067\
        );

    \I__2816\ : Odrv4
    port map (
            O => \N__23067\,
            I => n22629
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__23064\,
            I => \N__23061\
        );

    \I__2814\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23057\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__23060\,
            I => \N__23054\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__23057\,
            I => \N__23050\
        );

    \I__2811\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23047\
        );

    \I__2810\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23044\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__23050\,
            I => cmd_rdadctmp_14_adj_1478
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__23047\,
            I => cmd_rdadctmp_14_adj_1478
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__23044\,
            I => cmd_rdadctmp_14_adj_1478
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__23037\,
            I => \N__23034\
        );

    \I__2805\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__23027\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__23030\,
            I => \N__23024\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__23027\,
            I => \N__23020\
        );

    \I__2801\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23015\
        );

    \I__2800\ : InMux
    port map (
            O => \N__23023\,
            I => \N__23015\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__23020\,
            I => cmd_rdadctmp_15_adj_1477
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__23015\,
            I => cmd_rdadctmp_15_adj_1477
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__23010\,
            I => \N__23002\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__23009\,
            I => \N__22999\
        );

    \I__2795\ : InMux
    port map (
            O => \N__23008\,
            I => \N__22995\
        );

    \I__2794\ : InMux
    port map (
            O => \N__23007\,
            I => \N__22992\
        );

    \I__2793\ : InMux
    port map (
            O => \N__23006\,
            I => \N__22989\
        );

    \I__2792\ : InMux
    port map (
            O => \N__23005\,
            I => \N__22980\
        );

    \I__2791\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22980\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22980\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22980\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__22995\,
            I => \RTD.n13090\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22992\,
            I => \RTD.n13090\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22989\,
            I => \RTD.n13090\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__22980\,
            I => \RTD.n13090\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__22971\,
            I => \N__22964\
        );

    \I__2783\ : CascadeMux
    port map (
            O => \N__22970\,
            I => \N__22961\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__22969\,
            I => \N__22957\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__22968\,
            I => \N__22954\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__22967\,
            I => \N__22951\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22945\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22942\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22939\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22936\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22954\,
            I => \N__22925\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22925\
        );

    \I__2773\ : InMux
    port map (
            O => \N__22950\,
            I => \N__22925\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22925\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22925\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__22945\,
            I => \N__22916\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__22942\,
            I => \N__22916\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__22939\,
            I => \N__22916\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22936\,
            I => \N__22916\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22913\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__22916\,
            I => \N__22910\
        );

    \I__2764\ : Span4Mux_h
    port map (
            O => \N__22913\,
            I => \N__22907\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__22910\,
            I => \RTD.n21061\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__22907\,
            I => \RTD.n21061\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22902\,
            I => \N__22898\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22895\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__22898\,
            I => \N__22892\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22895\,
            I => \RTD.cfg_buf_0\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__22892\,
            I => \RTD.cfg_buf_0\
        );

    \I__2756\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22883\
        );

    \I__2755\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22880\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__22883\,
            I => \buf_readRTD_9\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__22880\,
            I => \buf_readRTD_9\
        );

    \I__2752\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22871\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__22874\,
            I => \N__22868\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22865\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__2748\ : Odrv12
    port map (
            O => \N__22865\,
            I => buf_adcdata_vdc_3
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__22862\,
            I => buf_adcdata_vdc_3
        );

    \I__2746\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22854\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22854\,
            I => \N__22850\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22847\
        );

    \I__2743\ : Span12Mux_v
    port map (
            O => \N__22850\,
            I => \N__22843\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__22847\,
            I => \N__22840\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22837\
        );

    \I__2740\ : Span12Mux_h
    port map (
            O => \N__22843\,
            I => \N__22834\
        );

    \I__2739\ : Span4Mux_h
    port map (
            O => \N__22840\,
            I => \N__22831\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22837\,
            I => buf_adcdata_iac_3
        );

    \I__2737\ : Odrv12
    port map (
            O => \N__22834\,
            I => buf_adcdata_iac_3
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__22831\,
            I => buf_adcdata_iac_3
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__22824\,
            I => \n19_adj_1609_cascade_\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__22821\,
            I => \N__22818\
        );

    \I__2733\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22811\
        );

    \I__2731\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22808\
        );

    \I__2730\ : Odrv12
    port map (
            O => \N__22811\,
            I => \buf_readRTD_14\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22808\,
            I => \buf_readRTD_14\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__22803\,
            I => \N__22800\
        );

    \I__2727\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22796\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__22799\,
            I => \N__22793\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22789\
        );

    \I__2724\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22786\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22783\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__22789\,
            I => \N__22780\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__22786\,
            I => cmd_rdadctmp_10_adj_1482
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__22783\,
            I => cmd_rdadctmp_10_adj_1482
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__22780\,
            I => cmd_rdadctmp_10_adj_1482
        );

    \I__2718\ : IoInMux
    port map (
            O => \N__22773\,
            I => \N__22770\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__2716\ : Span12Mux_s5_v
    port map (
            O => \N__22767\,
            I => \N__22763\
        );

    \I__2715\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22760\
        );

    \I__2714\ : Odrv12
    port map (
            O => \N__22763\,
            I => \DDS_MOSI1\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__22760\,
            I => \DDS_MOSI1\
        );

    \I__2712\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22749\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22754\,
            I => \N__22749\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__22749\,
            I => \RTD.cfg_buf_5\
        );

    \I__2709\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22743\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__22743\,
            I => \RTD.n11_adj_1444\
        );

    \I__2707\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22734\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22734\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__22734\,
            I => \RTD.cfg_buf_3\
        );

    \I__2704\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22725\
        );

    \I__2703\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22725\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__22725\,
            I => \RTD.cfg_buf_4\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22722\,
            I => \N__22716\
        );

    \I__2700\ : InMux
    port map (
            O => \N__22721\,
            I => \N__22716\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__22716\,
            I => \RTD.cfg_buf_2\
        );

    \I__2698\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22710\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__22710\,
            I => \RTD.n10\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22703\
        );

    \I__2695\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22700\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__22703\,
            I => \RTD.n11\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22700\,
            I => \RTD.n11\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__22695\,
            I => \N__22688\
        );

    \I__2691\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22680\
        );

    \I__2690\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22674\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__22692\,
            I => \N__22671\
        );

    \I__2688\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22663\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22663\
        );

    \I__2686\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22663\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22660\
        );

    \I__2684\ : InMux
    port map (
            O => \N__22685\,
            I => \N__22653\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22684\,
            I => \N__22653\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22653\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22649\
        );

    \I__2680\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22646\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__22678\,
            I => \N__22641\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__22677\,
            I => \N__22636\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22632\
        );

    \I__2676\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22627\
        );

    \I__2675\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22627\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__22663\,
            I => \N__22620\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__22660\,
            I => \N__22620\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22620\
        );

    \I__2671\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22617\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__22649\,
            I => \N__22614\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__22646\,
            I => \N__22611\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__22645\,
            I => \N__22606\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22600\
        );

    \I__2666\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22597\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22640\,
            I => \N__22594\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22587\
        );

    \I__2663\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22587\
        );

    \I__2662\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22587\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__22632\,
            I => \N__22580\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22580\
        );

    \I__2659\ : Span4Mux_v
    port map (
            O => \N__22620\,
            I => \N__22580\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22573\
        );

    \I__2657\ : Span4Mux_h
    port map (
            O => \N__22614\,
            I => \N__22573\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__22611\,
            I => \N__22573\
        );

    \I__2655\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22560\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22560\
        );

    \I__2653\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22560\
        );

    \I__2652\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22560\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22560\
        );

    \I__2650\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22560\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22600\,
            I => \RTD.adc_state_3\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__22597\,
            I => \RTD.adc_state_3\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22594\,
            I => \RTD.adc_state_3\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__22587\,
            I => \RTD.adc_state_3\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__22580\,
            I => \RTD.adc_state_3\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__22573\,
            I => \RTD.adc_state_3\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__22560\,
            I => \RTD.adc_state_3\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__22545\,
            I => \N__22541\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22538\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22535\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22532\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__22535\,
            I => \RTD.n21036\
        );

    \I__2637\ : Odrv12
    port map (
            O => \N__22532\,
            I => \RTD.n21036\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22523\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22526\,
            I => \N__22520\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22523\,
            I => \N__22517\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22513\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__22517\,
            I => \N__22509\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22506\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__22513\,
            I => \N__22503\
        );

    \I__2629\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22500\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__22509\,
            I => \RTD.n21199\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__22506\,
            I => \RTD.n21199\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__22503\,
            I => \RTD.n21199\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__22500\,
            I => \RTD.n21199\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__22491\,
            I => \RTD.n13090_cascade_\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22484\
        );

    \I__2622\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22481\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__22484\,
            I => \RTD.cfg_buf_1\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__22481\,
            I => \RTD.cfg_buf_1\
        );

    \I__2619\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22473\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__22473\,
            I => \RTD.n12\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22464\
        );

    \I__2616\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22464\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__22464\,
            I => \RTD.cfg_buf_7\
        );

    \I__2614\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__22458\,
            I => \RTD.cfg_tmp_1\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__22455\,
            I => \N__22452\
        );

    \I__2611\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__22449\,
            I => \RTD.cfg_tmp_2\
        );

    \I__2609\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22443\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__22443\,
            I => \RTD.cfg_tmp_3\
        );

    \I__2607\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22437\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__22437\,
            I => \RTD.cfg_tmp_4\
        );

    \I__2605\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22431\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__22431\,
            I => \RTD.cfg_tmp_5\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22425\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22425\,
            I => \RTD.cfg_tmp_6\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__22422\,
            I => \N__22418\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__22421\,
            I => \N__22415\
        );

    \I__2599\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22406\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22383\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22383\
        );

    \I__2596\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22383\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22383\
        );

    \I__2594\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22383\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22410\,
            I => \N__22383\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22409\,
            I => \N__22383\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22380\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22370\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22370\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22361\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22402\,
            I => \N__22361\
        );

    \I__2586\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22361\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22361\
        );

    \I__2584\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22356\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22356\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22353\
        );

    \I__2581\ : Span4Mux_v
    port map (
            O => \N__22380\,
            I => \N__22347\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22344\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__22378\,
            I => \N__22333\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__22377\,
            I => \N__22328\
        );

    \I__2577\ : InMux
    port map (
            O => \N__22376\,
            I => \N__22324\
        );

    \I__2576\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22321\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22314\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__22361\,
            I => \N__22314\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__22356\,
            I => \N__22314\
        );

    \I__2572\ : Span4Mux_v
    port map (
            O => \N__22353\,
            I => \N__22311\
        );

    \I__2571\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22308\
        );

    \I__2570\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22305\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22302\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__22347\,
            I => \N__22297\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22297\
        );

    \I__2566\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22284\
        );

    \I__2565\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22284\
        );

    \I__2564\ : InMux
    port map (
            O => \N__22341\,
            I => \N__22284\
        );

    \I__2563\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22284\
        );

    \I__2562\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22284\
        );

    \I__2561\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22284\
        );

    \I__2560\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22269\
        );

    \I__2559\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22269\
        );

    \I__2558\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22269\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22269\
        );

    \I__2556\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22269\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22269\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22269\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22262\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__22321\,
            I => \N__22262\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__22314\,
            I => \N__22262\
        );

    \I__2550\ : Sp12to4
    port map (
            O => \N__22311\,
            I => \N__22257\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__22308\,
            I => \N__22257\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__22305\,
            I => \RTD.adc_state_0\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__22302\,
            I => \RTD.adc_state_0\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__22297\,
            I => \RTD.adc_state_0\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__22284\,
            I => \RTD.adc_state_0\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__22269\,
            I => \RTD.adc_state_0\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__22262\,
            I => \RTD.adc_state_0\
        );

    \I__2542\ : Odrv12
    port map (
            O => \N__22257\,
            I => \RTD.adc_state_0\
        );

    \I__2541\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__22239\,
            I => \N__22236\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__22236\,
            I => \N__22232\
        );

    \I__2538\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22229\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__22232\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__22229\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2535\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22198\
        );

    \I__2534\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22198\
        );

    \I__2533\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22198\
        );

    \I__2532\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22198\
        );

    \I__2531\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22198\
        );

    \I__2530\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22198\
        );

    \I__2529\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22198\
        );

    \I__2528\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22198\
        );

    \I__2527\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22189\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__22215\,
            I => \N__22183\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__22198\,
            I => \N__22170\
        );

    \I__2524\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22157\
        );

    \I__2523\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22157\
        );

    \I__2522\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22157\
        );

    \I__2521\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22157\
        );

    \I__2520\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22157\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__22192\,
            I => \N__22149\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__22189\,
            I => \N__22146\
        );

    \I__2517\ : InMux
    port map (
            O => \N__22188\,
            I => \N__22141\
        );

    \I__2516\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22141\
        );

    \I__2515\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22138\
        );

    \I__2514\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22135\
        );

    \I__2513\ : InMux
    port map (
            O => \N__22182\,
            I => \N__22130\
        );

    \I__2512\ : InMux
    port map (
            O => \N__22181\,
            I => \N__22130\
        );

    \I__2511\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22125\
        );

    \I__2510\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22125\
        );

    \I__2509\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22116\
        );

    \I__2508\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22116\
        );

    \I__2507\ : InMux
    port map (
            O => \N__22176\,
            I => \N__22116\
        );

    \I__2506\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22116\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__22174\,
            I => \N__22112\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__22173\,
            I => \N__22108\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__22170\,
            I => \N__22105\
        );

    \I__2502\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22102\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__22168\,
            I => \N__22099\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__22157\,
            I => \N__22091\
        );

    \I__2499\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22080\
        );

    \I__2498\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22080\
        );

    \I__2497\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22080\
        );

    \I__2496\ : InMux
    port map (
            O => \N__22153\,
            I => \N__22080\
        );

    \I__2495\ : InMux
    port map (
            O => \N__22152\,
            I => \N__22080\
        );

    \I__2494\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22077\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__22146\,
            I => \N__22074\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__22141\,
            I => \N__22069\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__22138\,
            I => \N__22069\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__22135\,
            I => \N__22063\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22058\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__22125\,
            I => \N__22058\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__22116\,
            I => \N__22055\
        );

    \I__2486\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22052\
        );

    \I__2485\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22047\
        );

    \I__2484\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22047\
        );

    \I__2483\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22044\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__22105\,
            I => \N__22039\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__22102\,
            I => \N__22039\
        );

    \I__2480\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22034\
        );

    \I__2479\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22034\
        );

    \I__2478\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22025\
        );

    \I__2477\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22025\
        );

    \I__2476\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22025\
        );

    \I__2475\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22025\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__22091\,
            I => \N__22014\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22014\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__22077\,
            I => \N__22014\
        );

    \I__2471\ : Span4Mux_h
    port map (
            O => \N__22074\,
            I => \N__22014\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__22069\,
            I => \N__22014\
        );

    \I__2469\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22007\
        );

    \I__2468\ : InMux
    port map (
            O => \N__22067\,
            I => \N__22007\
        );

    \I__2467\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22007\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__22063\,
            I => \N__22000\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__22058\,
            I => \N__22000\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__22055\,
            I => \N__22000\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__22052\,
            I => adc_state_2
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__22047\,
            I => adc_state_2
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__22044\,
            I => adc_state_2
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__22039\,
            I => adc_state_2
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__22034\,
            I => adc_state_2
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__22025\,
            I => adc_state_2
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__22014\,
            I => adc_state_2
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__22007\,
            I => adc_state_2
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__22000\,
            I => adc_state_2
        );

    \I__2454\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21978\,
            I => \RTD.cfg_tmp_0\
        );

    \I__2452\ : CEMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__21972\,
            I => \RTD.n13137\
        );

    \I__2450\ : SRMux
    port map (
            O => \N__21969\,
            I => \N__21966\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__21966\,
            I => \RTD.n15115\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__21963\,
            I => \N__21959\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21962\,
            I => \N__21956\
        );

    \I__2446\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21953\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21956\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__21953\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21948\,
            I => \ADC_IAC.n19833\
        );

    \I__2442\ : InMux
    port map (
            O => \N__21945\,
            I => \ADC_IAC.n19834\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21938\
        );

    \I__2440\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21935\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__21938\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21935\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__2437\ : CEMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__21927\,
            I => \N__21924\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__21924\,
            I => \N__21921\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__21921\,
            I => \ADC_IAC.n12698\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__21918\,
            I => \ADC_IAC.n12698_cascade_\
        );

    \I__2432\ : SRMux
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__21912\,
            I => \N__21909\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__21909\,
            I => \N__21906\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__21906\,
            I => \ADC_IAC.n15014\
        );

    \I__2428\ : IoInMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__21900\,
            I => \N__21897\
        );

    \I__2426\ : IoSpan4Mux
    port map (
            O => \N__21897\,
            I => \N__21894\
        );

    \I__2425\ : IoSpan4Mux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__2424\ : Span4Mux_s3_v
    port map (
            O => \N__21891\,
            I => \N__21888\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__21888\,
            I => \N__21885\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__21885\,
            I => \AC_ADC_SYNC\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__21882\,
            I => \n14_adj_1662_cascade_\
        );

    \I__2420\ : IoInMux
    port map (
            O => \N__21879\,
            I => \N__21876\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__2418\ : Span4Mux_s3_v
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__21870\,
            I => \N__21866\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21863\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__21866\,
            I => \IAC_CS\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21863\,
            I => \IAC_CS\
        );

    \I__2413\ : IoInMux
    port map (
            O => \N__21858\,
            I => \N__21855\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21855\,
            I => \N__21852\
        );

    \I__2411\ : Span4Mux_s3_v
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__21849\,
            I => \N__21846\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__21846\,
            I => \N__21843\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__21843\,
            I => \DDS_CS1\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__21840\,
            I => \ADC_IAC.n21458_cascade_\
        );

    \I__2406\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__21834\,
            I => \ADC_IAC.n16\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21827\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21830\,
            I => \N__21824\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__21827\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21824\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__2400\ : InMux
    port map (
            O => \N__21819\,
            I => \bfn_6_18_0_\
        );

    \I__2399\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21812\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21809\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__21812\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21809\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__2395\ : InMux
    port map (
            O => \N__21804\,
            I => \ADC_IAC.n19828\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21797\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21794\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21797\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__21794\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21789\,
            I => \ADC_IAC.n19829\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21782\
        );

    \I__2388\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21779\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__21782\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21779\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__2385\ : InMux
    port map (
            O => \N__21774\,
            I => \ADC_IAC.n19830\
        );

    \I__2384\ : InMux
    port map (
            O => \N__21771\,
            I => \N__21767\
        );

    \I__2383\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21764\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21767\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__21764\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21759\,
            I => \ADC_IAC.n19831\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__21756\,
            I => \N__21752\
        );

    \I__2378\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21749\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21746\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__21749\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__21746\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__2374\ : InMux
    port map (
            O => \N__21741\,
            I => \ADC_IAC.n19832\
        );

    \I__2373\ : CEMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__21732\,
            I => \ADC_VAC.n12\
        );

    \I__2370\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21726\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__21726\,
            I => n21050
        );

    \I__2368\ : CascadeMux
    port map (
            O => \N__21723\,
            I => \N__21719\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__21722\,
            I => \N__21716\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21710\
        );

    \I__2365\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21707\
        );

    \I__2364\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21704\
        );

    \I__2363\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21701\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__21713\,
            I => \N__21698\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__21710\,
            I => \N__21695\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21707\,
            I => \N__21692\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__21704\,
            I => \N__21689\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21686\
        );

    \I__2357\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21683\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__21695\,
            I => \N__21678\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__21692\,
            I => \N__21678\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__21689\,
            I => \N__21671\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__21686\,
            I => \N__21671\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21671\
        );

    \I__2351\ : Sp12to4
    port map (
            O => \N__21678\,
            I => \N__21666\
        );

    \I__2350\ : Sp12to4
    port map (
            O => \N__21671\,
            I => \N__21666\
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__21666\,
            I => \VAC_DRDY\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__21663\,
            I => \n21050_cascade_\
        );

    \I__2347\ : IoInMux
    port map (
            O => \N__21660\,
            I => \N__21657\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__21657\,
            I => \N__21654\
        );

    \I__2345\ : Span4Mux_s3_h
    port map (
            O => \N__21654\,
            I => \N__21651\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__21651\,
            I => \N__21647\
        );

    \I__2343\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21644\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__21647\,
            I => \N__21641\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__21644\,
            I => \N__21638\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__21641\,
            I => \VAC_CS\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__21638\,
            I => \VAC_CS\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21630\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21630\,
            I => n14_adj_1657
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__21627\,
            I => \N__21622\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__21626\,
            I => \N__21613\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__21625\,
            I => \N__21609\
        );

    \I__2333\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21604\
        );

    \I__2332\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21601\
        );

    \I__2331\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21598\
        );

    \I__2330\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21595\
        );

    \I__2329\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21592\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21587\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21587\
        );

    \I__2326\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21576\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21576\
        );

    \I__2324\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21576\
        );

    \I__2323\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21576\
        );

    \I__2322\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21576\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__21604\,
            I => \N__21569\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__21601\,
            I => \N__21569\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__21598\,
            I => \N__21569\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__21595\,
            I => \DTRIG_N_958_adj_1493\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__21592\,
            I => \DTRIG_N_958_adj_1493\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__21587\,
            I => \DTRIG_N_958_adj_1493\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__21576\,
            I => \DTRIG_N_958_adj_1493\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__21569\,
            I => \DTRIG_N_958_adj_1493\
        );

    \I__2313\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21547\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21547\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21544\
        );

    \I__2310\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21536\
        );

    \I__2309\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21533\
        );

    \I__2308\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21528\
        );

    \I__2307\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21528\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__21547\,
            I => \N__21523\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__21544\,
            I => \N__21523\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21543\,
            I => \N__21512\
        );

    \I__2303\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21512\
        );

    \I__2302\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21512\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21512\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21512\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__21536\,
            I => adc_state_1_adj_1459
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__21533\,
            I => adc_state_1_adj_1459
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__21528\,
            I => adc_state_1_adj_1459
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__21523\,
            I => adc_state_1_adj_1459
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21512\,
            I => adc_state_1_adj_1459
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__21501\,
            I => \N__21498\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21493\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__21497\,
            I => \N__21490\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__21496\,
            I => \N__21487\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21484\
        );

    \I__2289\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21479\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21479\
        );

    \I__2287\ : Odrv12
    port map (
            O => \N__21484\,
            I => cmd_rdadctmp_14
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__21479\,
            I => cmd_rdadctmp_14
        );

    \I__2285\ : InMux
    port map (
            O => \N__21474\,
            I => \N__21471\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__21471\,
            I => \ADC_VAC.n17\
        );

    \I__2283\ : IoInMux
    port map (
            O => \N__21468\,
            I => \N__21465\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21462\
        );

    \I__2281\ : IoSpan4Mux
    port map (
            O => \N__21462\,
            I => \N__21459\
        );

    \I__2280\ : Span4Mux_s2_h
    port map (
            O => \N__21459\,
            I => \N__21455\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__21458\,
            I => \N__21452\
        );

    \I__2278\ : Span4Mux_h
    port map (
            O => \N__21455\,
            I => \N__21449\
        );

    \I__2277\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21446\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__21449\,
            I => \VAC_SCLK\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__21446\,
            I => \VAC_SCLK\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__21441\,
            I => \N__21437\
        );

    \I__2273\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21429\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21429\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21429\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__21429\,
            I => cmd_rdadctmp_26_adj_1466
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__21426\,
            I => \N__21423\
        );

    \I__2268\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21420\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21417\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__21417\,
            I => \N__21413\
        );

    \I__2265\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21410\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__21413\,
            I => cmd_rdadctmp_3_adj_1489
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21410\,
            I => cmd_rdadctmp_3_adj_1489
        );

    \I__2262\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21402\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__21402\,
            I => \N__21399\
        );

    \I__2260\ : Span4Mux_h
    port map (
            O => \N__21399\,
            I => \N__21395\
        );

    \I__2259\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21391\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__21395\,
            I => \N__21388\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21385\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__21391\,
            I => buf_adcdata_iac_7
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__21388\,
            I => buf_adcdata_iac_7
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21385\,
            I => buf_adcdata_iac_7
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__21378\,
            I => \N__21374\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__21377\,
            I => \N__21371\
        );

    \I__2251\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__2250\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21364\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__21368\,
            I => \N__21361\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21358\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21364\,
            I => cmd_rdadctmp_8_adj_1484
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__21361\,
            I => cmd_rdadctmp_8_adj_1484
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__21358\,
            I => cmd_rdadctmp_8_adj_1484
        );

    \I__2244\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21348\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21345\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__21345\,
            I => \N__21342\
        );

    \I__2241\ : Sp12to4
    port map (
            O => \N__21342\,
            I => \N__21339\
        );

    \I__2240\ : Odrv12
    port map (
            O => \N__21339\,
            I => buf_data_iac_7
        );

    \I__2239\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__21333\,
            I => n22_adj_1598
        );

    \I__2237\ : InMux
    port map (
            O => \N__21330\,
            I => \N__21323\
        );

    \I__2236\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21323\
        );

    \I__2235\ : InMux
    port map (
            O => \N__21328\,
            I => \N__21320\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__21323\,
            I => cmd_rdadctmp_12_adj_1480
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21320\,
            I => cmd_rdadctmp_12_adj_1480
        );

    \I__2232\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21311\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__21314\,
            I => \N__21308\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__21311\,
            I => \N__21304\
        );

    \I__2229\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21301\
        );

    \I__2228\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21298\
        );

    \I__2227\ : Span12Mux_s9_h
    port map (
            O => \N__21304\,
            I => \N__21295\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__21301\,
            I => buf_adcdata_iac_4
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__21298\,
            I => buf_adcdata_iac_4
        );

    \I__2224\ : Odrv12
    port map (
            O => \N__21295\,
            I => buf_adcdata_iac_4
        );

    \I__2223\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21284\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__21287\,
            I => \N__21281\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__21284\,
            I => \N__21278\
        );

    \I__2220\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21274\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__21278\,
            I => \N__21271\
        );

    \I__2218\ : InMux
    port map (
            O => \N__21277\,
            I => \N__21268\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__21274\,
            I => buf_adcdata_vac_4
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__21271\,
            I => buf_adcdata_vac_4
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__21268\,
            I => buf_adcdata_vac_4
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__21261\,
            I => \n19_adj_1606_cascade_\
        );

    \I__2213\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21255\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__21252\,
            I => \N__21249\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__21249\,
            I => \N__21246\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__21246\,
            I => buf_data_iac_4
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__21243\,
            I => \n22_adj_1607_cascade_\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__2206\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21233\
        );

    \I__2205\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21230\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__21233\,
            I => cmd_rdadctmp_31_adj_1461
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__21230\,
            I => cmd_rdadctmp_31_adj_1461
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__2201\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__21219\,
            I => \N__21215\
        );

    \I__2199\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21212\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__21215\,
            I => \N__21206\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__21212\,
            I => \N__21206\
        );

    \I__2196\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21203\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__21206\,
            I => read_buf_0
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__21203\,
            I => read_buf_0
        );

    \I__2193\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21193\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__21197\,
            I => \N__21190\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__21196\,
            I => \N__21187\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__21193\,
            I => \N__21184\
        );

    \I__2189\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21179\
        );

    \I__2188\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21179\
        );

    \I__2187\ : Odrv12
    port map (
            O => \N__21184\,
            I => read_buf_2
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__21179\,
            I => read_buf_2
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__21174\,
            I => \N__21170\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__21173\,
            I => \N__21166\
        );

    \I__2183\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21156\
        );

    \I__2182\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21156\
        );

    \I__2181\ : InMux
    port map (
            O => \N__21166\,
            I => \N__21142\
        );

    \I__2180\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21142\
        );

    \I__2179\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21142\
        );

    \I__2178\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21137\
        );

    \I__2177\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21137\
        );

    \I__2176\ : InMux
    port map (
            O => \N__21161\,
            I => \N__21134\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21131\
        );

    \I__2174\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21126\
        );

    \I__2173\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21126\
        );

    \I__2172\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21115\
        );

    \I__2171\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21115\
        );

    \I__2170\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21115\
        );

    \I__2169\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21115\
        );

    \I__2168\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21115\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__21142\,
            I => n11856
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__21137\,
            I => n11856
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__21134\,
            I => n11856
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__21131\,
            I => n11856
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__21126\,
            I => n11856
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__21115\,
            I => n11856
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__21102\,
            I => \N__21097\
        );

    \I__2160\ : InMux
    port map (
            O => \N__21101\,
            I => \N__21092\
        );

    \I__2159\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21092\
        );

    \I__2158\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21089\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__21092\,
            I => read_buf_1
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__21089\,
            I => read_buf_1
        );

    \I__2155\ : InMux
    port map (
            O => \N__21084\,
            I => \N__21079\
        );

    \I__2154\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21074\
        );

    \I__2153\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21074\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__21079\,
            I => read_buf_12
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__21074\,
            I => read_buf_12
        );

    \I__2150\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21064\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__21068\,
            I => \N__21061\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__21067\,
            I => \N__21058\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21055\
        );

    \I__2146\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21050\
        );

    \I__2145\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21050\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__21055\,
            I => read_buf_13
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__21050\,
            I => read_buf_13
        );

    \I__2142\ : InMux
    port map (
            O => \N__21045\,
            I => \N__21035\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__21044\,
            I => \N__21032\
        );

    \I__2140\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21018\
        );

    \I__2139\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21018\
        );

    \I__2138\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21018\
        );

    \I__2137\ : InMux
    port map (
            O => \N__21040\,
            I => \N__21011\
        );

    \I__2136\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21011\
        );

    \I__2135\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21011\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__21035\,
            I => \N__21008\
        );

    \I__2133\ : InMux
    port map (
            O => \N__21032\,
            I => \N__21005\
        );

    \I__2132\ : InMux
    port map (
            O => \N__21031\,
            I => \N__20996\
        );

    \I__2131\ : InMux
    port map (
            O => \N__21030\,
            I => \N__20996\
        );

    \I__2130\ : InMux
    port map (
            O => \N__21029\,
            I => \N__20996\
        );

    \I__2129\ : InMux
    port map (
            O => \N__21028\,
            I => \N__20996\
        );

    \I__2128\ : InMux
    port map (
            O => \N__21027\,
            I => \N__20989\
        );

    \I__2127\ : InMux
    port map (
            O => \N__21026\,
            I => \N__20989\
        );

    \I__2126\ : InMux
    port map (
            O => \N__21025\,
            I => \N__20989\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__21018\,
            I => n13212
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__21011\,
            I => n13212
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__21008\,
            I => n13212
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__21005\,
            I => n13212
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__20996\,
            I => n13212
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20989\,
            I => n13212
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__20976\,
            I => \N__20971\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__20975\,
            I => \N__20965\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__20974\,
            I => \N__20962\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20952\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20952\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20952\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20946\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20935\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20935\
        );

    \I__2110\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20935\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20935\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20935\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20932\
        );

    \I__2106\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20925\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20925\
        );

    \I__2104\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20925\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20918\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20935\,
            I => \N__20915\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__20932\,
            I => \N__20910\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20910\
        );

    \I__2099\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20903\
        );

    \I__2098\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20903\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20903\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20900\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__20918\,
            I => \N__20895\
        );

    \I__2094\ : Span4Mux_v
    port map (
            O => \N__20915\,
            I => \N__20895\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__20910\,
            I => \N__20892\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20887\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20900\,
            I => \N__20887\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__20895\,
            I => n1_adj_1592
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__20892\,
            I => n1_adj_1592
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__20887\,
            I => n1_adj_1592
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__20880\,
            I => \N__20877\
        );

    \I__2086\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20873\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20869\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20866\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20863\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20869\,
            I => read_buf_6
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__20866\,
            I => read_buf_6
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__20863\,
            I => read_buf_6
        );

    \I__2079\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20851\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20846\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20846\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__20851\,
            I => read_buf_7
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__20846\,
            I => read_buf_7
        );

    \I__2074\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20838\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20838\,
            I => \N__20835\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__20835\,
            I => \N__20831\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20827\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__20831\,
            I => \N__20824\
        );

    \I__2069\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20821\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__20827\,
            I => buf_adcdata_iac_6
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__20824\,
            I => buf_adcdata_iac_6
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__20821\,
            I => buf_adcdata_iac_6
        );

    \I__2065\ : SRMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__20811\,
            I => \N__20807\
        );

    \I__2063\ : SRMux
    port map (
            O => \N__20810\,
            I => \N__20804\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__20807\,
            I => \N__20801\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__20804\,
            I => \N__20798\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__20801\,
            I => \N__20795\
        );

    \I__2059\ : Span4Mux_h
    port map (
            O => \N__20798\,
            I => \N__20790\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__20795\,
            I => \N__20790\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__20790\,
            I => \RTD.n20370\
        );

    \I__2056\ : InMux
    port map (
            O => \N__20787\,
            I => \N__20783\
        );

    \I__2055\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20780\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__20783\,
            I => \RTD.cfg_buf_6\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__20780\,
            I => \RTD.cfg_buf_6\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__20775\,
            I => \N__20771\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__20774\,
            I => \N__20768\
        );

    \I__2050\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20764\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20759\
        );

    \I__2048\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20759\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__20764\,
            I => read_buf_9
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__20759\,
            I => read_buf_9
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__20754\,
            I => \N__20745\
        );

    \I__2044\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20735\
        );

    \I__2043\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20735\
        );

    \I__2042\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20735\
        );

    \I__2041\ : InMux
    port map (
            O => \N__20750\,
            I => \N__20730\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20749\,
            I => \N__20730\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20718\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20718\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20718\
        );

    \I__2036\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20713\
        );

    \I__2035\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20713\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__20735\,
            I => \N__20706\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__20730\,
            I => \N__20706\
        );

    \I__2032\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20697\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20697\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20697\
        );

    \I__2029\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20697\
        );

    \I__2028\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20694\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__20718\,
            I => \N__20691\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20688\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20680\
        );

    \I__2024\ : InMux
    port map (
            O => \N__20711\,
            I => \N__20680\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__20706\,
            I => \N__20674\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20674\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__20694\,
            I => \N__20666\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__20691\,
            I => \N__20666\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__20688\,
            I => \N__20663\
        );

    \I__2018\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20656\
        );

    \I__2017\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20656\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20685\,
            I => \N__20656\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20653\
        );

    \I__2014\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20650\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__20674\,
            I => \N__20647\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20640\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20640\
        );

    \I__2010\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20640\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__20666\,
            I => \RTD.adc_state_1\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__20663\,
            I => \RTD.adc_state_1\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__20656\,
            I => \RTD.adc_state_1\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__20653\,
            I => \RTD.adc_state_1\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__20650\,
            I => \RTD.adc_state_1\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__20647\,
            I => \RTD.adc_state_1\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__20640\,
            I => \RTD.adc_state_1\
        );

    \I__2002\ : CEMux
    port map (
            O => \N__20625\,
            I => \N__20622\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__20619\,
            I => \N__20616\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__20616\,
            I => \N__20613\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__20613\,
            I => \RTD.n11829\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__20610\,
            I => \N__20605\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__20609\,
            I => \N__20602\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__20608\,
            I => \N__20599\
        );

    \I__1994\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20592\
        );

    \I__1993\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20592\
        );

    \I__1992\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20592\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__20592\,
            I => read_buf_8
        );

    \I__1990\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20583\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__20583\,
            I => \N__20576\
        );

    \I__1987\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20571\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20571\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20566\
        );

    \I__1984\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20566\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__20576\,
            I => \RTD.bit_cnt_3\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__20571\,
            I => \RTD.bit_cnt_3\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20566\,
            I => \RTD.bit_cnt_3\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20556\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__20556\,
            I => \N__20551\
        );

    \I__1978\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20548\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20545\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__20551\,
            I => \RTD.n18043\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__20548\,
            I => \RTD.n18043\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__20545\,
            I => \RTD.n18043\
        );

    \I__1973\ : InMux
    port map (
            O => \N__20538\,
            I => \N__20535\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20531\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20528\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__20531\,
            I => \N__20525\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20522\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__20525\,
            I => \RTD.n19026\
        );

    \I__1967\ : Odrv12
    port map (
            O => \N__20522\,
            I => \RTD.n19026\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \N__20513\
        );

    \I__1965\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20510\
        );

    \I__1964\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20507\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__20510\,
            I => adress_6
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__20507\,
            I => adress_6
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__20502\,
            I => \RTD.n9_cascade_\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__20499\,
            I => \RTD.adress_7_N_1086_7_cascade_\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20491\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20488\
        );

    \I__1957\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20485\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__20491\,
            I => \N__20482\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N__20479\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__20485\,
            I => \N__20476\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__20482\,
            I => \N__20469\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__20479\,
            I => \N__20469\
        );

    \I__1951\ : Span4Mux_v
    port map (
            O => \N__20476\,
            I => \N__20469\
        );

    \I__1950\ : Sp12to4
    port map (
            O => \N__20469\,
            I => \N__20466\
        );

    \I__1949\ : Span12Mux_v
    port map (
            O => \N__20466\,
            I => \N__20463\
        );

    \I__1948\ : Odrv12
    port map (
            O => \N__20463\,
            I => \RTD_DRDY\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__20460\,
            I => \RTD.n11_cascade_\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__20457\,
            I => \RTD.n19_cascade_\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__20454\,
            I => \N__20451\
        );

    \I__1944\ : InMux
    port map (
            O => \N__20451\,
            I => \N__20447\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__20450\,
            I => \N__20444\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__20447\,
            I => \N__20441\
        );

    \I__1941\ : InMux
    port map (
            O => \N__20444\,
            I => \N__20438\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__20441\,
            I => \N__20435\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__20438\,
            I => \RTD.adress_7\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__20435\,
            I => \RTD.adress_7\
        );

    \I__1937\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20424\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20419\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20419\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20427\,
            I => \N__20416\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20424\,
            I => \RTD.adress_7_N_1086_7\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20419\,
            I => \RTD.adress_7_N_1086_7\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__20416\,
            I => \RTD.adress_7_N_1086_7\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__20409\,
            I => \N__20406\
        );

    \I__1929\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__20400\,
            I => adress_0
        );

    \I__1926\ : CEMux
    port map (
            O => \N__20397\,
            I => \N__20394\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__20394\,
            I => \N__20385\
        );

    \I__1924\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20372\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20372\
        );

    \I__1922\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20372\
        );

    \I__1921\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20372\
        );

    \I__1920\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20372\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20372\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__20385\,
            I => n13054
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__20372\,
            I => n13054
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__20367\,
            I => \ADC_VAC.n21157_cascade_\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20364\,
            I => \N__20361\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20361\,
            I => \ADC_VAC.n21468\
        );

    \I__1913\ : CEMux
    port map (
            O => \N__20358\,
            I => \N__20355\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__20355\,
            I => \N__20352\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__20352\,
            I => \N__20349\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__20349\,
            I => \ADC_VAC.n21158\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__20346\,
            I => \N__20342\
        );

    \I__1908\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20339\
        );

    \I__1907\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20336\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__20339\,
            I => \N__20333\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20330\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__20333\,
            I => \N__20327\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__20330\,
            I => \RTD.n16766\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__20327\,
            I => \RTD.n16766\
        );

    \I__1901\ : IoInMux
    port map (
            O => \N__20322\,
            I => \N__20319\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__20319\,
            I => \N__20316\
        );

    \I__1899\ : IoSpan4Mux
    port map (
            O => \N__20316\,
            I => \N__20313\
        );

    \I__1898\ : IoSpan4Mux
    port map (
            O => \N__20313\,
            I => \N__20310\
        );

    \I__1897\ : Span4Mux_s3_h
    port map (
            O => \N__20310\,
            I => \N__20307\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__20307\,
            I => \N__20304\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__20304\,
            I => \N__20301\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__20301\,
            I => \RTD_CS\
        );

    \I__1893\ : InMux
    port map (
            O => \N__20298\,
            I => \N__20295\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20292\
        );

    \I__1891\ : Span4Mux_h
    port map (
            O => \N__20292\,
            I => \N__20289\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__20289\,
            I => \RTD.n14\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__20286\,
            I => \RTD.n21181_cascade_\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__20283\,
            I => \RTD.n13137_cascade_\
        );

    \I__1887\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20276\
        );

    \I__1886\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20273\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__20276\,
            I => \N__20268\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__20273\,
            I => \N__20268\
        );

    \I__1883\ : Span4Mux_v
    port map (
            O => \N__20268\,
            I => \N__20265\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__20265\,
            I => \RTD.n7889\
        );

    \I__1881\ : InMux
    port map (
            O => \N__20262\,
            I => \ADC_VAC.n19838\
        );

    \I__1880\ : InMux
    port map (
            O => \N__20259\,
            I => \ADC_VAC.n19839\
        );

    \I__1879\ : InMux
    port map (
            O => \N__20256\,
            I => \ADC_VAC.n19840\
        );

    \I__1878\ : InMux
    port map (
            O => \N__20253\,
            I => \ADC_VAC.n19841\
        );

    \I__1877\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20246\
        );

    \I__1876\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20243\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__20246\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__20243\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__1873\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20234\
        );

    \I__1872\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20231\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__20234\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__20231\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__20226\,
            I => \N__20222\
        );

    \I__1868\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20219\
        );

    \I__1867\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20216\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__20219\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__20216\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__1864\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20207\
        );

    \I__1863\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20204\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__20207\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__20204\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__1860\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20195\
        );

    \I__1859\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20192\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20189\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__20192\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__20189\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__1855\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20180\
        );

    \I__1854\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20177\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__20180\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__20177\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__20172\,
            I => \ADC_VAC.n21224_cascade_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20165\
        );

    \I__1849\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20162\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__20165\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__20162\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__1846\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20153\
        );

    \I__1845\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20150\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__20153\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__20150\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__20145\,
            I => \ADC_VAC.n21234_cascade_\
        );

    \I__1841\ : CEMux
    port map (
            O => \N__20142\,
            I => \N__20139\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20135\
        );

    \I__1839\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20132\
        );

    \I__1838\ : Sp12to4
    port map (
            O => \N__20135\,
            I => \N__20127\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__20132\,
            I => \N__20127\
        );

    \I__1836\ : Odrv12
    port map (
            O => \N__20127\,
            I => \ADC_VAC.n12803\
        );

    \I__1835\ : SRMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__1833\ : Span4Mux_h
    port map (
            O => \N__20118\,
            I => \N__20115\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__20115\,
            I => \ADC_VAC.n15052\
        );

    \I__1831\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20106\
        );

    \I__1830\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20106\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__20106\,
            I => cmd_rdadctmp_7_adj_1485
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__20103\,
            I => \N__20100\
        );

    \I__1827\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20097\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__20097\,
            I => \N__20094\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__20094\,
            I => \N__20091\
        );

    \I__1824\ : Sp12to4
    port map (
            O => \N__20091\,
            I => \N__20088\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__20088\,
            I => \VAC_MISO\
        );

    \I__1822\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20079\
        );

    \I__1821\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20079\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__20079\,
            I => cmd_rdadctmp_0_adj_1492
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__20076\,
            I => \N__20073\
        );

    \I__1818\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20067\
        );

    \I__1817\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20067\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__20067\,
            I => cmd_rdadctmp_1_adj_1491
        );

    \I__1815\ : InMux
    port map (
            O => \N__20064\,
            I => \N__20058\
        );

    \I__1814\ : InMux
    port map (
            O => \N__20063\,
            I => \N__20058\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__20058\,
            I => cmd_rdadctmp_2_adj_1490
        );

    \I__1812\ : InMux
    port map (
            O => \N__20055\,
            I => \bfn_5_14_0_\
        );

    \I__1811\ : InMux
    port map (
            O => \N__20052\,
            I => \ADC_VAC.n19835\
        );

    \I__1810\ : InMux
    port map (
            O => \N__20049\,
            I => \ADC_VAC.n19836\
        );

    \I__1809\ : InMux
    port map (
            O => \N__20046\,
            I => \ADC_VAC.n19837\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__20043\,
            I => \n19_adj_1597_cascade_\
        );

    \I__1807\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20037\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__20034\,
            I => \N__20029\
        );

    \I__1804\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20024\
        );

    \I__1803\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20024\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__20029\,
            I => buf_adcdata_vac_7
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__20024\,
            I => buf_adcdata_vac_7
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__20019\,
            I => \N__20014\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__20018\,
            I => \N__20011\
        );

    \I__1798\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20004\
        );

    \I__1797\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20004\
        );

    \I__1796\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20004\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__20004\,
            I => read_buf_4
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__20001\,
            I => \N__19996\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__20000\,
            I => \N__19993\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19988\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19988\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19985\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19982\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__19985\,
            I => read_buf_11
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19982\,
            I => read_buf_11
        );

    \I__1786\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19969\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19964\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19964\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__19969\,
            I => read_buf_5
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__19964\,
            I => read_buf_5
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__19959\,
            I => \N__19955\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__19958\,
            I => \N__19951\
        );

    \I__1778\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19948\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19943\
        );

    \I__1776\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19943\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__19948\,
            I => read_buf_3
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__19943\,
            I => read_buf_3
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__19938\,
            I => \n19_adj_1600_cascade_\
        );

    \I__1772\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__19932\,
            I => \N__19927\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19922\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19930\,
            I => \N__19922\
        );

    \I__1768\ : Odrv12
    port map (
            O => \N__19927\,
            I => read_buf_10
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__19922\,
            I => read_buf_10
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__19917\,
            I => \n13212_cascade_\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__19914\,
            I => \N__19911\
        );

    \I__1764\ : InMux
    port map (
            O => \N__19911\,
            I => \N__19905\
        );

    \I__1763\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19905\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__19905\,
            I => read_buf_15
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__19902\,
            I => \n11856_cascade_\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__19899\,
            I => \N__19894\
        );

    \I__1759\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19889\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19889\
        );

    \I__1757\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19886\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__19889\,
            I => read_buf_14
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__19886\,
            I => read_buf_14
        );

    \I__1754\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__19875\,
            I => \RTD.n12_adj_1445\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__19872\,
            I => \N__19869\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19863\
        );

    \I__1749\ : InMux
    port map (
            O => \N__19868\,
            I => \N__19858\
        );

    \I__1748\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19858\
        );

    \I__1747\ : InMux
    port map (
            O => \N__19866\,
            I => \N__19855\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19852\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19847\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__19855\,
            I => \N__19847\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__19852\,
            I => \N__19844\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__19847\,
            I => \RTD.mode\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__19844\,
            I => \RTD.mode\
        );

    \I__1740\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19833\
        );

    \I__1739\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19833\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__19833\,
            I => adress_5
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__19830\,
            I => \N__19827\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19824\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__19815\,
            I => \N__19812\
        );

    \I__1731\ : Sp12to4
    port map (
            O => \N__19812\,
            I => \N__19809\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__19809\,
            I => \RTD_SDO\
        );

    \I__1729\ : CEMux
    port map (
            O => \N__19806\,
            I => \N__19803\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__1727\ : Odrv12
    port map (
            O => \N__19800\,
            I => \RTD.n11915\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__19797\,
            I => \N__19792\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \N__19789\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19783\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19792\,
            I => \N__19772\
        );

    \I__1722\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19772\
        );

    \I__1721\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19772\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19787\,
            I => \N__19772\
        );

    \I__1719\ : InMux
    port map (
            O => \N__19786\,
            I => \N__19772\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__19783\,
            I => n14692
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19772\,
            I => n14692
        );

    \I__1716\ : SRMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__19764\,
            I => \N__19761\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__19761\,
            I => \RTD.n15280\
        );

    \I__1713\ : CEMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19752\
        );

    \I__1711\ : Span12Mux_v
    port map (
            O => \N__19752\,
            I => \N__19749\
        );

    \I__1710\ : Odrv12
    port map (
            O => \N__19749\,
            I => \RTD.n11860\
        );

    \I__1709\ : CEMux
    port map (
            O => \N__19746\,
            I => \N__19743\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__19740\,
            I => \RTD.n8\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__1705\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19730\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19727\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__19730\,
            I => adress_1
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__19727\,
            I => adress_1
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__1700\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19713\
        );

    \I__1699\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19713\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__19710\,
            I => adress_2
        );

    \I__1696\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19701\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19701\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__19701\,
            I => adress_3
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__19698\,
            I => \N__19695\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19689\
        );

    \I__1691\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19689\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__19689\,
            I => adress_4
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__1688\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19680\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__19680\,
            I => \RTD.n19032\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__19677\,
            I => \RTD.n4_cascade_\
        );

    \I__1685\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19671\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__19671\,
            I => \RTD.n21387\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__19668\,
            I => \RTD.n21199_cascade_\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19662\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19658\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19655\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__19658\,
            I => \RTD.adc_state_3_N_1114_1\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__19655\,
            I => \RTD.adc_state_3_N_1114_1\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__19650\,
            I => \RTD.n7_cascade_\
        );

    \I__1676\ : CEMux
    port map (
            O => \N__19647\,
            I => \N__19644\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__19644\,
            I => \N__19640\
        );

    \I__1674\ : CEMux
    port map (
            O => \N__19643\,
            I => \N__19637\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__19640\,
            I => \N__19632\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19637\,
            I => \N__19632\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__19632\,
            I => \RTD.n11868\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__19629\,
            I => \RTD.n21492_cascade_\
        );

    \I__1669\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__19620\,
            I => \RTD.n7_adj_1435\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__19617\,
            I => \N__19614\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19607\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19607\
        );

    \I__1663\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19604\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19607\,
            I => \RTD.bit_cnt_2\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__19604\,
            I => \RTD.bit_cnt_2\
        );

    \I__1660\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19589\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19589\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19589\
        );

    \I__1657\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19586\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__19589\,
            I => \RTD.bit_cnt_1\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__19586\,
            I => \RTD.bit_cnt_1\
        );

    \I__1654\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19568\
        );

    \I__1653\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19568\
        );

    \I__1652\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19568\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19568\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19565\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19568\,
            I => \RTD.bit_cnt_0\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__19565\,
            I => \RTD.bit_cnt_0\
        );

    \I__1647\ : IoInMux
    port map (
            O => \N__19560\,
            I => \N__19557\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__1645\ : Span4Mux_s2_h
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__1644\ : Sp12to4
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__1643\ : Span12Mux_v
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__1642\ : Odrv12
    port map (
            O => \N__19545\,
            I => \RTD_SDI\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__19542\,
            I => \RTD.n21471_cascade_\
        );

    \I__1640\ : IoInMux
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__1638\ : IoSpan4Mux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1637\ : Span4Mux_s3_h
    port map (
            O => \N__19530\,
            I => \N__19527\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__19527\,
            I => \N__19524\
        );

    \I__1635\ : Span4Mux_v
    port map (
            O => \N__19524\,
            I => \N__19521\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__19521\,
            I => \RTD_SCLK\
        );

    \I__1633\ : SRMux
    port map (
            O => \N__19518\,
            I => \N__19515\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__19515\,
            I => \CLK_DDS.n16974\
        );

    \I__1631\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19501\
        );

    \I__1630\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19501\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19501\
        );

    \I__1628\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19496\
        );

    \I__1627\ : InMux
    port map (
            O => \N__19508\,
            I => \N__19496\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__19501\,
            I => bit_cnt_0_adj_1498
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__19496\,
            I => bit_cnt_0_adj_1498
        );

    \I__1624\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19487\
        );

    \I__1623\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19484\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__19487\,
            I => bit_cnt_3
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__19484\,
            I => bit_cnt_3
        );

    \I__1620\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19474\
        );

    \I__1619\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19471\
        );

    \I__1618\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19468\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__19474\,
            I => bit_cnt_2
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__19471\,
            I => bit_cnt_2
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__19468\,
            I => bit_cnt_2
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__1613\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19450\
        );

    \I__1612\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19450\
        );

    \I__1611\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19447\
        );

    \I__1610\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19444\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__19450\,
            I => bit_cnt_1
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__19447\,
            I => bit_cnt_1
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__19444\,
            I => bit_cnt_1
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \n8_adj_1680_cascade_\
        );

    \I__1605\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19431\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__19431\,
            I => n21625
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__19428\,
            I => \RTD.n18043_cascade_\
        );

    \I__1602\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__19422\,
            I => \RTD.n21494\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19416\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__19416\,
            I => \RTD.n18092\
        );

    \I__1598\ : IoInMux
    port map (
            O => \N__19413\,
            I => \N__19410\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__1596\ : IoSpan4Mux
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__1595\ : IoSpan4Mux
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__19401\,
            I => \ICE_SYSCLK\
        );

    \I__1593\ : IoInMux
    port map (
            O => \N__19398\,
            I => \N__19395\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__1591\ : IoSpan4Mux
    port map (
            O => \N__19392\,
            I => \N__19389\
        );

    \I__1590\ : Span4Mux_s3_v
    port map (
            O => \N__19389\,
            I => \N__19386\
        );

    \I__1589\ : Sp12to4
    port map (
            O => \N__19386\,
            I => \N__19383\
        );

    \I__1588\ : Span12Mux_h
    port map (
            O => \N__19383\,
            I => \N__19380\
        );

    \I__1587\ : Odrv12
    port map (
            O => \N__19380\,
            I => \ICE_GPMO_2\
        );

    \INVADC_VDC.genclk.t0on_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i8C_net\,
            I => \N__50798\
        );

    \INVADC_VDC.genclk.t0on_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i0C_net\,
            I => \N__50797\
        );

    \INVADC_VDC.genclk.div_state_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i0C_net\,
            I => \N__50796\
        );

    \INVADC_VDC.genclk.t0off_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i8C_net\,
            I => \N__50795\
        );

    \INVADC_VDC.genclk.t0off_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i0C_net\,
            I => \N__50794\
        );

    \INVADC_VDC.genclk.div_state_i1C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i1C_net\,
            I => \N__50793\
        );

    \INVdds0_mclkcnt_i7_3772__i0C\ : INV
    port map (
            O => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            I => \N__50803\
        );

    \INVdds0_mclk_294C\ : INV
    port map (
            O => \INVdds0_mclk_294C_net\,
            I => \N__50799\
        );

    \INVcomm_spi.data_valid_85C\ : INV
    port map (
            O => \INVcomm_spi.data_valid_85C_net\,
            I => \N__55969\
        );

    \INVcomm_spi.MISO_48_12291_12292_setC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12291_12292_setC_net\,
            I => \N__55941\
        );

    \INVcomm_spi.MISO_48_12291_12292_resetC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12291_12292_resetC_net\,
            I => \N__55939\
        );

    \INVcomm_spi.imiso_83_12297_12298_setC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12297_12298_setC_net\,
            I => \N__58307\
        );

    \INVdata_cntvec_i0_i8C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i8C_net\,
            I => \N__56006\
        );

    \INVdata_cntvec_i0_i0C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i0C_net\,
            I => \N__55992\
        );

    \INVcomm_spi.bit_cnt_3767__i3C\ : INV
    port map (
            O => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            I => \N__58391\
        );

    \INVADC_VDC.genclk.t_clk_24C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t_clk_24C_net\,
            I => \N__50781\
        );

    \INVcomm_spi.imiso_83_12297_12298_resetC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12297_12298_resetC_net\,
            I => \N__58357\
        );

    \INVacadc_skipcnt_i0_i9C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i9C_net\,
            I => \N__56078\
        );

    \INVacadc_skipcnt_i0_i1C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i1C_net\,
            I => \N__56065\
        );

    \INVacadc_skipcnt_i0_i0C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i0C_net\,
            I => \N__56052\
        );

    \INVdata_count_i0_i8C\ : INV
    port map (
            O => \INVdata_count_i0_i8C_net\,
            I => \N__56045\
        );

    \INVdata_count_i0_i0C\ : INV
    port map (
            O => \INVdata_count_i0_i0C_net\,
            I => \N__56029\
        );

    \INVeis_state_i0C\ : INV
    port map (
            O => \INVeis_state_i0C_net\,
            I => \N__55990\
        );

    \INVeis_state_i1C\ : INV
    port map (
            O => \INVeis_state_i1C_net\,
            I => \N__56020\
        );

    \INVacadc_trig_300C\ : INV
    port map (
            O => \INVacadc_trig_300C_net\,
            I => \N__56003\
        );

    \INViac_raw_buf_vac_raw_buf_merged2WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            I => \N__56043\
        );

    \INViac_raw_buf_vac_raw_buf_merged7WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            I => \N__56103\
        );

    \INViac_raw_buf_vac_raw_buf_merged1WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            I => \N__55961\
        );

    \INViac_raw_buf_vac_raw_buf_merged6WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            I => \N__56101\
        );

    \INViac_raw_buf_vac_raw_buf_merged0WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            I => \N__55949\
        );

    \INViac_raw_buf_vac_raw_buf_merged5WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            I => \N__56098\
        );

    \INViac_raw_buf_vac_raw_buf_merged9WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            I => \N__55998\
        );

    \INViac_raw_buf_vac_raw_buf_merged4WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            I => \N__56091\
        );

    \INViac_raw_buf_vac_raw_buf_merged8WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            I => \N__55973\
        );

    \INViac_raw_buf_vac_raw_buf_merged10WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            I => \N__55985\
        );

    \INViac_raw_buf_vac_raw_buf_merged3WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            I => \N__56072\
        );

    \INViac_raw_buf_vac_raw_buf_merged11WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            I => \N__56013\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19939,
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19947,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19955,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19963,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19971,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_18_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_16_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \n19789_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_13_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19797,
            carryinitout => \bfn_13_20_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19781,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19772,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19820,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19811,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_19_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_7_0_\
        );

    \IN_MUX_bfv_19_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19895\,
            carryinitout => \bfn_19_8_0_\
        );

    \IN_MUX_bfv_22_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_7_0_\
        );

    \IN_MUX_bfv_22_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19910\,
            carryinitout => \bfn_22_8_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19884\,
            carryinitout => \bfn_10_7_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19849\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19857\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19865\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19873\,
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_18_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i3_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__19479\,
            in1 => \N__19512\,
            in2 => \N__19461\,
            in3 => \N__19491\,
            lcout => bit_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56028\,
            ce => \N__29821\,
            sr => \N__19518\
        );

    \CLK_DDS.bit_cnt_i2_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19457\,
            in1 => \N__19478\,
            in2 => \_gnd_net_\,
            in3 => \N__19511\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56028\,
            ce => \N__29821\,
            sr => \N__19518\
        );

    \CLK_DDS.bit_cnt_i1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19456\,
            in2 => \_gnd_net_\,
            in3 => \N__19510\,
            lcout => bit_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56028\,
            ce => \N__29821\,
            sr => \N__19518\
        );

    \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__22350\,
            in1 => \N__20279\,
            in2 => \N__22173\,
            in3 => \N__19425\,
            lcout => \RTD.n18092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i2_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30007\,
            in2 => \_gnd_net_\,
            in3 => \N__29819\,
            lcout => dds_state_2_adj_1494,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i0_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__22693\,
            in1 => \N__19419\,
            in2 => \_gnd_net_\,
            in3 => \N__19626\,
            lcout => \RTD.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40617\,
            ce => \N__19647\,
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100111"
        )
    port map (
            in0 => \N__22640\,
            in1 => \N__22111\,
            in2 => \N__19686\,
            in3 => \N__20538\,
            lcout => \RTD.adc_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40617\,
            ce => \N__19647\,
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i2_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__19674\,
            in1 => \N__20280\,
            in2 => \N__22174\,
            in3 => \N__22644\,
            lcout => adc_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40617\,
            ce => \N__19647\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__52285\,
            in1 => \N__54857\,
            in2 => \_gnd_net_\,
            in3 => \N__54554\,
            lcout => n14_adj_1578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.SCLK_51_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101111010100"
        )
    port map (
            in0 => \N__22351\,
            in1 => \N__20725\,
            in2 => \N__22678\,
            in3 => \N__22115\,
            lcout => \RTD_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40615\,
            ce => \N__19746\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i0_LC_3_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010101010"
        )
    port map (
            in0 => \N__19509\,
            in1 => \N__29910\,
            in2 => \N__30045\,
            in3 => \N__29791\,
            lcout => bit_cnt_0_adj_1498,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55996\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i1_3_lut_LC_3_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__30016\,
            in1 => \N__29909\,
            in2 => \_gnd_net_\,
            in3 => \N__29790\,
            lcout => \CLK_DDS.n16974\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19325_2_lut_LC_3_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19508\,
            in2 => \_gnd_net_\,
            in3 => \N__19490\,
            lcout => n21625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i3_3_lut_4_lut_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29907\,
            in1 => \N__19477\,
            in2 => \N__30031\,
            in3 => \N__19455\,
            lcout => OPEN,
            ltout => \n8_adj_1680_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i0_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000100010001"
        )
    port map (
            in0 => \N__29820\,
            in1 => \N__29908\,
            in2 => \N__19437\,
            in3 => \N__19434\,
            lcout => dds_state_0_adj_1496,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56014\,
            ce => \N__29718\,
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19612\,
            in1 => \N__19577\,
            in2 => \_gnd_net_\,
            in3 => \N__19596\,
            lcout => \RTD.n18043\,
            ltout => \RTD.n18043_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19370_3_lut_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__20580\,
            in1 => \_gnd_net_\,
            in2 => \N__19428\,
            in3 => \N__20711\,
            lcout => \RTD.n21494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19209_4_lut_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20579\,
            in1 => \N__20712\,
            in2 => \N__19872\,
            in3 => \N__20554\,
            lcout => OPEN,
            ltout => \RTD.n21492_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100110001"
        )
    port map (
            in0 => \N__22379\,
            in1 => \N__22169\,
            in2 => \N__19629\,
            in3 => \N__20534\,
            lcout => \RTD.n7_adj_1435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.bit_cnt_3769__i3_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__19599\,
            in1 => \N__20582\,
            in2 => \N__19617\,
            in3 => \N__19581\,
            lcout => \RTD.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40623\,
            ce => \N__19806\,
            sr => \N__19767\
        );

    \RTD.bit_cnt_3769__i2_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__19580\,
            in1 => \N__19613\,
            in2 => \_gnd_net_\,
            in3 => \N__19598\,
            lcout => \RTD.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40623\,
            ce => \N__19806\,
            sr => \N__19767\
        );

    \RTD.i1_2_lut_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__20555\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20581\,
            lcout => \RTD.adc_state_3_N_1114_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.bit_cnt_3769__i1_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19579\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19597\,
            lcout => \RTD.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40623\,
            ce => \N__19806\,
            sr => \N__19767\
        );

    \RTD.bit_cnt_3769__i0_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19578\,
            lcout => \RTD.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40623\,
            ce => \N__19806\,
            sr => \N__19767\
        );

    \i15467_2_lut_3_lut_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45479\,
            in1 => \N__54893\,
            in2 => \_gnd_net_\,
            in3 => \N__54514\,
            lcout => n14_adj_1548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.MOSI_59_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__22097\,
            in1 => \N__22343\,
            in2 => \N__20454\,
            in3 => \N__22242\,
            lcout => \RTD_SDI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40616\,
            ce => \N__19758\,
            sr => \N__20810\
        );

    \RTD.i19122_3_lut_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__22339\,
            in1 => \N__22512\,
            in2 => \_gnd_net_\,
            in3 => \N__20494\,
            lcout => OPEN,
            ltout => \RTD.n21471_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_10_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000000000"
        )
    port map (
            in0 => \N__22095\,
            in1 => \N__22639\,
            in2 => \N__19542\,
            in3 => \N__19868\,
            lcout => \RTD.n12_adj_1445\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i16510_3_lut_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011101"
        )
    port map (
            in0 => \N__22342\,
            in1 => \N__19866\,
            in2 => \_gnd_net_\,
            in3 => \N__22096\,
            lcout => \RTD.n19032\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_adj_19_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__22094\,
            in1 => \N__22635\,
            in2 => \_gnd_net_\,
            in3 => \N__22338\,
            lcout => n1_adj_1592,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_4_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22341\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => OPEN,
            ltout => \RTD.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19032_4_lut_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__22652\,
            in1 => \N__19867\,
            in2 => \N__19677\,
            in3 => \N__19661\,
            lcout => \RTD.n21387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_21_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22340\,
            in1 => \_gnd_net_\,
            in2 => \N__22677\,
            in3 => \_gnd_net_\,
            lcout => \RTD.n21061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i18472_2_lut_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20671\,
            in2 => \_gnd_net_\,
            in3 => \N__22066\,
            lcout => \RTD.n21199\,
            ltout => \RTD.n21199_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i3_4_lut_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__22331\,
            in1 => \N__22605\,
            in2 => \N__19668\,
            in3 => \N__20345\,
            lcout => \RTD.n11868\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011010110"
        )
    port map (
            in0 => \N__20685\,
            in1 => \N__22336\,
            in2 => \N__22168\,
            in3 => \N__19665\,
            lcout => OPEN,
            ltout => \RTD.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i1_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__22337\,
            in1 => \N__22610\,
            in2 => \N__19650\,
            in3 => \N__22516\,
            lcout => \RTD.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40538\,
            ce => \N__19643\,
            sr => \_gnd_net_\
        );

    \RTD.i27_4_lut_4_lut_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000110"
        )
    port map (
            in0 => \N__22098\,
            in1 => \N__20673\,
            in2 => \N__22645\,
            in3 => \N__22332\,
            lcout => \RTD.n11860\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19474_4_lut_4_lut_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111110111"
        )
    port map (
            in0 => \N__22068\,
            in1 => \N__22609\,
            in2 => \N__22378\,
            in3 => \N__20687\,
            lcout => \RTD.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i31_4_lut_3_lut_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22603\,
            in1 => \N__22327\,
            in2 => \_gnd_net_\,
            in3 => \N__20672\,
            lcout => \RTD.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__22067\,
            in1 => \N__22604\,
            in2 => \N__22377\,
            in3 => \N__20686\,
            lcout => \RTD.n20370\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i1_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19733\,
            in1 => \N__19786\,
            in2 => \N__20409\,
            in3 => \N__20388\,
            lcout => adress_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__20389\,
            in1 => \N__19718\,
            in2 => \N__19737\,
            in3 => \N__19795\,
            lcout => adress_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19706\,
            in1 => \N__19787\,
            in2 => \N__19722\,
            in3 => \N__20390\,
            lcout => adress_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i4_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__20391\,
            in1 => \N__19694\,
            in2 => \N__19796\,
            in3 => \N__19707\,
            lcout => adress_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19838\,
            in1 => \N__19788\,
            in2 => \N__19698\,
            in3 => \N__20392\,
            lcout => adress_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i6_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__20393\,
            in1 => \N__19839\,
            in2 => \N__19797\,
            in3 => \N__20516\,
            lcout => adress_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i0_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21211\,
            in1 => \N__20968\,
            in2 => \N__19830\,
            in3 => \N__21045\,
            lcout => read_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i11_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19931\,
            in1 => \N__20950\,
            in2 => \N__20000\,
            in3 => \N__21042\,
            lcout => read_buf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_8_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20495\,
            in2 => \_gnd_net_\,
            in3 => \N__20427\,
            lcout => \RTD.n16766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i14_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21069\,
            in1 => \N__20951\,
            in2 => \N__19899\,
            in3 => \N__21043\,
            lcout => read_buf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19471_4_lut_4_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011000111100"
        )
    port map (
            in0 => \N__22404\,
            in1 => \N__20748\,
            in2 => \N__22695\,
            in3 => \N__22188\,
            lcout => \RTD.n11915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i10_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19930\,
            in1 => \N__20949\,
            in2 => \N__20775\,
            in3 => \N__21041\,
            lcout => read_buf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12177_2_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20744\,
            lcout => n14692,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_3_lut_4_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010010100"
        )
    port map (
            in0 => \N__22187\,
            in1 => \N__22691\,
            in2 => \N__20754\,
            in3 => \N__22405\,
            lcout => \RTD.n15280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i6_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__43472\,
            in1 => \N__21165\,
            in2 => \N__20880\,
            in3 => \N__22156\,
            lcout => \buf_readRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i10_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__22153\,
            in1 => \N__19935\,
            in2 => \N__21173\,
            in3 => \N__23348\,
            lcout => \buf_readRTD_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010100000001"
        )
    port map (
            in0 => \N__20743\,
            in1 => \N__22375\,
            in2 => \N__22192\,
            in3 => \N__22670\,
            lcout => n13212,
            ltout => \n13212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i15_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__19898\,
            in1 => \N__19910\,
            in2 => \N__19917\,
            in3 => \N__20921\,
            lcout => read_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i15_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__27149\,
            in1 => \N__21164\,
            in2 => \N__19914\,
            in3 => \N__22155\,
            lcout => \buf_readRTD_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_16_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__22152\,
            in1 => \N__22376\,
            in2 => \N__22692\,
            in3 => \N__20742\,
            lcout => n11856,
            ltout => \n11856_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i14_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__22814\,
            in1 => \N__22154\,
            in2 => \N__19902\,
            in3 => \N__19897\,
            lcout => \buf_readRTD_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.mode_53_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__19881\,
            in1 => \N__22527\,
            in2 => \N__22971\,
            in3 => \N__20430\,
            lcout => \RTD.mode\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i4_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__22179\,
            in1 => \N__30620\,
            in2 => \N__20019\,
            in3 => \N__21161\,
            lcout => \buf_readRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i6_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__21029\,
            in1 => \N__19973\,
            in2 => \N__20975\,
            in3 => \N__20872\,
            lcout => read_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i12_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__21082\,
            in1 => \N__20959\,
            in2 => \N__21044\,
            in3 => \N__19999\,
            lcout => read_buf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i5_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__21028\,
            in1 => \N__19972\,
            in2 => \N__20974\,
            in3 => \N__20017\,
            lcout => read_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i4_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19954\,
            in1 => \N__20961\,
            in2 => \N__20018\,
            in3 => \N__21031\,
            lcout => read_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i12_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__35021\,
            in1 => \N__21155\,
            in2 => \N__22215\,
            in3 => \N__21083\,
            lcout => \buf_readRTD_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i3_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21198\,
            in1 => \N__20960\,
            in2 => \N__19958\,
            in3 => \N__21030\,
            lcout => read_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i11_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__25907\,
            in1 => \N__21154\,
            in2 => \N__20001\,
            in3 => \N__22180\,
            lcout => \buf_readRTD_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40569\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i5_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__22181\,
            in1 => \N__19977\,
            in2 => \N__21174\,
            in3 => \N__28283\,
            lcout => \buf_readRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__40805\,
            in1 => \N__21169\,
            in2 => \N__19959\,
            in3 => \N__22182\,
            lcout => \buf_readRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40612\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i19_3_lut_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25404\,
            in1 => \N__23138\,
            in2 => \_gnd_net_\,
            in3 => \N__57151\,
            lcout => OPEN,
            ltout => \n19_adj_1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i22_3_lut_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20830\,
            in2 => \N__19938\,
            in3 => \N__47515\,
            lcout => n22_adj_1601,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27974\,
            in1 => \N__27804\,
            in2 => \N__21377\,
            in3 => \N__27259\,
            lcout => buf_adcdata_vac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i19_3_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26766\,
            in1 => \N__20032\,
            in2 => \_gnd_net_\,
            in3 => \N__57260\,
            lcout => OPEN,
            ltout => \n19_adj_1597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i22_3_lut_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21394\,
            in2 => \N__20043\,
            in3 => \N__47694\,
            lcout => n22_adj_1598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i7_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27802\,
            in1 => \N__27977\,
            in2 => \N__23037\,
            in3 => \N__20033\,
            lcout => buf_adcdata_vac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i4_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27976\,
            in1 => \N__27805\,
            in2 => \N__21287\,
            in3 => \N__21330\,
            lcout => buf_adcdata_vac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i11_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__27803\,
            in1 => \N__23284\,
            in2 => \N__22799\,
            in3 => \N__28244\,
            lcout => cmd_rdadctmp_11_adj_1481,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i13_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__28245\,
            in1 => \N__21329\,
            in2 => \N__23227\,
            in3 => \N__27806\,
            lcout => cmd_rdadctmp_13_adj_1479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i23_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27801\,
            in1 => \N__27975\,
            in2 => \N__21240\,
            in3 => \N__27100\,
            lcout => buf_adcdata_vac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56059\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i3_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__28213\,
            in1 => \N__20064\,
            in2 => \N__27758\,
            in3 => \N__21416\,
            lcout => cmd_rdadctmp_3_adj_1489,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100010"
        )
    port map (
            in0 => \N__21620\,
            in1 => \N__27655\,
            in2 => \N__21722\,
            in3 => \N__21556\,
            lcout => \ADC_VAC.n12803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i8_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__28215\,
            in1 => \N__20112\,
            in2 => \N__27759\,
            in3 => \N__21367\,
            lcout => cmd_rdadctmp_8_adj_1484,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i7_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20111\,
            in1 => \N__27658\,
            in2 => \N__24690\,
            in3 => \N__28214\,
            lcout => cmd_rdadctmp_7_adj_1485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20084\,
            in1 => \N__27656\,
            in2 => \N__20103\,
            in3 => \N__28210\,
            lcout => cmd_rdadctmp_0_adj_1492,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28211\,
            in1 => \N__20072\,
            in2 => \N__27757\,
            in3 => \N__20085\,
            lcout => cmd_rdadctmp_1_adj_1491,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i2_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__20063\,
            in1 => \N__27657\,
            in2 => \N__20076\,
            in3 => \N__28212\,
            lcout => cmd_rdadctmp_2_adj_1490,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56073\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.bit_cnt_i0_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20184\,
            in2 => \_gnd_net_\,
            in3 => \N__20055\,
            lcout => \ADC_VAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \ADC_VAC.n19835\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i1_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20225\,
            in2 => \_gnd_net_\,
            in3 => \N__20052\,
            lcout => \ADC_VAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19835\,
            carryout => \ADC_VAC.n19836\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i2_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20211\,
            in2 => \_gnd_net_\,
            in3 => \N__20049\,
            lcout => \ADC_VAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19836\,
            carryout => \ADC_VAC.n19837\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20238\,
            in2 => \_gnd_net_\,
            in3 => \N__20046\,
            lcout => \ADC_VAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19837\,
            carryout => \ADC_VAC.n19838\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i4_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20250\,
            in2 => \_gnd_net_\,
            in3 => \N__20262\,
            lcout => \ADC_VAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19838\,
            carryout => \ADC_VAC.n19839\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i5_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20157\,
            in2 => \_gnd_net_\,
            in3 => \N__20259\,
            lcout => \ADC_VAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19839\,
            carryout => \ADC_VAC.n19840\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i6_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20198\,
            in2 => \_gnd_net_\,
            in3 => \N__20256\,
            lcout => \ADC_VAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19840\,
            carryout => \ADC_VAC.n19841\,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.bit_cnt_i7_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20169\,
            in2 => \_gnd_net_\,
            in3 => \N__20253\,
            lcout => \ADC_VAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56083\,
            ce => \N__20142\,
            sr => \N__20124\
        );

    \ADC_VAC.i18497_4_lut_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20249\,
            in1 => \N__20237\,
            in2 => \N__20226\,
            in3 => \N__20210\,
            lcout => OPEN,
            ltout => \ADC_VAC.n21224_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i18507_4_lut_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20199\,
            in1 => \N__20183\,
            in2 => \N__20172\,
            in3 => \N__20168\,
            lcout => OPEN,
            ltout => \ADC_VAC.n21234_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19109_4_lut_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27670\,
            in1 => \N__20156\,
            in2 => \N__20145\,
            in3 => \N__21552\,
            lcout => \ADC_VAC.n21468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i12536_2_lut_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__21617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20138\,
            lcout => \ADC_VAC.n15052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_adj_36_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111101111"
        )
    port map (
            in0 => \N__27668\,
            in1 => \N__21616\,
            in2 => \N__21723\,
            in3 => \N__28713\,
            lcout => OPEN,
            ltout => \ADC_VAC.n21157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_adj_37_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__21553\,
            in1 => \_gnd_net_\,
            in2 => \N__20367\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VAC.n21158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19419_2_lut_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27669\,
            in2 => \_gnd_net_\,
            in3 => \N__21474\,
            lcout => \ADC_VAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i0_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__21618\,
            in1 => \N__21555\,
            in2 => \N__27756\,
            in3 => \N__20364\,
            lcout => adc_state_0_adj_1460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56095\,
            ce => \N__20358\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30103\,
            in2 => \_gnd_net_\,
            in3 => \N__29941\,
            lcout => dds_state_1_adj_1495,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55955\,
            ce => \N__29711\,
            sr => \N__29844\
        );

    \RTD.CS_52_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101011111"
        )
    port map (
            in0 => \N__22399\,
            in1 => \N__20729\,
            in2 => \N__20346\,
            in3 => \N__22685\,
            lcout => \RTD_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40614\,
            ce => \N__20625\,
            sr => \_gnd_net_\
        );

    \RTD.i18454_2_lut_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22683\,
            in2 => \_gnd_net_\,
            in3 => \N__20726\,
            lcout => OPEN,
            ltout => \RTD.n21181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i30_4_lut_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110001000"
        )
    port map (
            in0 => \N__20298\,
            in1 => \N__22186\,
            in2 => \N__20286\,
            in3 => \N__22706\,
            lcout => \RTD.n13137\,
            ltout => \RTD.n13137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12599_2_lut_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20283\,
            in3 => \N__22684\,
            lcout => \RTD.n15115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_9_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__20728\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22398\,
            lcout => \RTD.n7889\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_adj_22_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__20727\,
            in1 => \N__20589\,
            in2 => \_gnd_net_\,
            in3 => \N__20559\,
            lcout => \RTD.n19026\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i7_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__22403\,
            in1 => \N__20753\,
            in2 => \N__20517\,
            in3 => \N__20429\,
            lcout => \RTD.adress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40608\,
            ce => \N__20397\,
            sr => \N__20814\
        );

    \RTD.i1_4_lut_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__25739\,
            in1 => \N__20786\,
            in2 => \N__27078\,
            in3 => \N__22902\,
            lcout => OPEN,
            ltout => \RTD.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i7_4_lut_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22476\,
            in1 => \N__22713\,
            in2 => \N__20502\,
            in3 => \N__22746\,
            lcout => \RTD.adress_7_N_1086_7\,
            ltout => \RTD.adress_7_N_1086_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_6_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20499\,
            in3 => \N__22400\,
            lcout => \RTD.n11\,
            ltout => \RTD.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i34_4_lut_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110011"
        )
    port map (
            in0 => \N__22401\,
            in1 => \N__20496\,
            in2 => \N__20460\,
            in3 => \N__20751\,
            lcout => OPEN,
            ltout => \RTD.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i35_4_lut_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__22544\,
            in1 => \N__22686\,
            in2 => \N__20457\,
            in3 => \N__22216\,
            lcout => n13054,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111110011"
        )
    port map (
            in0 => \N__22402\,
            in1 => \N__20752\,
            in2 => \N__20450\,
            in3 => \N__20428\,
            lcout => adress_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40608\,
            ce => \N__20397\,
            sr => \N__20814\
        );

    \RTD.i1_2_lut_3_lut_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__22352\,
            in1 => \N__20749\,
            in2 => \_gnd_net_\,
            in3 => \N__22175\,
            lcout => \RTD.n21036\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i8_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__22177\,
            in1 => \N__25817\,
            in2 => \N__20609\,
            in3 => \N__21163\,
            lcout => \buf_readRTD_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i9_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__21162\,
            in1 => \N__22886\,
            in2 => \N__20774\,
            in3 => \N__22178\,
            lcout => \buf_readRTD_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i6_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__22960\,
            in1 => \N__23008\,
            in2 => \N__27070\,
            in3 => \N__20787\,
            lcout => \RTD.cfg_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21038\,
            in1 => \N__21218\,
            in2 => \N__21102\,
            in3 => \N__20922\,
            lcout => read_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i9_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__20924\,
            in1 => \N__20767\,
            in2 => \N__20610\,
            in3 => \N__21040\,
            lcout => read_buf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19396_3_lut_3_lut_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__22679\,
            in1 => \N__20750\,
            in2 => \_gnd_net_\,
            in3 => \N__22176\,
            lcout => \RTD.n11829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i8_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20923\,
            in1 => \N__20856\,
            in2 => \N__20608\,
            in3 => \N__21039\,
            lcout => read_buf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i13_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__22193\,
            in1 => \N__34892\,
            in2 => \N__21068\,
            in3 => \N__21152\,
            lcout => \buf_readRTD_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i7_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__21151\,
            in1 => \N__22196\,
            in2 => \N__23723\,
            in3 => \N__20855\,
            lcout => \buf_readRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i2_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21101\,
            in1 => \N__20970\,
            in2 => \N__21196\,
            in3 => \N__21027\,
            lcout => read_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i0_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__21149\,
            in1 => \N__43697\,
            in2 => \N__21225\,
            in3 => \N__22197\,
            lcout => \buf_readRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__22194\,
            in1 => \N__35159\,
            in2 => \N__21197\,
            in3 => \N__21153\,
            lcout => \buf_readRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i1_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__21150\,
            in1 => \N__22195\,
            in2 => \N__28337\,
            in3 => \N__21100\,
            lcout => \buf_readRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i13_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__21084\,
            in1 => \N__20969\,
            in2 => \N__21067\,
            in3 => \N__21026\,
            lcout => read_buf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i7_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__21025\,
            in1 => \N__20854\,
            in2 => \N__20976\,
            in3 => \N__20876\,
            lcout => read_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40582\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38590\,
            in1 => \N__38751\,
            in2 => \N__23496\,
            in3 => \N__27223\,
            lcout => buf_adcdata_iac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i11_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38592\,
            in1 => \N__23527\,
            in2 => \N__24326\,
            in3 => \N__29392\,
            lcout => cmd_rdadctmp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i6_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38591\,
            in1 => \N__38753\,
            in2 => \N__21497\,
            in3 => \N__20834\,
            lcout => buf_adcdata_iac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i3_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38752\,
            in1 => \N__38594\,
            in2 => \N__23534\,
            in3 => \N__22846\,
            lcout => buf_adcdata_iac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i14_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38593\,
            in1 => \N__24353\,
            in2 => \N__21496\,
            in3 => \N__29393\,
            lcout => cmd_rdadctmp_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i22_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27973\,
            in1 => \N__27800\,
            in2 => \N__23099\,
            in3 => \N__23202\,
            lcout => buf_adcdata_vac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56016\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19316_2_lut_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__57187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31974\,
            lcout => n21705,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i19_3_lut_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__25608\,
            in1 => \_gnd_net_\,
            in2 => \N__57259\,
            in3 => \N__21277\,
            lcout => OPEN,
            ltout => \n19_adj_1606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i22_3_lut_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__21307\,
            in1 => \_gnd_net_\,
            in2 => \N__21261\,
            in3 => \N__47695\,
            lcout => OPEN,
            ltout => \n22_adj_1607_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i30_3_lut_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21258\,
            in2 => \N__21243\,
            in3 => \N__47091\,
            lcout => n30_adj_1608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i31_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__28191\,
            in1 => \N__23201\,
            in2 => \N__27847\,
            in3 => \N__21236\,
            lcout => cmd_rdadctmp_31_adj_1461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i14_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23053\,
            in1 => \N__27796\,
            in2 => \N__23228\,
            in3 => \N__28190\,
            lcout => cmd_rdadctmp_14_adj_1478,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i7_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38764\,
            in1 => \N__38598\,
            in2 => \N__26301\,
            in3 => \N__21398\,
            lcout => buf_adcdata_iac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i10_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22792\,
            in1 => \N__27723\,
            in2 => \N__23423\,
            in3 => \N__28187\,
            lcout => cmd_rdadctmp_10_adj_1482,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i9_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29383\,
            in1 => \N__36331\,
            in2 => \N__23489\,
            in3 => \N__38562\,
            lcout => cmd_rdadctmp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i9_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23416\,
            in1 => \N__27725\,
            in2 => \N__21378\,
            in3 => \N__28189\,
            lcout => cmd_rdadctmp_9_adj_1483,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i30_3_lut_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21351\,
            in1 => \N__21336\,
            in2 => \_gnd_net_\,
            in3 => \N__47048\,
            lcout => n30_adj_1599,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i12_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21328\,
            in1 => \N__27724\,
            in2 => \N__23297\,
            in3 => \N__28188\,
            lcout => cmd_rdadctmp_12_adj_1480,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i13_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38560\,
            in1 => \N__24346\,
            in2 => \N__23514\,
            in3 => \N__29384\,
            lcout => cmd_rdadctmp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i4_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38763\,
            in1 => \N__38561\,
            in2 => \N__21314\,
            in3 => \N__23513\,
            lcout => buf_adcdata_iac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i4_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__29452\,
            in1 => \N__46909\,
            in2 => \N__42714\,
            in3 => \N__46733\,
            lcout => buf_dds1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i3_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__50982\,
            in1 => \N__37536\,
            in2 => \N__47131\,
            in3 => \N__49878\,
            lcout => comm_cmd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i30_4_lut_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000010001"
        )
    port map (
            in0 => \N__28698\,
            in1 => \N__21621\,
            in2 => \N__21713\,
            in3 => \N__21557\,
            lcout => \ADC_VAC.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.DTRIG_39_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101000"
        )
    port map (
            in0 => \N__28846\,
            in1 => \N__21558\,
            in2 => \N__21627\,
            in3 => \N__27722\,
            lcout => acadc_dtrig_v,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i16_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__27721\,
            in1 => \N__26181\,
            in2 => \N__27964\,
            in3 => \N__25762\,
            lcout => buf_adcdata_vac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.CS_37_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__21729\,
            in1 => \N__21633\,
            in2 => \N__27755\,
            in3 => \N__21714\,
            lcout => \VAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i26_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21436\,
            in1 => \N__27645\,
            in2 => \N__26207\,
            in3 => \N__28130\,
            lcout => cmd_rdadctmp_26_adj_1466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.SCLK_35_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__27644\,
            in1 => \N__21619\,
            in2 => \N__21458\,
            in3 => \N__21554\,
            lcout => \VAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i27_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__25996\,
            in1 => \N__27646\,
            in2 => \N__21441\,
            in3 => \N__28131\,
            lcout => cmd_rdadctmp_27_adj_1465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i18_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27883\,
            in1 => \N__27650\,
            in2 => \N__24130\,
            in3 => \N__21440\,
            lcout => buf_adcdata_vac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28132\,
            in1 => \N__24713\,
            in2 => \N__21426\,
            in3 => \N__27651\,
            lcout => cmd_rdadctmp_4_adj_1488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i10_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24313\,
            in1 => \N__29380\,
            in2 => \N__36344\,
            in3 => \N__38563\,
            lcout => cmd_rdadctmp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i2_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__27630\,
            in1 => \N__21612\,
            in2 => \_gnd_net_\,
            in3 => \N__21542\,
            lcout => \DTRIG_N_958_adj_1493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56084\,
            ce => \N__21738\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i1_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__21543\,
            in1 => \_gnd_net_\,
            in2 => \N__21626\,
            in3 => \N__27631\,
            lcout => adc_state_1_adj_1459,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56084\,
            ce => \N__21738\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21607\,
            in2 => \_gnd_net_\,
            in3 => \N__21539\,
            lcout => n21050,
            ltout => \n21050_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_3_lut_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21715\,
            in2 => \N__21663\,
            in3 => \N__27628\,
            lcout => n12850,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_223_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110010"
        )
    port map (
            in0 => \N__21541\,
            in1 => \N__21650\,
            in2 => \N__21625\,
            in3 => \N__27629\,
            lcout => n14_adj_1657,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_61_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21608\,
            in2 => \_gnd_net_\,
            in3 => \N__21540\,
            lcout => n21076,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i15_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38408\,
            in1 => \N__26281\,
            in2 => \N__21501\,
            in3 => \N__29337\,
            lcout => cmd_rdadctmp_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i6_4_lut_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__24828\,
            in1 => \N__21830\,
            in2 => \N__21963\,
            in3 => \N__38406\,
            lcout => \ADC_IAC.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19194_4_lut_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21770\,
            in1 => \N__21785\,
            in2 => \N__21756\,
            in3 => \N__21800\,
            lcout => OPEN,
            ltout => \ADC_IAC.n21458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19307_4_lut_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21941\,
            in1 => \N__21816\,
            in2 => \N__21840\,
            in3 => \N__21837\,
            lcout => \ADC_IAC.n21457\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19411_2_lut_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38407\,
            in2 => \_gnd_net_\,
            in3 => \N__23757\,
            lcout => \ADC_IAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.bit_cnt_i0_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21831\,
            in2 => \_gnd_net_\,
            in3 => \N__21819\,
            lcout => \ADC_IAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_6_18_0_\,
            carryout => \ADC_IAC.n19828\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i1_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21815\,
            in2 => \_gnd_net_\,
            in3 => \N__21804\,
            lcout => \ADC_IAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19828\,
            carryout => \ADC_IAC.n19829\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i2_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21801\,
            in2 => \_gnd_net_\,
            in3 => \N__21789\,
            lcout => \ADC_IAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19829\,
            carryout => \ADC_IAC.n19830\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i3_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21786\,
            in2 => \_gnd_net_\,
            in3 => \N__21774\,
            lcout => \ADC_IAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19830\,
            carryout => \ADC_IAC.n19831\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i4_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21771\,
            in2 => \_gnd_net_\,
            in3 => \N__21759\,
            lcout => \ADC_IAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19831\,
            carryout => \ADC_IAC.n19832\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i5_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21755\,
            in2 => \_gnd_net_\,
            in3 => \N__21741\,
            lcout => \ADC_IAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19832\,
            carryout => \ADC_IAC.n19833\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i6_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21962\,
            in2 => \_gnd_net_\,
            in3 => \N__21948\,
            lcout => \ADC_IAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19833\,
            carryout => \ADC_IAC.n19834\,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.bit_cnt_i7_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21942\,
            in2 => \_gnd_net_\,
            in3 => \N__21945\,
            lcout => \ADC_IAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56096\,
            ce => \N__21930\,
            sr => \N__21915\
        );

    \ADC_IAC.i1_4_lut_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000100"
        )
    port map (
            in0 => \N__38457\,
            in1 => \N__24935\,
            in2 => \N__24615\,
            in3 => \N__24852\,
            lcout => \ADC_IAC.n12698\,
            ltout => \ADC_IAC.n12698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i12498_2_lut_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__24939\,
            in1 => \_gnd_net_\,
            in2 => \N__21918\,
            in3 => \_gnd_net_\,
            lcout => \ADC_IAC.n15014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_I_0_1_lut_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \AC_ADC_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_225_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110010"
        )
    port map (
            in0 => \N__24853\,
            in1 => \N__21869\,
            in2 => \N__24942\,
            in3 => \N__38458\,
            lcout => OPEN,
            ltout => \n14_adj_1662_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.CS_37_LC_6_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__38459\,
            in1 => \N__24606\,
            in2 => \N__21882\,
            in3 => \N__23799\,
            lcout => \IAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i3_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__24057\,
            in1 => \N__51413\,
            in2 => \N__22874\,
            in3 => \N__31626\,
            lcout => buf_adcdata_vdc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.CS_28_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__30102\,
            in1 => \N__29767\,
            in2 => \_gnd_net_\,
            in3 => \N__29942\,
            lcout => \DDS_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55951\,
            ce => \N__30123\,
            sr => \_gnd_net_\
        );

    \RTD.cfg_tmp_i1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__22217\,
            in1 => \N__22412\,
            in2 => \N__39600\,
            in3 => \N__21981\,
            lcout => \RTD.cfg_tmp_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__22410\,
            in1 => \N__22461\,
            in2 => \N__23334\,
            in3 => \N__22223\,
            lcout => \RTD.cfg_tmp_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__22218\,
            in1 => \N__22413\,
            in2 => \N__22455\,
            in3 => \N__25946\,
            lcout => \RTD.cfg_tmp_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i4_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__35010\,
            in1 => \N__22446\,
            in2 => \N__22421\,
            in3 => \N__22224\,
            lcout => \RTD.cfg_tmp_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i5_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__22221\,
            in1 => \N__22440\,
            in2 => \N__22422\,
            in3 => \N__34939\,
            lcout => \RTD.cfg_tmp_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__22411\,
            in1 => \N__22220\,
            in2 => \N__27077\,
            in3 => \N__22434\,
            lcout => \RTD.cfg_tmp_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i7_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__22219\,
            in1 => \N__22414\,
            in2 => \N__27024\,
            in3 => \N__22428\,
            lcout => \RTD.cfg_tmp_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_tmp_i0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__22409\,
            in1 => \N__22235\,
            in2 => \N__25740\,
            in3 => \N__22222\,
            lcout => \RTD.cfg_tmp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40622\,
            ce => \N__21975\,
            sr => \N__21969\
        );

    \RTD.cfg_buf_i4_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__22731\,
            in1 => \N__22949\,
            in2 => \N__23009\,
            in3 => \N__35008\,
            lcout => \RTD.cfg_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i5_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22755\,
            in1 => \N__23005\,
            in2 => \N__22968\,
            in3 => \N__34940\,
            lcout => \RTD.cfg_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i3_4_lut_adj_7_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__34941\,
            in1 => \N__22754\,
            in2 => \N__25947\,
            in3 => \N__22739\,
            lcout => \RTD.n11_adj_1444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i3_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__22740\,
            in1 => \N__22998\,
            in2 => \N__22967\,
            in3 => \N__25942\,
            lcout => \RTD.cfg_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i2_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__22722\,
            in1 => \N__22950\,
            in2 => \N__23010\,
            in3 => \N__23323\,
            lcout => \RTD.cfg_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_4_lut_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__35009\,
            in1 => \N__22730\,
            in2 => \N__23330\,
            in3 => \N__22721\,
            lcout => \RTD.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i22_4_lut_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__22707\,
            in1 => \N__22694\,
            in2 => \N__22545\,
            in3 => \N__22526\,
            lcout => \RTD.n13090\,
            ltout => \RTD.n13090_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__22948\,
            in1 => \N__39596\,
            in2 => \N__22491\,
            in3 => \N__22488\,
            lcout => \RTD.cfg_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4_4_lut_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__27017\,
            in1 => \N__22469\,
            in2 => \N__39595\,
            in3 => \N__22487\,
            lcout => \RTD.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i7_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22470\,
            in1 => \N__27016\,
            in2 => \N__22970\,
            in3 => \N__23007\,
            lcout => \RTD.cfg_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__25735\,
            in1 => \N__23006\,
            in2 => \N__22969\,
            in3 => \N__22901\,
            lcout => \RTD.cfg_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_1_i20_3_lut_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22887\,
            in1 => \N__39585\,
            in2 => \_gnd_net_\,
            in3 => \N__57196\,
            lcout => n20_adj_1693,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i19_3_lut_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57198\,
            in1 => \N__22875\,
            in2 => \_gnd_net_\,
            in3 => \N__23258\,
            lcout => OPEN,
            ltout => \n19_adj_1609_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i22_3_lut_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22853\,
            in2 => \N__22824\,
            in3 => \N__47500\,
            lcout => n22_adj_1610,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22407_bdd_4_lut_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__47501\,
            in1 => \N__23706\,
            in2 => \N__23697\,
            in3 => \N__23175\,
            lcout => n22410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19857_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__27060\,
            in1 => \N__57197\,
            in2 => \N__22821\,
            in3 => \N__46256\,
            lcout => n22629,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__28001\,
            in1 => \N__27850\,
            in2 => \N__22803\,
            in3 => \N__23159\,
            lcout => buf_adcdata_vac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55987\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i19_3_lut_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25437\,
            in1 => \N__23561\,
            in2 => \_gnd_net_\,
            in3 => \N__57091\,
            lcout => n19_adj_1652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.MOSI_31_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24396\,
            in1 => \N__22766\,
            in2 => \_gnd_net_\,
            in3 => \N__29822\,
            lcout => \DDS_MOSI1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55987\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19678_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__24099\,
            in1 => \N__46257\,
            in2 => \N__23184\,
            in3 => \N__47451\,
            lcout => n22407,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i19_3_lut_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57092\,
            in1 => \N__25647\,
            in2 => \_gnd_net_\,
            in3 => \N__23158\,
            lcout => OPEN,
            ltout => \n19_adj_1612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i22_3_lut_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24283\,
            in2 => \N__23145\,
            in3 => \N__47452\,
            lcout => n22_adj_1613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i6_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__28002\,
            in1 => \N__27851\,
            in2 => \N__23064\,
            in3 => \N__23137\,
            lcout => buf_adcdata_vac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55987\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15464_2_lut_3_lut_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45848\,
            in1 => \N__54884\,
            in2 => \_gnd_net_\,
            in3 => \N__54555\,
            lcout => n14_adj_1574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22629_bdd_4_lut_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__23092\,
            in1 => \N__23073\,
            in2 => \N__25686\,
            in3 => \N__46159\,
            lcout => n21237,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__23314\,
            in1 => \N__49312\,
            in2 => \N__45868\,
            in3 => \N__39663\,
            lcout => \buf_cfgRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i16_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__27848\,
            in1 => \N__26221\,
            in2 => \N__23030\,
            in3 => \N__28268\,
            lcout => cmd_rdadctmp_16_adj_1476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28267\,
            in1 => \N__23023\,
            in2 => \N__23060\,
            in3 => \N__27849\,
            lcout => cmd_rdadctmp_15_adj_1477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56000\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i30_3_lut_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47158\,
            in1 => \N__23403\,
            in2 => \_gnd_net_\,
            in3 => \N__23388\,
            lcout => n30_adj_1602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i30_3_lut_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23379\,
            in1 => \N__23358\,
            in2 => \_gnd_net_\,
            in3 => \N__47159\,
            lcout => n30_adj_1614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i20_3_lut_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56937\,
            in1 => \N__23352\,
            in2 => \_gnd_net_\,
            in3 => \N__23313\,
            lcout => n20_adj_1684,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i17_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23461\,
            in1 => \N__27794\,
            in2 => \N__26234\,
            in3 => \N__28246\,
            lcout => cmd_rdadctmp_17_adj_1475,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i3_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27791\,
            in1 => \N__27989\,
            in2 => \N__23298\,
            in3 => \N__23257\,
            lcout => buf_adcdata_vac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i5_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27990\,
            in1 => \N__27792\,
            in2 => \N__23235\,
            in3 => \N__24257\,
            lcout => buf_adcdata_vac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__50981\,
            in1 => \N__37522\,
            in2 => \N__49745\,
            in3 => \N__46224\,
            lcout => comm_cmd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i30_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__23200\,
            in1 => \N__27795\,
            in2 => \N__23448\,
            in3 => \N__28247\,
            lcout => cmd_rdadctmp_30_adj_1462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i21_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27790\,
            in1 => \N__27988\,
            in2 => \N__27421\,
            in3 => \N__23447\,
            lcout => buf_adcdata_vac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i9_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27991\,
            in1 => \N__27793\,
            in2 => \N__23466\,
            in3 => \N__23560\,
            lcout => buf_adcdata_vac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i12_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38558\,
            in1 => \N__23509\,
            in2 => \N__23538\,
            in3 => \N__29363\,
            lcout => cmd_rdadctmp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i8_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29362\,
            in1 => \N__23482\,
            in2 => \N__23667\,
            in3 => \N__38559\,
            lcout => cmd_rdadctmp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_dtrig_i_I_0_2_lut_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28826\,
            in2 => \_gnd_net_\,
            in3 => \N__28785\,
            lcout => \iac_raw_buf_N_776\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__27821\,
            in1 => \N__23465\,
            in2 => \N__26126\,
            in3 => \N__28254\,
            lcout => cmd_rdadctmp_18_adj_1474,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.DTRIG_39_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001000000"
        )
    port map (
            in0 => \N__38557\,
            in1 => \N__24854\,
            in2 => \N__24940\,
            in3 => \N__28786\,
            lcout => acadc_dtrig_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i29_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__27822\,
            in1 => \N__24412\,
            in2 => \N__23443\,
            in3 => \N__28256\,
            lcout => cmd_rdadctmp_29_adj_1463,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i28_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__28255\,
            in1 => \N__27823\,
            in2 => \N__24416\,
            in3 => \N__26003\,
            lcout => cmd_rdadctmp_28_adj_1464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27820\,
            in1 => \N__27965\,
            in2 => \N__23424\,
            in3 => \N__32162\,
            lcout => buf_adcdata_vac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i10_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30094\,
            in1 => \N__29845\,
            in2 => \N__23586\,
            in3 => \N__30873\,
            lcout => \CLK_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i11_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__29846\,
            in1 => \N__30098\,
            in2 => \N__23634\,
            in3 => \N__26442\,
            lcout => \CLK_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i12_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30095\,
            in1 => \N__29847\,
            in2 => \N__23625\,
            in3 => \N__36287\,
            lcout => \CLK_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i13_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__34960\,
            in1 => \N__23616\,
            in2 => \N__29872\,
            in3 => \N__30101\,
            lcout => \CLK_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i14_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30096\,
            in1 => \N__29851\,
            in2 => \N__23607\,
            in3 => \N__35637\,
            lcout => \CLK_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i15_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__29852\,
            in1 => \N__30099\,
            in2 => \N__23595\,
            in3 => \N__30897\,
            lcout => tmp_buf_15_adj_1497,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i9_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30097\,
            in1 => \N__29854\,
            in2 => \N__23577\,
            in3 => \N__32526\,
            lcout => \CLK_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i8_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__29853\,
            in1 => \N__30100\,
            in2 => \N__24540\,
            in3 => \N__39103\,
            lcout => \CLK_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56047\,
            ce => \N__30147\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i3_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__24474\,
            in1 => \N__24441\,
            in2 => \N__24498\,
            in3 => \N__36605\,
            lcout => \SIG_DDS.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56061\,
            ce => \N__44517\,
            sr => \N__24645\
        );

    \SIG_DDS.bit_cnt_i1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24439\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24497\,
            lcout => \SIG_DDS.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56061\,
            ce => \N__44517\,
            sr => \N__24645\
        );

    \i18636_3_lut_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23733\,
            in1 => \N__28389\,
            in2 => \_gnd_net_\,
            in3 => \N__46258\,
            lcout => n21363,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i2_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__24473\,
            in1 => \N__24493\,
            in2 => \_gnd_net_\,
            in3 => \N__24440\,
            lcout => \SIG_DDS.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56061\,
            ce => \N__44517\,
            sr => \N__24645\
        );

    \mux_128_Mux_1_i16_3_lut_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57269\,
            in1 => \N__32525\,
            in2 => \_gnd_net_\,
            in3 => \N__31253\,
            lcout => n16_adj_1690,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_1_i17_3_lut_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24749\,
            in1 => \N__26090\,
            in2 => \_gnd_net_\,
            in3 => \N__57268\,
            lcout => n17_adj_1691,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__38447\,
            in1 => \N__24908\,
            in2 => \_gnd_net_\,
            in3 => \N__24840\,
            lcout => \DTRIG_N_958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => \N__23682\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i1_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__24841\,
            in1 => \_gnd_net_\,
            in2 => \N__24927\,
            in3 => \N__38448\,
            lcout => adc_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56075\,
            ce => \N__23682\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_52_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24904\,
            in2 => \_gnd_net_\,
            in3 => \N__24839\,
            lcout => n21079,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i0_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__38446\,
            in1 => \N__24846\,
            in2 => \N__24928\,
            in3 => \N__23673\,
            lcout => adc_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56085\,
            ce => \N__25008\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i7_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23657\,
            in1 => \N__29328\,
            in2 => \N__23646\,
            in3 => \N__38401\,
            lcout => cmd_rdadctmp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i6_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__38399\,
            in1 => \N__23642\,
            in2 => \N__29374\,
            in3 => \N__23766\,
            lcout => cmd_rdadctmp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23789\,
            in1 => \N__29326\,
            in2 => \N__38564\,
            in3 => \N__24989\,
            lcout => cmd_rdadctmp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_226_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24918\,
            in2 => \_gnd_net_\,
            in3 => \N__24850\,
            lcout => n21082,
            ltout => \n21082_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_3_lut_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24616\,
            in2 => \N__23793\,
            in3 => \N__38397\,
            lcout => n12771,
            ltout => \n12771_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__38398\,
            in1 => \N__23790\,
            in2 => \N__23781\,
            in3 => \N__23774\,
            lcout => cmd_rdadctmp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__23765\,
            in1 => \N__29327\,
            in2 => \N__23778\,
            in3 => \N__38400\,
            lcout => cmd_rdadctmp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i30_4_lut_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001010001"
        )
    port map (
            in0 => \N__24926\,
            in1 => \N__24851\,
            in2 => \N__24623\,
            in3 => \N__28708\,
            lcout => \ADC_IAC.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_main.i19991_1_lut_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50810\,
            lcout => \DDS_MCLK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i18_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51476\,
            in1 => \N__31620\,
            in2 => \N__24155\,
            in3 => \N__24198\,
            lcout => buf_adcdata_vdc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i16_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__29082\,
            in1 => \N__24029\,
            in2 => \N__51758\,
            in3 => \N__25469\,
            lcout => cmd_rdadctmp_16_adj_1507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i17_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__24028\,
            in1 => \N__29084\,
            in2 => \N__51708\,
            in3 => \N__24004\,
            lcout => cmd_rdadctmp_17_adj_1506,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i19_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__23974\,
            in1 => \N__51640\,
            in2 => \N__29117\,
            in3 => \N__25258\,
            lcout => cmd_rdadctmp_19_adj_1504,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__51639\,
            in1 => \N__25301\,
            in2 => \N__23909\,
            in3 => \N__29093\,
            lcout => cmd_rdadctmp_6_adj_1517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__29083\,
            in1 => \N__23831\,
            in2 => \N__25074\,
            in3 => \N__51648\,
            lcout => cmd_rdadctmp_1_adj_1522,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__23830\,
            in1 => \N__51942\,
            in2 => \N__51707\,
            in3 => \N__29091\,
            lcout => cmd_rdadctmp_0_adj_1523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__23902\,
            in1 => \N__51641\,
            in2 => \N__29118\,
            in3 => \N__25277\,
            lcout => cmd_rdadctmp_7_adj_1516,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i18_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__51638\,
            in1 => \N__24005\,
            in2 => \N__23981\,
            in3 => \N__29092\,
            lcout => cmd_rdadctmp_18_adj_1505,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42365\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23814\,
            in2 => \N__23835\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.cmd_rdadcbuf_0\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \ADC_VDC.n19842\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23808\,
            in2 => \N__25072\,
            in3 => \N__23802\,
            lcout => \ADC_VDC.cmd_rdadcbuf_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19842\,
            carryout => \ADC_VDC.n19843\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23952\,
            in2 => \N__25047\,
            in3 => \N__23946\,
            lcout => \ADC_VDC.cmd_rdadcbuf_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19843\,
            carryout => \ADC_VDC.n19844\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23943\,
            in2 => \N__25029\,
            in3 => \N__23937\,
            lcout => \ADC_VDC.cmd_rdadcbuf_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19844\,
            carryout => \ADC_VDC.n19845\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25315\,
            in2 => \N__23934\,
            in3 => \N__23922\,
            lcout => \ADC_VDC.cmd_rdadcbuf_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19845\,
            carryout => \ADC_VDC.n19846\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23919\,
            in2 => \N__25302\,
            in3 => \N__23913\,
            lcout => \ADC_VDC.cmd_rdadcbuf_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19846\,
            carryout => \ADC_VDC.n19847\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23883\,
            in2 => \N__23910\,
            in3 => \N__23877\,
            lcout => \ADC_VDC.cmd_rdadcbuf_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19847\,
            carryout => \ADC_VDC.n19848\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25276\,
            in2 => \N__23874\,
            in3 => \N__23865\,
            lcout => \ADC_VDC.cmd_rdadcbuf_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19848\,
            carryout => \ADC_VDC.n19849\,
            clk => \N__42394\,
            ce => \N__26908\,
            sr => \N__26856\
        );

    \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23862\,
            in2 => \N__25238\,
            in3 => \N__23856\,
            lcout => \ADC_VDC.cmd_rdadcbuf_8\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \ADC_VDC.n19850\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23853\,
            in2 => \N__25215\,
            in3 => \N__23847\,
            lcout => \ADC_VDC.cmd_rdadcbuf_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19850\,
            carryout => \ADC_VDC.n19851\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23844\,
            in2 => \N__25194\,
            in3 => \N__23838\,
            lcout => \ADC_VDC.cmd_rdadcbuf_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19851\,
            carryout => \ADC_VDC.n19852\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25379\,
            in2 => \N__25167\,
            in3 => \N__24066\,
            lcout => cmd_rdadcbuf_11,
            ltout => OPEN,
            carryin => \ADC_VDC.n19852\,
            carryout => \ADC_VDC.n19853\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25147\,
            in2 => \N__31493\,
            in3 => \N__24063\,
            lcout => cmd_rdadcbuf_12,
            ltout => OPEN,
            carryin => \ADC_VDC.n19853\,
            carryout => \ADC_VDC.n19854\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25658\,
            in2 => \N__25126\,
            in3 => \N__24060\,
            lcout => cmd_rdadcbuf_13,
            ltout => OPEN,
            carryin => \ADC_VDC.n19854\,
            carryout => \ADC_VDC.n19855\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24050\,
            in2 => \N__25488\,
            in3 => \N__24039\,
            lcout => cmd_rdadcbuf_14,
            ltout => OPEN,
            carryin => \ADC_VDC.n19855\,
            carryout => \ADC_VDC.n19856\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25619\,
            in2 => \N__25470\,
            in3 => \N__24036\,
            lcout => cmd_rdadcbuf_15,
            ltout => OPEN,
            carryin => \ADC_VDC.n19856\,
            carryout => \ADC_VDC.n19857\,
            clk => \N__42411\,
            ce => \N__26946\,
            sr => \N__26853\
        );

    \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25586\,
            in2 => \N__24033\,
            in3 => \N__24012\,
            lcout => cmd_rdadcbuf_16,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \ADC_VDC.n19858\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25419\,
            in2 => \N__24009\,
            in3 => \N__23988\,
            lcout => cmd_rdadcbuf_17,
            ltout => OPEN,
            carryin => \ADC_VDC.n19858\,
            carryout => \ADC_VDC.n19859\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26777\,
            in2 => \N__23985\,
            in3 => \N__23955\,
            lcout => cmd_rdadcbuf_18,
            ltout => OPEN,
            carryin => \ADC_VDC.n19859\,
            carryout => \ADC_VDC.n19860\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25260\,
            in2 => \N__29666\,
            in3 => \N__24093\,
            lcout => cmd_rdadcbuf_19,
            ltout => OPEN,
            carryin => \ADC_VDC.n19860\,
            carryout => \ADC_VDC.n19861\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25448\,
            in2 => \N__25554\,
            in3 => \N__24090\,
            lcout => cmd_rdadcbuf_20,
            ltout => OPEN,
            carryin => \ADC_VDC.n19861\,
            carryout => \ADC_VDC.n19862\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25343\,
            in2 => \N__25529\,
            in3 => \N__24087\,
            lcout => cmd_rdadcbuf_21,
            ltout => OPEN,
            carryin => \ADC_VDC.n19862\,
            carryout => \ADC_VDC.n19863\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26705\,
            in2 => \N__30279\,
            in3 => \N__24084\,
            lcout => cmd_rdadcbuf_22,
            ltout => OPEN,
            carryin => \ADC_VDC.n19863\,
            carryout => \ADC_VDC.n19864\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26792\,
            in2 => \N__30243\,
            in3 => \N__24081\,
            lcout => cmd_rdadcbuf_23,
            ltout => OPEN,
            carryin => \ADC_VDC.n19864\,
            carryout => \ADC_VDC.n19865\,
            clk => \N__42384\,
            ce => \N__26930\,
            sr => \N__26854\
        );

    \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29642\,
            in2 => \_gnd_net_\,
            in3 => \N__24078\,
            lcout => cmd_rdadcbuf_24,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \ADC_VDC.n19866\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26720\,
            in2 => \_gnd_net_\,
            in3 => \N__24075\,
            lcout => cmd_rdadcbuf_25,
            ltout => OPEN,
            carryin => \ADC_VDC.n19866\,
            carryout => \ADC_VDC.n19867\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26738\,
            in2 => \_gnd_net_\,
            in3 => \N__24072\,
            lcout => cmd_rdadcbuf_26,
            ltout => OPEN,
            carryin => \ADC_VDC.n19867\,
            carryout => \ADC_VDC.n19868\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25100\,
            in2 => \_gnd_net_\,
            in3 => \N__24069\,
            lcout => cmd_rdadcbuf_27,
            ltout => OPEN,
            carryin => \ADC_VDC.n19868\,
            carryout => \ADC_VDC.n19869\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29564\,
            in2 => \_gnd_net_\,
            in3 => \N__24201\,
            lcout => cmd_rdadcbuf_28,
            ltout => OPEN,
            carryin => \ADC_VDC.n19869\,
            carryout => \ADC_VDC.n19870\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24191\,
            in2 => \_gnd_net_\,
            in3 => \N__24180\,
            lcout => cmd_rdadcbuf_29,
            ltout => OPEN,
            carryin => \ADC_VDC.n19870\,
            carryout => \ADC_VDC.n19871\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29600\,
            in2 => \_gnd_net_\,
            in3 => \N__24177\,
            lcout => cmd_rdadcbuf_30,
            ltout => OPEN,
            carryin => \ADC_VDC.n19871\,
            carryout => \ADC_VDC.n19872\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29474\,
            in2 => \_gnd_net_\,
            in3 => \N__24174\,
            lcout => cmd_rdadcbuf_31,
            ltout => OPEN,
            carryin => \ADC_VDC.n19872\,
            carryout => \ADC_VDC.n19873\,
            clk => \N__42412\,
            ce => \N__26941\,
            sr => \N__26868\
        );

    \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29519\,
            in2 => \_gnd_net_\,
            in3 => \N__24171\,
            lcout => cmd_rdadcbuf_32,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \ADC_VDC.n19874\,
            clk => \N__42434\,
            ce => \N__26945\,
            sr => \N__26855\
        );

    \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25328\,
            in2 => \_gnd_net_\,
            in3 => \N__24168\,
            lcout => cmd_rdadcbuf_33,
            ltout => OPEN,
            carryin => \ADC_VDC.n19874\,
            carryout => \ADC_VDC.n19875\,
            clk => \N__42434\,
            ce => \N__26945\,
            sr => \N__26855\
        );

    \ADC_VDC.add_23_36_lut_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25861\,
            in2 => \_gnd_net_\,
            in3 => \N__24165\,
            lcout => \ADC_VDC.cmd_rdadcbuf_35_N_1296_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i19_3_lut_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57148\,
            in1 => \N__24162\,
            in2 => \_gnd_net_\,
            in3 => \N__24131\,
            lcout => n19_adj_1683,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_1_i19_3_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29553\,
            in1 => \N__24521\,
            in2 => \_gnd_net_\,
            in3 => \N__57149\,
            lcout => n19_adj_1692,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i5_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__24227\,
            in1 => \N__24357\,
            in2 => \N__38607\,
            in3 => \N__38775\,
            lcout => buf_adcdata_iac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55988\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38774\,
            in1 => \N__38602\,
            in2 => \N__24290\,
            in3 => \N__24330\,
            lcout => buf_adcdata_iac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55988\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i19_3_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57150\,
            in1 => \N__25575\,
            in2 => \_gnd_net_\,
            in3 => \N__24253\,
            lcout => OPEN,
            ltout => \n19_adj_1603_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i22_3_lut_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24226\,
            in2 => \N__24213\,
            in3 => \N__47453\,
            lcout => n22_adj_1604,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i20_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__27500\,
            in1 => \N__27458\,
            in2 => \N__27858\,
            in3 => \N__28269\,
            lcout => cmd_rdadctmp_20_adj_1472,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55988\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i2_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__50994\,
            in1 => \N__37532\,
            in2 => \N__47537\,
            in3 => \N__50157\,
            lcout => comm_cmd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55988\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000110011"
        )
    port map (
            in0 => \N__36591\,
            in1 => \N__44702\,
            in2 => \N__24453\,
            in3 => \N__44516\,
            lcout => dds_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56001\,
            ce => \N__44550\,
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19668_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__47190\,
            in2 => \N__32580\,
            in3 => \N__47457\,
            lcout => OPEN,
            ltout => \n22377_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22377_bdd_4_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47191\,
            in1 => \N__30735\,
            in2 => \N__24210\,
            in3 => \N__24207\,
            lcout => n22380,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i1_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__49973\,
            in1 => \N__55461\,
            in2 => \N__49746\,
            in3 => \N__53141\,
            lcout => comm_buf_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i13_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011111100"
        )
    port map (
            in0 => \N__30723\,
            in1 => \N__46916\,
            in2 => \N__34967\,
            in3 => \N__55462\,
            lcout => buf_dds1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i5_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__55460\,
            in1 => \N__25364\,
            in2 => \N__37257\,
            in3 => \N__46915\,
            lcout => buf_dds1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i10_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27966\,
            in1 => \N__27827\,
            in2 => \N__27325\,
            in3 => \N__26122\,
            lcout => buf_adcdata_vac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i20_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27826\,
            in1 => \N__27967\,
            in2 => \N__24417\,
            in3 => \N__31859\,
            lcout => buf_adcdata_vac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i14_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__38750\,
            in1 => \N__43378\,
            in2 => \N__24669\,
            in3 => \N__38606\,
            lcout => buf_adcdata_iac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56018\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__29873\,
            in1 => \N__30108\,
            in2 => \N__41736\,
            in3 => \N__24392\,
            lcout => \CLK_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30104\,
            in1 => \N__29874\,
            in2 => \N__24381\,
            in3 => \N__35607\,
            lcout => \CLK_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__29875\,
            in1 => \N__24372\,
            in2 => \N__30114\,
            in3 => \N__26265\,
            lcout => \CLK_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30105\,
            in1 => \N__29876\,
            in2 => \N__24366\,
            in3 => \N__32688\,
            lcout => \CLK_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__29877\,
            in1 => \N__30109\,
            in2 => \N__24576\,
            in3 => \N__29456\,
            lcout => \CLK_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i5_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30106\,
            in1 => \N__29878\,
            in2 => \N__24567\,
            in3 => \N__25363\,
            lcout => \CLK_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__29879\,
            in1 => \N__30110\,
            in2 => \N__24558\,
            in3 => \N__46965\,
            lcout => \CLK_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i7_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__30107\,
            in1 => \N__29880\,
            in2 => \N__24549\,
            in3 => \N__36576\,
            lcout => \CLK_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56032\,
            ce => \N__30143\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i17_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27978\,
            in1 => \N__27824\,
            in2 => \N__26208\,
            in3 => \N__24520\,
            lcout => buf_adcdata_vac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i4_4_lut_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24492\,
            in1 => \N__24437\,
            in2 => \N__24472\,
            in3 => \N__44709\,
            lcout => \SIG_DDS.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i0_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__44508\,
            in1 => \_gnd_net_\,
            in2 => \N__24641\,
            in3 => \N__24438\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i8_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__39104\,
            in1 => \N__46914\,
            in2 => \N__45647\,
            in3 => \N__46754\,
            lcout => buf_dds1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i22_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__28089\,
            in1 => \N__27825\,
            in2 => \N__26347\,
            in3 => \N__28237\,
            lcout => cmd_rdadctmp_22_adj_1470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_292_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__46454\,
            in1 => \N__47193\,
            in2 => \_gnd_net_\,
            in3 => \N__47532\,
            lcout => n69,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i5_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24698\,
            in1 => \N__24720\,
            in2 => \N__27855\,
            in3 => \N__28185\,
            lcout => cmd_rdadctmp_5_adj_1487,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i22_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24658\,
            in1 => \N__29386\,
            in2 => \N__33114\,
            in3 => \N__38456\,
            lcout => cmd_rdadctmp_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i6_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24680\,
            in1 => \N__27778\,
            in2 => \N__24702\,
            in3 => \N__28186\,
            lcout => cmd_rdadctmp_6_adj_1486,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i22_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38640\,
            in1 => \N__38455\,
            in2 => \N__30778\,
            in3 => \N__26585\,
            lcout => buf_adcdata_iac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__38454\,
            in1 => \N__24659\,
            in2 => \N__29394\,
            in3 => \N__28738\,
            lcout => cmd_rdadctmp_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i12572_3_lut_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__44667\,
            in1 => \N__44708\,
            in2 => \_gnd_net_\,
            in3 => \N__44504\,
            lcout => n15092,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i28_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38403\,
            in1 => \N__28900\,
            in2 => \N__26408\,
            in3 => \N__29325\,
            lcout => cmd_rdadctmp_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i29_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29323\,
            in1 => \N__28960\,
            in2 => \N__28907\,
            in3 => \N__38404\,
            lcout => cmd_rdadctmp_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_adj_3_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__24903\,
            in1 => \N__38402\,
            in2 => \N__24624\,
            in3 => \N__28709\,
            lcout => OPEN,
            ltout => \ADC_IAC.n21159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_2_lut_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25011\,
            in3 => \N__24842\,
            lcout => \ADC_IAC.n21160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__29324\,
            in1 => \N__38405\,
            in2 => \N__26586\,
            in3 => \N__28961\,
            lcout => cmd_rdadctmp_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i19_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38449\,
            in1 => \N__26383\,
            in2 => \N__38265\,
            in3 => \N__29334\,
            lcout => cmd_rdadctmp_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i1_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24998\,
            in1 => \N__29333\,
            in2 => \N__24954\,
            in3 => \N__38453\,
            lcout => cmd_rdadctmp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i2_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38451\,
            in1 => \N__24999\,
            in2 => \N__24990\,
            in3 => \N__29336\,
            lcout => cmd_rdadctmp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__24950\,
            in1 => \N__29332\,
            in2 => \N__24975\,
            in3 => \N__38452\,
            lcout => cmd_rdadctmp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i20_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38450\,
            in1 => \N__26384\,
            in2 => \N__29429\,
            in3 => \N__29335\,
            lcout => cmd_rdadctmp_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.SCLK_35_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__38588\,
            in1 => \N__24941\,
            in2 => \N__24776\,
            in3 => \N__24855\,
            lcout => \IAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i17_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38762\,
            in1 => \N__38589\,
            in2 => \N__28887\,
            in3 => \N__24742\,
            lcout => buf_adcdata_iac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i16_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51489\,
            in1 => \N__31625\,
            in2 => \N__25799\,
            in3 => \N__25107\,
            lcout => buf_adcdata_vdc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42429\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7791_3_lut_4_lut_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001011011010"
        )
    port map (
            in0 => \N__51908\,
            in1 => \N__51174\,
            in2 => \N__52004\,
            in3 => \N__31661\,
            lcout => OPEN,
            ltout => \ADC_VDC.n10309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_adj_29_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111110"
        )
    port map (
            in0 => \N__51637\,
            in1 => \N__51488\,
            in2 => \N__25089\,
            in3 => \N__29688\,
            lcout => \ADC_VDC.n13276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001100000110000"
        )
    port map (
            in0 => \N__51894\,
            in1 => \N__51500\,
            in2 => \N__51709\,
            in3 => \N__51179\,
            lcout => adc_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42399\,
            ce => \N__25086\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i22_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51696\,
            in1 => \N__29080\,
            in2 => \N__30274\,
            in3 => \N__25530\,
            lcout => cmd_rdadctmp_22_adj_1501,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i10_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__25213\,
            in1 => \N__29070\,
            in2 => \N__25193\,
            in3 => \N__51602\,
            lcout => cmd_rdadctmp_10_adj_1513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__25046\,
            in1 => \N__51698\,
            in2 => \N__29114\,
            in3 => \N__25027\,
            lcout => cmd_rdadctmp_3_adj_1520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51697\,
            in1 => \N__25045\,
            in2 => \N__25073\,
            in3 => \N__29081\,
            lcout => cmd_rdadctmp_2_adj_1521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i4_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51600\,
            in1 => \N__25316\,
            in2 => \N__29115\,
            in3 => \N__25028\,
            lcout => cmd_rdadctmp_4_adj_1519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010001000"
        )
    port map (
            in0 => \N__51412\,
            in1 => \N__51599\,
            in2 => \N__51910\,
            in3 => \N__51145\,
            lcout => \ADC_VDC.n13463\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51601\,
            in1 => \N__25300\,
            in2 => \N__29116\,
            in3 => \N__25317\,
            lcout => cmd_rdadctmp_5_adj_1518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i8_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51704\,
            in1 => \N__25234\,
            in2 => \N__25281\,
            in3 => \N__29136\,
            lcout => cmd_rdadctmp_8_adj_1515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51701\,
            in1 => \N__25549\,
            in2 => \N__29142\,
            in3 => \N__25259\,
            lcout => cmd_rdadctmp_20_adj_1503,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51705\,
            in1 => \N__25214\,
            in2 => \N__25239\,
            in3 => \N__29137\,
            lcout => cmd_rdadctmp_9_adj_1514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51699\,
            in1 => \N__25165\,
            in2 => \N__29139\,
            in3 => \N__25189\,
            lcout => cmd_rdadctmp_11_adj_1512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51703\,
            in1 => \N__25487\,
            in2 => \N__25134\,
            in3 => \N__29135\,
            lcout => cmd_rdadctmp_14_adj_1509,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51700\,
            in1 => \N__25149\,
            in2 => \N__29140\,
            in3 => \N__25166\,
            lcout => cmd_rdadctmp_12_adj_1511,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__25148\,
            in1 => \N__51702\,
            in2 => \N__25133\,
            in3 => \N__29134\,
            lcout => cmd_rdadctmp_13_adj_1510,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__25486\,
            in1 => \N__51706\,
            in2 => \N__29141\,
            in3 => \N__25468\,
            lcout => cmd_rdadctmp_15_adj_1508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42424\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7_4_lut_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__26975\,
            in1 => \N__26516\,
            in2 => \N__26631\,
            in3 => \N__26957\,
            lcout => \ADC_VDC.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i9_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__25449\,
            in1 => \N__51475\,
            in2 => \N__31624\,
            in3 => \N__25430\,
            lcout => buf_adcdata_vdc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i6_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51473\,
            in1 => \N__31610\,
            in2 => \N__25397\,
            in3 => \N__25418\,
            lcout => buf_adcdata_vdc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31609\,
            in1 => \N__51474\,
            in2 => \N__27293\,
            in3 => \N__25380\,
            lcout => buf_adcdata_vdc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22473_bdd_4_lut_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000010"
        )
    port map (
            in0 => \N__25970\,
            in1 => \N__25896\,
            in2 => \N__46469\,
            in3 => \N__29589\,
            lcout => n22476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i16_3_lut_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25368\,
            in1 => \N__33027\,
            in2 => \_gnd_net_\,
            in3 => \N__57105\,
            lcout => n16_adj_1628,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i12698_2_lut_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__51690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26900\,
            lcout => \ADC_VDC.n15175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i10_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31580\,
            in1 => \N__51496\,
            in2 => \N__27350\,
            in3 => \N__25344\,
            lcout => buf_adcdata_vdc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i22_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__25332\,
            in1 => \N__51498\,
            in2 => \N__25676\,
            in3 => \N__31585\,
            lcout => buf_adcdata_vdc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51494\,
            in1 => \N__31583\,
            in2 => \N__25643\,
            in3 => \N__25659\,
            lcout => buf_adcdata_vdc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__51497\,
            in2 => \N__25604\,
            in3 => \N__25620\,
            lcout => buf_adcdata_vdc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__51495\,
            in1 => \N__25587\,
            in2 => \N__25571\,
            in3 => \N__31584\,
            lcout => buf_adcdata_vdc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i23_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31581\,
            in1 => \N__51499\,
            in2 => \N__27138\,
            in3 => \N__25863\,
            lcout => buf_adcdata_vdc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i21_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51746\,
            in1 => \N__25525\,
            in2 => \N__29138\,
            in3 => \N__25553\,
            lcout => cmd_rdadctmp_21_adj_1502,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i34_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__51478\,
            in1 => \N__25506\,
            in2 => \N__25842\,
            in3 => \N__51744\,
            lcout => cmd_rdadcbuf_34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42430\,
            ce => \N__25833\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i9_4_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26649\,
            in1 => \N__26610\,
            in2 => \N__26673\,
            in3 => \N__26694\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i11_3_lut_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25500\,
            in2 => \N__25491\,
            in3 => \N__30159\,
            lcout => \ADC_VDC.n18780\,
            ltout => \ADC_VDC.n18780_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25862\,
            in2 => \N__25845\,
            in3 => \N__51212\,
            lcout => \ADC_VDC.n4_adj_1451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011110000"
        )
    port map (
            in0 => \N__51211\,
            in1 => \N__51477\,
            in2 => \N__51759\,
            in3 => \N__51911\,
            lcout => \ADC_VDC.n13503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19823_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__46301\,
            in1 => \N__25824\,
            in2 => \N__56960\,
            in3 => \N__25715\,
            lcout => OPEN,
            ltout => \n22575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22575_bdd_4_lut_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__25806\,
            in1 => \N__25778\,
            in2 => \N__25743\,
            in3 => \N__46302\,
            lcout => n22578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40448\,
            in1 => \N__39639\,
            in2 => \_gnd_net_\,
            in3 => \N__25716\,
            lcout => \buf_cfgRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__47450\,
            in1 => \N__56787\,
            in2 => \_gnd_net_\,
            in3 => \N__46300\,
            lcout => OPEN,
            ltout => \n10902_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_279_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__49383\,
            in1 => \N__30477\,
            in2 => \N__25692\,
            in3 => \N__55430\,
            lcout => n12624,
            ltout => \n12624_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__25928\,
            in1 => \N__45348\,
            in2 => \N__25689\,
            in3 => \N__49384\,
            lcout => \buf_cfgRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55964\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i36_4_lut_4_lut_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001011001110"
        )
    port map (
            in0 => \N__46299\,
            in1 => \N__47165\,
            in2 => \N__56959\,
            in3 => \N__47449\,
            lcout => n30_adj_1499,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19809_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__25927\,
            in1 => \N__56783\,
            in2 => \N__25914\,
            in3 => \N__46298\,
            lcout => n22473,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_idxvec_i0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__43206\,
            in1 => \N__55402\,
            in2 => \N__43865\,
            in3 => \N__25887\,
            lcout => data_idxvec_0,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => n19813,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36170\,
            in1 => \N__44213\,
            in2 => \N__55465\,
            in3 => \N__25884\,
            lcout => data_idxvec_1,
            ltout => OPEN,
            carryin => n19813,
            carryout => n19814,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__34859\,
            in1 => \N__55406\,
            in2 => \N__35423\,
            in3 => \N__25881\,
            lcout => data_idxvec_2,
            ltout => OPEN,
            carryin => n19814,
            carryout => n19815,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i3_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__36486\,
            in1 => \N__41237\,
            in2 => \N__55466\,
            in3 => \N__25878\,
            lcout => data_idxvec_3,
            ltout => OPEN,
            carryin => n19815,
            carryout => n19816,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i4_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__36198\,
            in1 => \N__55410\,
            in2 => \N__30677\,
            in3 => \N__25875\,
            lcout => data_idxvec_4,
            ltout => OPEN,
            carryin => n19816,
            carryout => n19817,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i5_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37249\,
            in1 => \N__32327\,
            in2 => \N__55467\,
            in3 => \N__25872\,
            lcout => data_idxvec_5,
            ltout => OPEN,
            carryin => n19817,
            carryout => n19818,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i6_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__31727\,
            in1 => \N__55414\,
            in2 => \N__43457\,
            in3 => \N__25869\,
            lcout => data_idxvec_6,
            ltout => OPEN,
            carryin => n19818,
            carryout => n19819,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i7_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__32274\,
            in1 => \N__46544\,
            in2 => \N__55468\,
            in3 => \N__25866\,
            lcout => data_idxvec_7,
            ltout => OPEN,
            carryin => n19819,
            carryout => n19820,
            clk => \N__55975\,
            ce => \N__26156\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i8_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__40452\,
            in1 => \N__55420\,
            in2 => \N__40925\,
            in3 => \N__26034\,
            lcout => data_idxvec_8,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => n19821,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i9_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37452\,
            in1 => \N__55427\,
            in2 => \N__43106\,
            in3 => \N__26031\,
            lcout => data_idxvec_9,
            ltout => OPEN,
            carryin => n19821,
            carryout => n19822,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i10_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__32042\,
            in1 => \N__55421\,
            in2 => \N__40703\,
            in3 => \N__26028\,
            lcout => data_idxvec_10,
            ltout => OPEN,
            carryin => n19822,
            carryout => n19823,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i11_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__35253\,
            in1 => \N__55428\,
            in2 => \N__26061\,
            in3 => \N__26025\,
            lcout => data_idxvec_11,
            ltout => OPEN,
            carryin => n19823,
            carryout => n19824,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i12_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37206\,
            in1 => \N__55422\,
            in2 => \N__40379\,
            in3 => \N__26022\,
            lcout => data_idxvec_12,
            ltout => OPEN,
            carryin => n19824,
            carryout => n19825,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i13_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__30721\,
            in1 => \N__55429\,
            in2 => \N__32411\,
            in3 => \N__26019\,
            lcout => data_idxvec_13,
            ltout => OPEN,
            carryin => n19825,
            carryout => n19826,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i14_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__30359\,
            in1 => \N__55423\,
            in2 => \N__32600\,
            in3 => \N__26016\,
            lcout => data_idxvec_14,
            ltout => OPEN,
            carryin => n19826,
            carryout => n19827,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i15_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__28481\,
            in2 => \N__55469\,
            in3 => \N__26013\,
            lcout => data_idxvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55989\,
            ce => \N__26160\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i19_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27999\,
            in1 => \N__27839\,
            in2 => \N__26010\,
            in3 => \N__25969\,
            lcout => buf_adcdata_vac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_295_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110111"
        )
    port map (
            in0 => \N__55419\,
            in1 => \N__41124\,
            in2 => \N__49389\,
            in3 => \N__38946\,
            lcout => n12493,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15461_2_lut_3_lut_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__54863\,
            in1 => \N__49567\,
            in2 => \_gnd_net_\,
            in3 => \N__54573\,
            lcout => n14_adj_1571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22509_bdd_4_lut_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__26139\,
            in1 => \N__47536\,
            in2 => \N__32538\,
            in3 => \N__26040\,
            lcout => n22512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i7_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__49568\,
            in1 => \N__30806\,
            in2 => \N__49390\,
            in3 => \N__39515\,
            lcout => \VAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i19_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__28265\,
            in1 => \N__27445\,
            in2 => \N__26127\,
            in3 => \N__27840\,
            lcout => cmd_rdadctmp_19_adj_1473,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i2_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49365\,
            in1 => \N__39514\,
            in2 => \N__53458\,
            in3 => \N__26080\,
            lcout => \IAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15228_2_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28839\,
            in2 => \_gnd_net_\,
            in3 => \N__28801\,
            lcout => n17728,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__26264\,
            in1 => \N__46889\,
            in2 => \N__45480\,
            in3 => \N__46766\,
            lcout => buf_dds1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_3_i26_3_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56913\,
            in1 => \N__26060\,
            in2 => \_gnd_net_\,
            in3 => \N__37955\,
            lcout => OPEN,
            ltout => \n26_adj_1678_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19760_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__45753\,
            in1 => \N__47563\,
            in2 => \N__26043\,
            in3 => \N__46317\,
            lcout => n22509,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__31448\,
            in2 => \_gnd_net_\,
            in3 => \N__41666\,
            lcout => buf_dds0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56019\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i16_3_lut_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56914\,
            in1 => \N__26263\,
            in2 => \_gnd_net_\,
            in3 => \N__31447\,
            lcout => n16_adj_1645,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18607_3_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26418\,
            in1 => \N__47564\,
            in2 => \_gnd_net_\,
            in3 => \N__26250\,
            lcout => n21334,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27981\,
            in1 => \N__27833\,
            in2 => \N__43741\,
            in3 => \N__26238\,
            lcout => buf_adcdata_vac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i25_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__28240\,
            in1 => \N__26174\,
            in2 => \N__27856\,
            in3 => \N__26194\,
            lcout => cmd_rdadctmp_25_adj_1467,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i23_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__26323\,
            in1 => \N__27834\,
            in2 => \N__26354\,
            in3 => \N__28238\,
            lcout => cmd_rdadctmp_23_adj_1469,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_327_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45870\,
            in1 => \N__28046\,
            in2 => \_gnd_net_\,
            in3 => \N__35706\,
            lcout => acadc_rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i24_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__26173\,
            in1 => \N__27835\,
            in2 => \N__26328\,
            in3 => \N__28239\,
            lcout => cmd_rdadctmp_24_adj_1468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i9_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49369\,
            in1 => \N__31252\,
            in2 => \N__53462\,
            in3 => \N__41663\,
            lcout => buf_dds0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i14_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27979\,
            in1 => \N__27832\,
            in2 => \N__26355\,
            in3 => \N__32461\,
            lcout => buf_adcdata_vac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i15_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27831\,
            in1 => \N__27980\,
            in2 => \N__28432\,
            in3 => \N__26327\,
            lcout => buf_adcdata_vac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_293_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001000"
        )
    port map (
            in0 => \N__26313\,
            in1 => \N__55464\,
            in2 => \N__49370\,
            in3 => \N__44114\,
            lcout => n12654,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i11_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__26441\,
            in1 => \N__46885\,
            in2 => \N__45357\,
            in3 => \N__46732\,
            lcout => buf_dds1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i16_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__33796\,
            in1 => \N__29385\,
            in2 => \N__26300\,
            in3 => \N__38553\,
            lcout => cmd_rdadctmp_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i6_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__27373\,
            in1 => \N__49305\,
            in2 => \N__52290\,
            in3 => \N__39538\,
            lcout => \VAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i10_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49304\,
            in1 => \N__41664\,
            in2 => \N__45879\,
            in3 => \N__31081\,
            lcout => buf_dds0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i19_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__38500\,
            in1 => \N__26409\,
            in2 => \N__38770\,
            in3 => \N__26461\,
            lcout => buf_adcdata_iac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i17_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__38501\,
            in1 => \N__33803\,
            in2 => \N__33776\,
            in3 => \N__29382\,
            lcout => cmd_rdadctmp_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i4_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__26486\,
            in1 => \N__45352\,
            in2 => \N__49391\,
            in3 => \N__39539\,
            lcout => \IAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_start_329_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45648\,
            in1 => \N__28050\,
            in2 => \_gnd_net_\,
            in3 => \N__31028\,
            lcout => eis_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19842_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__26485\,
            in1 => \N__57097\,
            in2 => \N__26465\,
            in3 => \N__46406\,
            lcout => OPEN,
            ltout => \n22605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22605_bdd_4_lut_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__46407\,
            in1 => \N__31366\,
            in2 => \N__26445\,
            in3 => \N__26431\,
            lcout => n22608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i18_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__29381\,
            in1 => \N__38502\,
            in2 => \N__38264\,
            in3 => \N__33772\,
            lcout => cmd_rdadctmp_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56063\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i27_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38583\,
            in1 => \N__26401\,
            in2 => \N__32786\,
            in3 => \N__29372\,
            lcout => cmd_rdadctmp_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i11_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__38742\,
            in1 => \N__26385\,
            in2 => \N__41296\,
            in3 => \N__38584\,
            lcout => buf_adcdata_iac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__28879\,
            in1 => \N__29373\,
            in2 => \N__26370\,
            in3 => \N__38586\,
            lcout => cmd_rdadctmp_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i16_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38582\,
            in1 => \N__38743\,
            in2 => \N__39142\,
            in3 => \N__26369\,
            lcout => buf_adcdata_iac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i24_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__26365\,
            in1 => \N__38585\,
            in2 => \N__29390\,
            in3 => \N__28745\,
            lcout => cmd_rdadctmp_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i31_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__29213\,
            in1 => \N__38587\,
            in2 => \N__29391\,
            in3 => \N__26584\,
            lcout => cmd_rdadctmp_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56077\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16257_3_lut_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101100110"
        )
    port map (
            in0 => \N__51154\,
            in1 => \N__51882\,
            in2 => \_gnd_net_\,
            in3 => \N__26565\,
            lcout => OPEN,
            ltout => \ADC_VDC.n18783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i1_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51329\,
            in1 => \N__51636\,
            in2 => \N__26553\,
            in3 => \N__29148\,
            lcout => \ADC_VDC.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42398\,
            ce => \N__26550\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19425_4_lut_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011011111"
        )
    port map (
            in0 => \N__51635\,
            in1 => \N__51328\,
            in2 => \N__31398\,
            in3 => \N__26544\,
            lcout => \ADC_VDC.n16_adj_1450\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i39_3_lut_4_lut_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000110011"
        )
    port map (
            in0 => \N__51153\,
            in1 => \N__51975\,
            in2 => \N__31662\,
            in3 => \N__51881\,
            lcout => \ADC_VDC.n18\,
            ltout => \ADC_VDC.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19428_4_lut_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111101111"
        )
    port map (
            in0 => \N__51327\,
            in1 => \N__51634\,
            in2 => \N__26538\,
            in3 => \N__29687\,
            lcout => \ADC_VDC.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18466_2_lut_3_lut_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__51152\,
            in1 => \N__51974\,
            in2 => \_gnd_net_\,
            in3 => \N__51880\,
            lcout => \ADC_VDC.n21193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i7_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26535\,
            lcout => buf_control_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55940\,
            ce => \N__42069\,
            sr => \N__42093\
        );

    \ADC_VDC.avg_cnt_i0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26517\,
            in2 => \_gnd_net_\,
            in3 => \N__26505\,
            lcout => \ADC_VDC.avg_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \ADC_VDC.n19877\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26690\,
            in2 => \_gnd_net_\,
            in3 => \N__26676\,
            lcout => \ADC_VDC.avg_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19877\,
            carryout => \ADC_VDC.n19878\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26669\,
            in2 => \_gnd_net_\,
            in3 => \N__26655\,
            lcout => \ADC_VDC.avg_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19878\,
            carryout => \ADC_VDC.n19879\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30171\,
            in2 => \_gnd_net_\,
            in3 => \N__26652\,
            lcout => \ADC_VDC.avg_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19879\,
            carryout => \ADC_VDC.n19880\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26648\,
            in2 => \_gnd_net_\,
            in3 => \N__26634\,
            lcout => \ADC_VDC.avg_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19880\,
            carryout => \ADC_VDC.n19881\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26630\,
            in2 => \_gnd_net_\,
            in3 => \N__26616\,
            lcout => \ADC_VDC.avg_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19881\,
            carryout => \ADC_VDC.n19882\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30185\,
            in2 => \_gnd_net_\,
            in3 => \N__26613\,
            lcout => \ADC_VDC.avg_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19882\,
            carryout => \ADC_VDC.n19883\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i7_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26609\,
            in2 => \_gnd_net_\,
            in3 => \N__26595\,
            lcout => \ADC_VDC.avg_cnt_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19883\,
            carryout => \ADC_VDC.n19884\,
            clk => \N__42362\,
            ce => \N__26940\,
            sr => \N__26864\
        );

    \ADC_VDC.avg_cnt_i8_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30198\,
            in2 => \_gnd_net_\,
            in3 => \N__26592\,
            lcout => \ADC_VDC.avg_cnt_8\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \ADC_VDC.n19885\,
            clk => \N__42409\,
            ce => \N__26929\,
            sr => \N__26863\
        );

    \ADC_VDC.avg_cnt_i9_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30210\,
            in2 => \_gnd_net_\,
            in3 => \N__26589\,
            lcout => \ADC_VDC.avg_cnt_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19885\,
            carryout => \ADC_VDC.n19886\,
            clk => \N__42409\,
            ce => \N__26929\,
            sr => \N__26863\
        );

    \ADC_VDC.avg_cnt_i10_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26976\,
            in2 => \_gnd_net_\,
            in3 => \N__26964\,
            lcout => \ADC_VDC.avg_cnt_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19886\,
            carryout => \ADC_VDC.n19887\,
            clk => \N__42409\,
            ce => \N__26929\,
            sr => \N__26863\
        );

    \ADC_VDC.avg_cnt_i11_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26958\,
            in2 => \_gnd_net_\,
            in3 => \N__26961\,
            lcout => \ADC_VDC.avg_cnt_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42409\,
            ce => \N__26929\,
            sr => \N__26863\
        );

    \ADC_VDC.ADC_DATA_i12_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31587\,
            in1 => \N__51483\,
            in2 => \N__28019\,
            in3 => \N__26796\,
            lcout => buf_adcdata_vdc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i7_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__26781\,
            in1 => \N__26759\,
            in2 => \N__51501\,
            in3 => \N__31589\,
            lcout => buf_adcdata_vdc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i23_3_lut_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57185\,
            in1 => \N__35996\,
            in2 => \_gnd_net_\,
            in3 => \N__33048\,
            lcout => n23_adj_1668,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_35_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__51480\,
            in1 => \N__51745\,
            in2 => \N__51915\,
            in3 => \N__51197\,
            lcout => n11891,
            ltout => \n11891_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i15_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__28403\,
            in1 => \N__51484\,
            in2 => \N__26748\,
            in3 => \N__26745\,
            lcout => buf_adcdata_vdc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i14_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51481\,
            in1 => \N__31588\,
            in2 => \N__32489\,
            in3 => \N__26727\,
            lcout => buf_adcdata_vdc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i11_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31586\,
            in1 => \N__51482\,
            in2 => \N__35069\,
            in3 => \N__26709\,
            lcout => buf_adcdata_vdc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i23_3_lut_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27198\,
            in1 => \N__56957\,
            in2 => \_gnd_net_\,
            in3 => \N__31184\,
            lcout => n23_adj_1658,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.SCLK_27_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000110001"
        )
    port map (
            in0 => \N__29840\,
            in1 => \N__30093\,
            in2 => \N__27179\,
            in3 => \N__29951\,
            lcout => \DDS_SCK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19833_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__27014\,
            in1 => \N__56958\,
            in2 => \N__27162\,
            in3 => \N__46308\,
            lcout => OPEN,
            ltout => \n22593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22593_bdd_4_lut_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__46309\,
            in1 => \N__27137\,
            in2 => \N__27123\,
            in3 => \N__27113\,
            lcout => n21240,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i6_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49377\,
            in1 => \N__39641\,
            in2 => \N__49569\,
            in3 => \N__27053\,
            lcout => \buf_cfgRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i7_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__27015\,
            in1 => \N__49378\,
            in2 => \N__42554\,
            in3 => \N__39642\,
            lcout => \buf_cfgRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55952\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_60_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__46307\,
            in1 => \N__37589\,
            in2 => \N__26985\,
            in3 => \N__47702\,
            lcout => \comm_state_3_N_460_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_59_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56867\,
            in2 => \_gnd_net_\,
            in3 => \N__46306\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i13_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__27998\,
            in1 => \N__27842\,
            in2 => \N__28313\,
            in3 => \N__28088\,
            lcout => buf_adcdata_vac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_307_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47164\,
            in2 => \_gnd_net_\,
            in3 => \N__32390\,
            lcout => n4_adj_1455,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i11_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__27841\,
            in1 => \N__27997\,
            in2 => \N__27465\,
            in3 => \N__35044\,
            lcout => buf_adcdata_vac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i4_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49385\,
            in1 => \N__39640\,
            in2 => \N__34999\,
            in3 => \N__47799\,
            lcout => \buf_cfgRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i19_3_lut_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29508\,
            in1 => \N__27425\,
            in2 => \_gnd_net_\,
            in3 => \N__56868\,
            lcout => n19_adj_1666,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i17_3_lut_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56869\,
            in1 => \N__28940\,
            in2 => \_gnd_net_\,
            in3 => \N__27383\,
            lcout => n17_adj_1665,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i19_3_lut_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27354\,
            in1 => \N__27329\,
            in2 => \_gnd_net_\,
            in3 => \N__57026\,
            lcout => n19_adj_1646,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i19_3_lut_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57025\,
            in1 => \N__27294\,
            in2 => \_gnd_net_\,
            in3 => \N__27272\,
            lcout => OPEN,
            ltout => \n19_adj_1534_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i22_3_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27230\,
            in2 => \N__27201\,
            in3 => \N__47519\,
            lcout => n22_adj_1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i0_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__57028\,
            in1 => \N__48696\,
            in2 => \N__50980\,
            in3 => \N__37531\,
            lcout => comm_cmd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55965\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19701_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__28359\,
            in1 => \N__46310\,
            in2 => \N__28347\,
            in3 => \N__47518\,
            lcout => n22431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i19_3_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57027\,
            in1 => \N__28312\,
            in2 => \_gnd_net_\,
            in3 => \N__29631\,
            lcout => OPEN,
            ltout => \n19_adj_1629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19653_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__28287\,
            in1 => \N__46311\,
            in2 => \N__28272\,
            in3 => \N__47520\,
            lcout => n22365,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_261_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__31154\,
            in1 => \N__55418\,
            in2 => \N__28062\,
            in3 => \N__54008\,
            lcout => n10695,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i21_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__27843\,
            in1 => \N__28078\,
            in2 => \N__27513\,
            in3 => \N__28266\,
            lcout => cmd_rdadctmp_21_adj_1471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_368_i8_2_lut_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46291\,
            in2 => \_gnd_net_\,
            in3 => \N__47601\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_stop_328_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__53448\,
            in1 => \N__28034\,
            in2 => \_gnd_net_\,
            in3 => \N__43028\,
            lcout => eis_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i19_3_lut_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28023\,
            in1 => \N__27481\,
            in2 => \_gnd_net_\,
            in3 => \N__56873\,
            lcout => n19_adj_1634,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i12_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__28000\,
            in1 => \N__27482\,
            in2 => \N__27857\,
            in3 => \N__27512\,
            lcout => buf_adcdata_vac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i12_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__36277\,
            in1 => \N__46898\,
            in2 => \N__47819\,
            in3 => \N__46746\,
            lcout => buf_dds1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19658_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__46369\,
            in1 => \N__28994\,
            in2 => \N__29202\,
            in3 => \N__56899\,
            lcout => n22371,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_4_lut_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30963\,
            in1 => \N__35709\,
            in2 => \N__28665\,
            in3 => \N__37771\,
            lcout => \iac_raw_buf_N_774\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1564638_i1_3_lut_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47245\,
            in1 => \N__28494\,
            in2 => \_gnd_net_\,
            in3 => \N__28488\,
            lcout => n30_adj_1679,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i26_3_lut_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28482\,
            in1 => \N__57205\,
            in2 => \_gnd_net_\,
            in3 => \N__28643\,
            lcout => OPEN,
            ltout => \n26_adj_1659_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18597_4_lut_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__46371\,
            in1 => \N__28467\,
            in2 => \N__28446\,
            in3 => \N__56900\,
            lcout => OPEN,
            ltout => \n21324_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19799_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__28365\,
            in1 => \N__47244\,
            in2 => \N__28443\,
            in3 => \N__47703\,
            lcout => n22401,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i19_3_lut_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28433\,
            in1 => \N__28407\,
            in2 => \_gnd_net_\,
            in3 => \N__56898\,
            lcout => n19_adj_1621,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18596_4_lut_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__34494\,
            in1 => \N__57204\,
            in2 => \N__28377\,
            in3 => \N__46370\,
            lcout => n21323,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22371_bdd_4_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__30889\,
            in1 => \N__28722\,
            in2 => \N__31299\,
            in3 => \N__46318\,
            lcout => n22374,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18_3_lut_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35874\,
            in1 => \N__35776\,
            in2 => \_gnd_net_\,
            in3 => \N__30968\,
            lcout => OPEN,
            ltout => \n12_adj_1454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_trig_300_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000100"
        )
    port map (
            in0 => \N__35733\,
            in1 => \N__28664\,
            in2 => \N__28716\,
            in3 => \N__28697\,
            lcout => acadc_trig,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_300C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_209_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35859\,
            in2 => \_gnd_net_\,
            in3 => \N__35775\,
            lcout => n21053,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15227_2_lut_3_lut_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__30966\,
            in1 => \N__28848\,
            in2 => \_gnd_net_\,
            in3 => \N__28806\,
            lcout => \eis_state_2_N_392_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_269_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35873\,
            in1 => \N__28862\,
            in2 => \_gnd_net_\,
            in3 => \N__30908\,
            lcout => OPEN,
            ltout => \n21042_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_286_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111110011"
        )
    port map (
            in0 => \N__30967\,
            in1 => \N__35800\,
            in2 => \N__28650\,
            in3 => \N__35875\,
            lcout => OPEN,
            ltout => \n21030_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_299_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__28644\,
            in1 => \N__35734\,
            in2 => \N__28647\,
            in3 => \N__35777\,
            lcout => eis_end,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_300C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_1__bdd_4_lut_19731_4_lut_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111000101010"
        )
    port map (
            in0 => \N__35866\,
            in1 => \N__35783\,
            in2 => \N__30981\,
            in3 => \N__28764\,
            lcout => n22437,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19465_3_lut_4_lut_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__35860\,
            in1 => \N__30955\,
            in2 => \N__35794\,
            in3 => \N__35707\,
            lcout => n11989,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__31029\,
            in1 => \N__43043\,
            in2 => \N__30980\,
            in3 => \N__28863\,
            lcout => OPEN,
            ltout => \n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19423_3_lut_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__35782\,
            in1 => \_gnd_net_\,
            in2 => \N__28851\,
            in3 => \N__35865\,
            lcout => n11908,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_adj_270_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__35708\,
            in1 => \N__30964\,
            in2 => \N__35876\,
            in3 => \N__35781\,
            lcout => n11933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15247_2_lut_3_lut_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__35861\,
            in1 => \N__28847\,
            in2 => \_gnd_net_\,
            in3 => \N__28802\,
            lcout => \eis_state_2_N_392_1\,
            ltout => \eis_state_2_N_392_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_2__I_0_371_Mux_1_i2_4_lut_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__31030\,
            in1 => \N__30965\,
            in2 => \N__28758\,
            in3 => \N__32815\,
            lcout => OPEN,
            ltout => \n2_adj_1696_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i1_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__35784\,
            in1 => \N__30962\,
            in2 => \N__28755\,
            in3 => \N__28752\,
            lcout => eis_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i1C_net\,
            ce => \N__30995\,
            sr => \N__35735\
        );

    \ADC_IAC.ADC_DATA_i15_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38737\,
            in1 => \N__38551\,
            in2 => \N__42046\,
            in3 => \N__28746\,
            lcout => buf_adcdata_iac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i9_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49302\,
            in1 => \N__47863\,
            in2 => \N__53466\,
            in3 => \N__42977\,
            lcout => \acadc_skipCount_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i12_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49303\,
            in1 => \N__36256\,
            in2 => \N__47820\,
            in3 => \N__41665\,
            lcout => buf_dds0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i8_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__42543\,
            in1 => \N__39516\,
            in2 => \N__49382\,
            in3 => \N__28990\,
            lcout => \VAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i15_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49301\,
            in1 => \N__47862\,
            in2 => \N__31185\,
            in3 => \N__42542\,
            lcout => \acadc_skipCount_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i21_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38738\,
            in1 => \N__38552\,
            in2 => \N__28971\,
            in3 => \N__28933\,
            lcout => buf_adcdata_iac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i20_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38746\,
            in1 => \N__38504\,
            in2 => \N__28911\,
            in3 => \N__32128\,
            lcout => buf_adcdata_iac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i3_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49337\,
            in1 => \N__39528\,
            in2 => \N__45878\,
            in3 => \N__30526\,
            lcout => \IAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i12_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38503\,
            in1 => \N__38745\,
            in2 => \N__29430\,
            in3 => \N__30601\,
            lcout => buf_adcdata_iac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i11_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49336\,
            in1 => \N__31367\,
            in2 => \N__45356\,
            in3 => \N__41667\,
            lcout => buf_dds0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i8_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49335\,
            in1 => \N__47864\,
            in2 => \N__45646\,
            in3 => \N__32719\,
            lcout => \acadc_skipCount_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i26_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__29364\,
            in1 => \N__32779\,
            in2 => \N__28886\,
            in3 => \N__38597\,
            lcout => cmd_rdadctmp_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i21_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__38595\,
            in1 => \N__33097\,
            in2 => \N__29428\,
            in3 => \N__29365\,
            lcout => cmd_rdadctmp_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i23_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38744\,
            in1 => \N__38596\,
            in2 => \N__29217\,
            in3 => \N__29188\,
            lcout => buf_adcdata_iac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i2_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__51867\,
            in1 => \N__51344\,
            in2 => \_gnd_net_\,
            in3 => \N__51180\,
            lcout => adc_state_2_adj_1500,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42364\,
            ce => \N__29166\,
            sr => \N__31383\
        );

    \ADC_VDC.i19237_4_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__34374\,
            in1 => \N__34338\,
            in2 => \N__34440\,
            in3 => \N__34401\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19248_4_lut_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__51892\,
            in1 => \N__31680\,
            in2 => \N__29154\,
            in3 => \N__34305\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.n22587_bdd_4_lut_4_lut_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101010000"
        )
    port map (
            in0 => \N__51356\,
            in1 => \N__51893\,
            in2 => \N__29151\,
            in3 => \N__30291\,
            lcout => \ADC_VDC.n22590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_34_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__51151\,
            in1 => \N__51355\,
            in2 => \N__51909\,
            in3 => \N__51711\,
            lcout => n13324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i24_3_lut_4_lut_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110000"
        )
    port map (
            in0 => \N__51710\,
            in1 => \N__51149\,
            in2 => \N__51414\,
            in3 => \N__51986\,
            lcout => \ADC_VDC.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51357\,
            in2 => \_gnd_net_\,
            in3 => \N__51713\,
            lcout => \ADC_VDC.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16264_3_lut_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001100110"
        )
    port map (
            in0 => \N__51856\,
            in1 => \N__51985\,
            in2 => \_gnd_net_\,
            in3 => \N__51150\,
            lcout => OPEN,
            ltout => \ADC_VDC.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_32_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111110"
        )
    port map (
            in0 => \N__51442\,
            in1 => \N__51712\,
            in2 => \N__29691\,
            in3 => \N__29686\,
            lcout => \ADC_VDC.n65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i8_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__43769\,
            in1 => \N__31601\,
            in2 => \N__51491\,
            in3 => \N__29670\,
            lcout => buf_adcdata_vdc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i13_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51361\,
            in1 => \N__29621\,
            in2 => \N__31617\,
            in3 => \N__29649\,
            lcout => buf_adcdata_vdc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i19_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__29582\,
            in1 => \N__31600\,
            in2 => \N__51490\,
            in3 => \N__29610\,
            lcout => buf_adcdata_vdc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i17_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51362\,
            in1 => \N__29540\,
            in2 => \N__31618\,
            in3 => \N__29571\,
            lcout => buf_adcdata_vdc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i21_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__29529\,
            in1 => \N__31590\,
            in2 => \N__29501\,
            in3 => \N__51364\,
            lcout => buf_adcdata_vdc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i20_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__51363\,
            in1 => \N__31895\,
            in2 => \N__31619\,
            in3 => \N__29484\,
            lcout => buf_adcdata_vdc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i16_3_lut_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29463\,
            in1 => \N__32255\,
            in2 => \_gnd_net_\,
            in3 => \N__57208\,
            lcout => n16_adj_1633,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110001101100"
        )
    port map (
            in0 => \N__51860\,
            in1 => \N__51175\,
            in2 => \N__51415\,
            in3 => \N__30285\,
            lcout => \ADC_VDC.n22587\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i3_4_lut_adj_30_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__34369\,
            in1 => \N__31470\,
            in2 => \N__34436\,
            in3 => \N__31671\,
            lcout => \ADC_VDC.n10708\,
            ltout => \ADC_VDC.n10708_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i23_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__30236\,
            in1 => \N__30278\,
            in2 => \N__30246\,
            in3 => \N__51203\,
            lcout => \ADC_VDC.cmd_rdadctmp_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42414\,
            ce => \N__31941\,
            sr => \N__30222\
        );

    \ADC_VDC.i8_4_lut_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30209\,
            in1 => \N__30197\,
            in2 => \N__30186\,
            in3 => \N__30170\,
            lcout => \ADC_VDC.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19393_4_lut_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100110"
        )
    port map (
            in0 => \N__30072\,
            in1 => \N__29947\,
            in2 => \N__38828\,
            in3 => \N__29792\,
            lcout => \CLK_DDS.n13005\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i23_4_lut_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000010101"
        )
    port map (
            in0 => \N__29794\,
            in1 => \N__38824\,
            in2 => \N__29952\,
            in3 => \N__30074\,
            lcout => \CLK_DDS.n9_adj_1433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19409_4_lut_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__30073\,
            in1 => \N__29946\,
            in2 => \N__38829\,
            in3 => \N__29793\,
            lcout => \CLK_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secclk_cnt_3765_3766__i1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34554\,
            in2 => \_gnd_net_\,
            in3 => \N__29694\,
            lcout => secclk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => n19956,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34610\,
            in2 => \_gnd_net_\,
            in3 => \N__30318\,
            lcout => secclk_cnt_1,
            ltout => OPEN,
            carryin => n19956,
            carryout => n19957,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31785\,
            in2 => \_gnd_net_\,
            in3 => \N__30315\,
            lcout => secclk_cnt_2,
            ltout => OPEN,
            carryin => n19957,
            carryout => n19958,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i4_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31803\,
            in2 => \_gnd_net_\,
            in3 => \N__30312\,
            lcout => secclk_cnt_3,
            ltout => OPEN,
            carryin => n19958,
            carryout => n19959,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34517\,
            in2 => \_gnd_net_\,
            in3 => \N__30309\,
            lcout => secclk_cnt_4,
            ltout => OPEN,
            carryin => n19959,
            carryout => n19960,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i6_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34592\,
            in2 => \_gnd_net_\,
            in3 => \N__30306\,
            lcout => secclk_cnt_5,
            ltout => OPEN,
            carryin => n19960,
            carryout => n19961,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i7_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31845\,
            in2 => \_gnd_net_\,
            in3 => \N__30303\,
            lcout => secclk_cnt_6,
            ltout => OPEN,
            carryin => n19961,
            carryout => n19962,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i8_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31760\,
            in2 => \_gnd_net_\,
            in3 => \N__30300\,
            lcout => secclk_cnt_7,
            ltout => OPEN,
            carryin => n19962,
            carryout => n19963,
            clk => \N__50782\,
            ce => 'H',
            sr => \N__34714\
        );

    \secclk_cnt_3765_3766__i9_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34625\,
            in2 => \_gnd_net_\,
            in3 => \N__30297\,
            lcout => secclk_cnt_8,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => n19964,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i10_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35144\,
            in2 => \_gnd_net_\,
            in3 => \N__30294\,
            lcout => secclk_cnt_9,
            ltout => OPEN,
            carryin => n19964,
            carryout => n19965,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i11_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31817\,
            in2 => \_gnd_net_\,
            in3 => \N__30345\,
            lcout => secclk_cnt_10,
            ltout => OPEN,
            carryin => n19965,
            carryout => n19966,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i12_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34532\,
            in2 => \_gnd_net_\,
            in3 => \N__30342\,
            lcout => secclk_cnt_11,
            ltout => OPEN,
            carryin => n19966,
            carryout => n19967,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i13_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30392\,
            in2 => \_gnd_net_\,
            in3 => \N__30339\,
            lcout => secclk_cnt_12,
            ltout => OPEN,
            carryin => n19967,
            carryout => n19968,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i14_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31773\,
            in2 => \_gnd_net_\,
            in3 => \N__30336\,
            lcout => secclk_cnt_13,
            ltout => OPEN,
            carryin => n19968,
            carryout => n19969,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i15_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31833\,
            in2 => \_gnd_net_\,
            in3 => \N__30333\,
            lcout => secclk_cnt_14,
            ltout => OPEN,
            carryin => n19969,
            carryout => n19970,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i16_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34643\,
            in2 => \_gnd_net_\,
            in3 => \N__30330\,
            lcout => secclk_cnt_15,
            ltout => OPEN,
            carryin => n19970,
            carryout => n19971,
            clk => \N__50786\,
            ce => 'H',
            sr => \N__34716\
        );

    \secclk_cnt_3765_3766__i17_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31746\,
            in2 => \_gnd_net_\,
            in3 => \N__30327\,
            lcout => secclk_cnt_16,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => n19972,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \secclk_cnt_3765_3766__i18_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35129\,
            in2 => \_gnd_net_\,
            in3 => \N__30324\,
            lcout => secclk_cnt_17,
            ltout => OPEN,
            carryin => n19972,
            carryout => n19973,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \secclk_cnt_3765_3766__i19_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34571\,
            in2 => \_gnd_net_\,
            in3 => \N__30321\,
            lcout => secclk_cnt_18,
            ltout => OPEN,
            carryin => n19973,
            carryout => n19974,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \secclk_cnt_3765_3766__i20_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30408\,
            in2 => \_gnd_net_\,
            in3 => \N__30435\,
            lcout => secclk_cnt_19,
            ltout => OPEN,
            carryin => n19974,
            carryout => n19975,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \secclk_cnt_3765_3766__i21_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31928\,
            in2 => \_gnd_net_\,
            in3 => \N__30432\,
            lcout => secclk_cnt_20,
            ltout => OPEN,
            carryin => n19975,
            carryout => n19976,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \secclk_cnt_3765_3766__i22_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30422\,
            in2 => \_gnd_net_\,
            in3 => \N__30429\,
            lcout => secclk_cnt_21,
            ltout => OPEN,
            carryin => n19976,
            carryout => n19977,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \secclk_cnt_3765_3766__i23_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30378\,
            in2 => \_gnd_net_\,
            in3 => \N__30426\,
            lcout => secclk_cnt_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50788\,
            ce => 'H',
            sr => \N__34715\
        );

    \i6_4_lut_adj_201_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30423\,
            in1 => \N__30407\,
            in2 => \N__30396\,
            in3 => \N__30377\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6751_2_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54500\,
            in2 => \_gnd_net_\,
            in3 => \N__54001\,
            lcout => n9269,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__49350\,
            in1 => \N__47923\,
            in2 => \N__32562\,
            in3 => \N__45335\,
            lcout => \acadc_skipCount_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i14_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__47924\,
            in1 => \N__49351\,
            in2 => \N__49586\,
            in3 => \N__32217\,
            lcout => \acadc_skipCount_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i8_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35561\,
            in1 => \N__40447\,
            in2 => \_gnd_net_\,
            in3 => \N__30841\,
            lcout => req_data_cnt_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31991\,
            in1 => \N__30366\,
            in2 => \_gnd_net_\,
            in3 => \N__35560\,
            lcout => req_data_cnt_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55953\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18602_4_lut_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__46455\,
            in1 => \N__56865\,
            in2 => \N__32226\,
            in3 => \N__31990\,
            lcout => n21329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i17_3_lut_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56866\,
            in1 => \N__32756\,
            in2 => \_gnd_net_\,
            in3 => \N__30542\,
            lcout => n17_adj_1682,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_310_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__56751\,
            in1 => \N__37572\,
            in2 => \_gnd_net_\,
            in3 => \N__47133\,
            lcout => n11570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22401_bdd_4_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__47136\,
            in1 => \N__30507\,
            in2 => \N__30498\,
            in3 => \N__30486\,
            lcout => n22404,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i15_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__42535\,
            in1 => \N__49325\,
            in2 => \N__31294\,
            in3 => \N__41668\,
            lcout => buf_dds0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_278_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__47134\,
            in1 => \_gnd_net_\,
            in2 => \N__37582\,
            in3 => \N__54007\,
            lcout => n21122,
            ltout => \n21122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_276_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__32637\,
            in1 => \N__49323\,
            in2 => \N__30465\,
            in3 => \N__55296\,
            lcout => n12610,
            ltout => \n12610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__49324\,
            in1 => \N__47787\,
            in2 => \N__30462\,
            in3 => \N__32090\,
            lcout => \VAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55957\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i30_3_lut_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30459\,
            in1 => \N__30444\,
            in2 => \_gnd_net_\,
            in3 => \N__47135\,
            lcout => n30_adj_1605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_53_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__37571\,
            in1 => \N__56752\,
            in2 => \_gnd_net_\,
            in3 => \N__54006\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i26_3_lut_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30678\,
            in1 => \N__56874\,
            in2 => \_gnd_net_\,
            in3 => \N__37695\,
            lcout => OPEN,
            ltout => \n26_adj_1635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19706_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__57318\,
            in1 => \N__46296\,
            in2 => \N__30651\,
            in3 => \N__47706\,
            lcout => OPEN,
            ltout => \n22443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22443_bdd_4_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47707\,
            in1 => \N__32667\,
            in2 => \N__30648\,
            in3 => \N__35335\,
            lcout => OPEN,
            ltout => \n22446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1569462_i1_3_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30564\,
            in2 => \N__30645\,
            in3 => \N__47269\,
            lcout => OPEN,
            ltout => \n30_adj_1636_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54571\,
            in1 => \_gnd_net_\,
            in2 => \N__30642\,
            in3 => \N__53644\,
            lcout => comm_buf_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55966\,
            ce => \N__45213\,
            sr => \N__44015\
        );

    \comm_cmd_1__bdd_4_lut_19736_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__30639\,
            in1 => \N__46295\,
            in2 => \N__30633\,
            in3 => \N__47704\,
            lcout => OPEN,
            ltout => \n22467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22467_bdd_4_lut_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__47705\,
            in1 => \N__30608\,
            in2 => \N__30579\,
            in3 => \N__30576\,
            lcout => n22470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19726_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__57203\,
            in1 => \N__46458\,
            in2 => \N__31045\,
            in3 => \N__30845\,
            lcout => OPEN,
            ltout => \n22395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22395_bdd_4_lut_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__46459\,
            in1 => \N__44791\,
            in2 => \N__30849\,
            in3 => \N__32727\,
            lcout => n22398,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_155_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__40905\,
            in1 => \N__37908\,
            in2 => \N__30846\,
            in3 => \N__34768\,
            lcout => n19_adj_1526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__46456\,
            in1 => \N__30805\,
            in2 => \N__30780\,
            in3 => \N__57202\,
            lcout => OPEN,
            ltout => \n22635_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22635_bdd_4_lut_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__31323\,
            in1 => \N__35630\,
            in2 => \N__30738\,
            in3 => \N__46457\,
            lcout => n21236,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i13_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__34769\,
            in1 => \_gnd_net_\,
            in2 => \N__30722\,
            in3 => \N__35570\,
            lcout => req_data_cnt_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55977\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35571\,
            in1 => \N__31728\,
            in2 => \_gnd_net_\,
            in3 => \N__43517\,
            lcout => req_data_cnt_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55977\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43199\,
            in1 => \N__35569\,
            in2 => \_gnd_net_\,
            in3 => \N__43648\,
            lcout => req_data_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55977\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_2__I_0_371_Mux_0_i2_4_lut_4_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111110111"
        )
    port map (
            in0 => \N__31047\,
            in1 => \N__32816\,
            in2 => \N__30984\,
            in3 => \N__37780\,
            lcout => OPEN,
            ltout => \n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i0_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000010001"
        )
    port map (
            in0 => \N__35792\,
            in1 => \N__30979\,
            in2 => \N__30681\,
            in3 => \N__31053\,
            lcout => eis_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30996\,
            sr => \N__35732\
        );

    \i19138_2_lut_4_lut_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__43042\,
            in1 => \N__32421\,
            in2 => \N__30982\,
            in3 => \N__32069\,
            lcout => OPEN,
            ltout => \n21501_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_1__bdd_4_lut_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__35791\,
            in1 => \N__35871\,
            in2 => \N__31062\,
            in3 => \N__31059\,
            lcout => n22479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i29_4_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100001101"
        )
    port map (
            in0 => \N__31046\,
            in1 => \N__32817\,
            in2 => \N__30983\,
            in3 => \N__37779\,
            lcout => OPEN,
            ltout => \n11_adj_1632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i2_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__35793\,
            in1 => \N__35872\,
            in2 => \N__30999\,
            in3 => \N__30909\,
            lcout => eis_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30996\,
            sr => \N__35732\
        );

    \i1_2_lut_4_lut_4_lut_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__30969\,
            in1 => \N__43041\,
            in2 => \N__32073\,
            in3 => \N__32420\,
            lcout => n21041,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i16_3_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57207\,
            in1 => \N__35603\,
            in2 => \_gnd_net_\,
            in3 => \N__31198\,
            lcout => n16_adj_1651,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i16_3_lut_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30862\,
            in1 => \N__31091\,
            in2 => \_gnd_net_\,
            in3 => \N__57206\,
            lcout => n16_adj_1681,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i15_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46755\,
            in1 => \N__42555\,
            in2 => \N__46899\,
            in3 => \N__30893\,
            lcout => buf_dds1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i10_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__30872\,
            in1 => \N__46874\,
            in2 => \N__45874\,
            in3 => \N__46756\,
            lcout => buf_dds1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_161_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__46453\,
            in1 => \N__47192\,
            in2 => \N__57261\,
            in3 => \N__47666\,
            lcout => n5_adj_1536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i6_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__36129\,
            in1 => \N__55433\,
            in2 => \N__49341\,
            in3 => \N__38033\,
            lcout => data_index_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31199\,
            in1 => \N__36171\,
            in2 => \_gnd_net_\,
            in3 => \N__41662\,
            lcout => buf_dds0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36780\,
            in1 => \N__31171\,
            in2 => \N__37065\,
            in3 => \N__42973\,
            lcout => n24_adj_1593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12382_2_lut_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__37808\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35870\,
            lcout => n14907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__46460\,
            in1 => \N__47665\,
            in2 => \N__31158\,
            in3 => \N__54009\,
            lcout => n8841,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \EIS_SYNCCLK_I_0_1_lut_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \IAC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i14_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49297\,
            in1 => \N__31318\,
            in2 => \N__49587\,
            in3 => \N__41658\,
            lcout => buf_dds0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56021\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i10_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44638\,
            in1 => \N__44492\,
            in2 => \N__31233\,
            in3 => \N__31092\,
            lcout => \SIG_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i11_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__44493\,
            in1 => \N__44642\,
            in2 => \N__31377\,
            in3 => \N__31368\,
            lcout => \SIG_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i12_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44639\,
            in1 => \N__44494\,
            in2 => \N__31350\,
            in3 => \N__36257\,
            lcout => \SIG_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i13_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__44495\,
            in1 => \N__44643\,
            in2 => \N__31341\,
            in3 => \N__35310\,
            lcout => \SIG_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i14_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44640\,
            in1 => \N__44496\,
            in2 => \N__31332\,
            in3 => \N__31319\,
            lcout => \SIG_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i15_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__44497\,
            in1 => \N__44644\,
            in2 => \N__31298\,
            in3 => \N__31263\,
            lcout => tmp_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i9_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44641\,
            in1 => \N__44499\,
            in2 => \N__31224\,
            in3 => \N__31257\,
            lcout => \SIG_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i8_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__44498\,
            in1 => \N__36621\,
            in2 => \N__39081\,
            in3 => \N__44645\,
            lcout => \SIG_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56035\,
            ce => \N__43910\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44646\,
            in1 => \N__44449\,
            in2 => \N__39005\,
            in3 => \N__41538\,
            lcout => \SIG_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__44450\,
            in1 => \N__44650\,
            in2 => \N__31212\,
            in3 => \N__31203\,
            lcout => \SIG_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i2_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44647\,
            in1 => \N__44451\,
            in2 => \N__31464\,
            in3 => \N__31455\,
            lcout => \SIG_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i3_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__44648\,
            in1 => \N__32996\,
            in2 => \N__31434\,
            in3 => \N__44452\,
            lcout => \SIG_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i4_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__44453\,
            in1 => \N__44651\,
            in2 => \N__31425\,
            in3 => \N__32256\,
            lcout => \SIG_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i5_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__44649\,
            in1 => \N__44454\,
            in2 => \N__31416\,
            in3 => \N__33023\,
            lcout => \SIG_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i6_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__44455\,
            in1 => \N__44652\,
            in2 => \N__31407\,
            in3 => \N__41463\,
            lcout => \SIG_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56051\,
            ce => \N__43911\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12301_12302_set_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36912\,
            in1 => \N__36887\,
            in2 => \_gnd_net_\,
            in3 => \N__45033\,
            lcout => \comm_spi.n14822\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58358\,
            ce => 'H',
            sr => \N__37170\
        );

    \ADC_VDC.adc_state_i0_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010100"
        )
    port map (
            in0 => \N__51859\,
            in1 => \N__51722\,
            in2 => \N__52000\,
            in3 => \N__51345\,
            lcout => \ADC_VDC.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42372\,
            ce => \N__31686\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_3_lut_adj_28_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__51993\,
            in1 => \N__51858\,
            in2 => \_gnd_net_\,
            in3 => \N__51184\,
            lcout => \ADC_VDC.n21007\,
            ltout => \ADC_VDC.n21007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19461_3_lut_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000000"
        )
    port map (
            in0 => \N__51331\,
            in1 => \_gnd_net_\,
            in2 => \N__31386\,
            in3 => \N__51721\,
            lcout => \ADC_VDC.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_27_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51720\,
            in2 => \_gnd_net_\,
            in3 => \N__51330\,
            lcout => \ADC_VDC.n21133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_3_lut_4_lut_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__31707\,
            in1 => \N__51385\,
            in2 => \N__51754\,
            in3 => \N__51857\,
            lcout => \ADC_VDC.n15273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_33_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101010"
        )
    port map (
            in0 => \N__31701\,
            in1 => \N__51210\,
            in2 => \N__31695\,
            in3 => \N__31632\,
            lcout => \ADC_VDC.n42_adj_1452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_3_lut_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__34253\,
            in1 => \N__34273\,
            in2 => \_gnd_net_\,
            in3 => \N__34751\,
            lcout => \ADC_VDC.n20998\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_4_lut_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34750\,
            in1 => \N__34252\,
            in2 => \N__34275\,
            in3 => \N__34393\,
            lcout => \ADC_VDC.n11494\,
            ltout => \ADC_VDC.n11494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i3_4_lut_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__34297\,
            in1 => \N__31947\,
            in2 => \N__31665\,
            in3 => \N__34333\,
            lcout => \ADC_VDC.n15\,
            ltout => \ADC_VDC.n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18458_2_lut_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__51904\,
            in1 => \_gnd_net_\,
            in2 => \N__31635\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.n21185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__31608\,
            in1 => \N__51456\,
            in2 => \N__31497\,
            in3 => \N__32195\,
            lcout => buf_adcdata_vdc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42334\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18476_2_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34326\,
            in2 => \_gnd_net_\,
            in3 => \N__34296\,
            lcout => \ADC_VDC.n21203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18484_2_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34422\,
            in2 => \_gnd_net_\,
            in3 => \N__34359\,
            lcout => \ADC_VDC.n21211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101000"
        )
    port map (
            in0 => \N__51455\,
            in1 => \N__51896\,
            in2 => \N__51762\,
            in3 => \N__51209\,
            lcout => \ADC_VDC.n13368\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12325_12326_reset_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34806\,
            in1 => \N__52632\,
            in2 => \_gnd_net_\,
            in3 => \N__57474\,
            lcout => \comm_spi.n14847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58400\,
            ce => 'H',
            sr => \N__35226\
        );

    \i15_4_lut_adj_203_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31734\,
            in1 => \N__31791\,
            in2 => \N__34503\,
            in3 => \N__34578\,
            lcout => OPEN,
            ltout => \n20048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_204_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__31932\,
            in1 => \N__35115\,
            in2 => \N__31914\,
            in3 => \N__31911\,
            lcout => n14899,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i19_3_lut_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31902\,
            in1 => \N__31871\,
            in2 => \_gnd_net_\,
            in3 => \N__57184\,
            lcout => n19_adj_1673,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_200_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31844\,
            in1 => \N__31832\,
            in2 => \N__31821\,
            in3 => \N__31802\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_199_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31784\,
            in1 => \N__31772\,
            in2 => \N__31761\,
            in3 => \N__31745\,
            lcout => n26_adj_1656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15472_2_lut_3_lut_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__49496\,
            in1 => \N__54851\,
            in2 => \_gnd_net_\,
            in3 => \N__54341\,
            lcout => n14_adj_1552,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_158_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31953\,
            in1 => \N__34866\,
            in2 => \N__34728\,
            in3 => \N__34461\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i10_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32046\,
            in1 => \N__35533\,
            in2 => \_gnd_net_\,
            in3 => \N__35206\,
            lcout => req_data_cnt_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i11_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__31967\,
            in1 => \_gnd_net_\,
            in2 => \N__35556\,
            in3 => \N__35246\,
            lcout => req_data_cnt_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i15_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37476\,
            in1 => \N__35537\,
            in2 => \_gnd_net_\,
            in3 => \N__34480\,
            lcout => req_data_cnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i7_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35538\,
            in1 => \N__32270\,
            in2 => \_gnd_net_\,
            in3 => \N__46571\,
            lcout => req_data_cnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i30_3_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32019\,
            in1 => \N__32001\,
            in2 => \_gnd_net_\,
            in3 => \N__47258\,
            lcout => n30_adj_1611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_149_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37887\,
            in1 => \N__37962\,
            in2 => \N__31992\,
            in3 => \N__31966\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i5_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__39649\,
            in1 => \N__49388\,
            in2 => \N__52275\,
            in3 => \N__34919\,
            lcout => \buf_cfgRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i5_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35558\,
            in1 => \N__37250\,
            in2 => \_gnd_net_\,
            in3 => \N__32305\,
            lcout => req_data_cnt_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15471_2_lut_3_lut_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44061\,
            in1 => \N__54825\,
            in2 => \_gnd_net_\,
            in3 => \N__54501\,
            lcout => n14_adj_1551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i3_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36481\,
            in1 => \N__35557\,
            in2 => \_gnd_net_\,
            in3 => \N__41192\,
            lcout => req_data_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i4_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49387\,
            in1 => \N__32245\,
            in2 => \N__42707\,
            in3 => \N__41669\,
            lcout => buf_dds0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55944\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14639_3_lut_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32216\,
            in1 => \N__50720\,
            in2 => \_gnd_net_\,
            in3 => \N__57093\,
            lcout => n23_adj_1661,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__37092\,
            in1 => \N__32215\,
            in2 => \N__36756\,
            in3 => \N__32554\,
            lcout => n23_adj_1591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i4_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35559\,
            in1 => \N__36197\,
            in2 => \_gnd_net_\,
            in3 => \N__35336\,
            lcout => req_data_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i19_3_lut_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32202\,
            in1 => \N__32174\,
            in2 => \_gnd_net_\,
            in3 => \N__57023\,
            lcout => n19_adj_1616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i17_3_lut_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57024\,
            in1 => \N__32141\,
            in2 => \_gnd_net_\,
            in3 => \N__32089\,
            lcout => n17_adj_1672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i4_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__50983\,
            in1 => \N__37523\,
            in2 => \N__32391\,
            in3 => \N__53640\,
            lcout => comm_cmd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_153_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37668\,
            in1 => \N__41223\,
            in2 => \N__32306\,
            in3 => \N__41188\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__48821\,
            in1 => \N__53342\,
            in2 => \N__50990\,
            in3 => \N__37524\,
            lcout => comm_cmd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55950\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__32377\,
            in1 => \N__48847\,
            in2 => \_gnd_net_\,
            in3 => \N__48820\,
            lcout => n16818,
            ltout => \n16818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32364\,
            in3 => \N__47132\,
            lcout => n12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22365_bdd_4_lut_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__32361\,
            in1 => \N__32346\,
            in2 => \N__33084\,
            in3 => \N__47671\,
            lcout => n22368,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i26_3_lut_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__32334\,
            in1 => \N__57194\,
            in2 => \_gnd_net_\,
            in3 => \N__37667\,
            lcout => OPEN,
            ltout => \n26_adj_1630_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19711_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__57336\,
            in1 => \N__46297\,
            in2 => \N__32313\,
            in3 => \N__47672\,
            lcout => OPEN,
            ltout => \n22449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22449_bdd_4_lut_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47673\,
            in1 => \N__32976\,
            in2 => \N__32310\,
            in3 => \N__32307\,
            lcout => OPEN,
            ltout => \n22452_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1570065_i1_3_lut_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32283\,
            in2 => \N__32277\,
            in3 => \N__47243\,
            lcout => OPEN,
            ltout => \n30_adj_1631_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i5_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__53343\,
            in1 => \_gnd_net_\,
            in2 => \N__32640\,
            in3 => \N__54572\,
            lcout => comm_buf_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55954\,
            ce => \N__45212\,
            sr => \N__44016\
        );

    \equal_188_i9_2_lut_3_lut_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__46410\,
            in1 => \N__47667\,
            in2 => \_gnd_net_\,
            in3 => \N__57132\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18603_4_lut_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__57133\,
            in1 => \N__32625\,
            in2 => \N__32604\,
            in3 => \N__46411\,
            lcout => n21330,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_3_i23_3_lut_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32561\,
            in1 => \N__36214\,
            in2 => \_gnd_net_\,
            in3 => \N__57134\,
            lcout => n23_adj_1677,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i9_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__32518\,
            in1 => \N__53435\,
            in2 => \N__46767\,
            in3 => \N__46873\,
            lcout => buf_dds1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55963\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i19_3_lut_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32499\,
            in1 => \N__32468\,
            in2 => \_gnd_net_\,
            in3 => \N__57135\,
            lcout => n19_adj_1625,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_157_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__43844\,
            in1 => \N__43437\,
            in2 => \N__43649\,
            in3 => \N__43513\,
            lcout => OPEN,
            ltout => \n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_adj_160_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35316\,
            in1 => \N__32439\,
            in2 => \N__32430\,
            in3 => \N__32427\,
            lcout => n29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19285_2_lut_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__57136\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32412\,
            lcout => n21671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_3_i16_3_lut_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32997\,
            in1 => \N__32683\,
            in2 => \_gnd_net_\,
            in3 => \N__57147\,
            lcout => n16_adj_1640,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49280\,
            in1 => \N__42001\,
            in2 => \N__45645\,
            in3 => \N__44792\,
            lcout => buf_control_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i3_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000101110"
        )
    port map (
            in0 => \N__32687\,
            in1 => \N__46872\,
            in2 => \N__55434\,
            in3 => \N__36485\,
            lcout => buf_dds1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i0_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43198\,
            in1 => \N__47905\,
            in2 => \_gnd_net_\,
            in3 => \N__43676\,
            lcout => \acadc_skipCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i4_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__47907\,
            in1 => \_gnd_net_\,
            in2 => \N__36196\,
            in3 => \N__32660\,
            lcout => \acadc_skipCount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44165\,
            in1 => \N__36165\,
            in2 => \_gnd_net_\,
            in3 => \N__47906\,
            lcout => \acadc_skipCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36726\,
            in1 => \N__32659\,
            in2 => \N__36660\,
            in3 => \N__44164\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i6_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49279\,
            in1 => \N__47908\,
            in2 => \N__49497\,
            in3 => \N__43538\,
            lcout => \acadc_skipCount_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55974\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i7_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__32646\,
            in1 => \N__55432\,
            in2 => \N__49316\,
            in3 => \N__37989\,
            lcout => data_index_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55986\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6314_3_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44059\,
            in1 => \N__38008\,
            in2 => \_gnd_net_\,
            in3 => \N__41096\,
            lcout => n8_adj_1560,
            ltout => \n8_adj_1560_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49203\,
            in1 => \N__55431\,
            in2 => \N__32949\,
            in3 => \N__37988\,
            lcout => \data_index_9_N_212_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i7_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__44060\,
            in1 => \N__46598\,
            in2 => \N__47922\,
            in3 => \N__49207\,
            lcout => \acadc_skipCount_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55986\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_63_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36702\,
            in1 => \N__46594\,
            in2 => \N__36825\,
            in3 => \N__35392\,
            lcout => OPEN,
            ltout => \n22_adj_1590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_75_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32844\,
            in1 => \N__32838\,
            in2 => \N__32829\,
            in3 => \N__50592\,
            lcout => OPEN,
            ltout => \n30_adj_1543_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_79_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32826\,
            in1 => \N__36021\,
            in2 => \N__32820\,
            in3 => \N__32694\,
            lcout => n31_adj_1537,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i2_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__35393\,
            in1 => \_gnd_net_\,
            in2 => \N__47921\,
            in3 => \N__34860\,
            lcout => \acadc_skipCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55986\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i18_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38599\,
            in1 => \N__38748\,
            in2 => \N__32796\,
            in3 => \N__32749\,
            lcout => buf_adcdata_iac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_61_i14_2_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37113\,
            in2 => \_gnd_net_\,
            in3 => \N__33040\,
            lcout => OPEN,
            ltout => \n14_adj_1538_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__36801\,
            in1 => \N__32726\,
            in2 => \N__32697\,
            in3 => \N__32955\,
            lcout => n26_adj_1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i13_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38747\,
            in1 => \N__38600\,
            in2 => \N__33083\,
            in3 => \N__33113\,
            lcout => buf_adcdata_iac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i13_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__33041\,
            in1 => \N__49318\,
            in2 => \N__52286\,
            in3 => \N__47909\,
            lcout => \acadc_skipCount_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6324_3_lut_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41079\,
            in1 => \N__49494\,
            in2 => \_gnd_net_\,
            in3 => \N__38050\,
            lcout => n8_adj_1562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i5_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49134\,
            in1 => \N__33016\,
            in2 => \N__50424\,
            in3 => \N__41613\,
            lcout => buf_dds0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i5_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__47910\,
            in1 => \N__50418\,
            in2 => \N__49376\,
            in3 => \N__32975\,
            lcout => \acadc_skipCount_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55999\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i2_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__44515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44653\,
            lcout => dds_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i3_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36465\,
            in1 => \N__32995\,
            in2 => \_gnd_net_\,
            in3 => \N__41657\,
            lcout => buf_dds0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i3_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41162\,
            in1 => \N__36466\,
            in2 => \_gnd_net_\,
            in3 => \N__47916\,
            lcout => \acadc_skipCount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36681\,
            in1 => \N__32971\,
            in2 => \N__36867\,
            in3 => \N__41161\,
            lcout => n20_adj_1670,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i8_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38505\,
            in1 => \N__38771\,
            in2 => \N__41701\,
            in3 => \N__33810\,
            lcout => buf_adcdata_iac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i9_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__38506\,
            in1 => \N__38772\,
            in2 => \N__33783\,
            in3 => \N__43601\,
            lcout => buf_adcdata_iac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i8_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__39076\,
            in1 => \N__49322\,
            in2 => \N__41670\,
            in3 => \N__45634\,
            lcout => buf_dds0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56015\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_count_i0_i0_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33673\,
            in2 => \N__37785\,
            in3 => \_gnd_net_\,
            lcout => data_count_0,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => n19765,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33571\,
            in2 => \_gnd_net_\,
            in3 => \N__33549\,
            lcout => data_count_1,
            ltout => OPEN,
            carryin => n19765,
            carryout => n19766,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i2_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33460\,
            in2 => \_gnd_net_\,
            in3 => \N__33438\,
            lcout => data_count_2,
            ltout => OPEN,
            carryin => n19766,
            carryout => n19767,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i3_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33349\,
            in2 => \_gnd_net_\,
            in3 => \N__33327\,
            lcout => data_count_3,
            ltout => OPEN,
            carryin => n19767,
            carryout => n19768,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i4_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33247\,
            in2 => \_gnd_net_\,
            in3 => \N__33225\,
            lcout => data_count_4,
            ltout => OPEN,
            carryin => n19768,
            carryout => n19769,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i5_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33142\,
            in2 => \_gnd_net_\,
            in3 => \N__33117\,
            lcout => data_count_5,
            ltout => OPEN,
            carryin => n19769,
            carryout => n19770,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i6_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34153\,
            in2 => \_gnd_net_\,
            in3 => \N__34131\,
            lcout => data_count_6,
            ltout => OPEN,
            carryin => n19770,
            carryout => n19771,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i7_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34045\,
            in2 => \_gnd_net_\,
            in3 => \N__34023\,
            lcout => data_count_7,
            ltout => OPEN,
            carryin => n19771,
            carryout => n19772,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__37843\,
            sr => \N__38139\
        );

    \data_count_i0_i8_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33937\,
            in2 => \_gnd_net_\,
            in3 => \N__33915\,
            lcout => data_count_8,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => n19773,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__37845\,
            sr => \N__38149\
        );

    \data_count_i0_i9_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33835\,
            in2 => \_gnd_net_\,
            in3 => \N__33912\,
            lcout => data_count_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__37845\,
            sr => \N__38149\
        );

    \comm_spi.imosi_44_12287_12288_reset_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50884\,
            lcout => \comm_spi.n14809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55937\,
            ce => 'H',
            sr => \N__50832\
        );

    \comm_spi.data_rx_i0_12301_12302_reset_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36911\,
            in1 => \N__36886\,
            in2 => \_gnd_net_\,
            in3 => \N__45032\,
            lcout => \comm_spi.n14823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58352\,
            ce => 'H',
            sr => \N__39774\
        );

    \comm_spi.i19525_4_lut_3_lut_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36970\,
            in1 => \N__50466\,
            in2 => \_gnd_net_\,
            in3 => \N__58121\,
            lcout => \comm_spi.n23083\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19500_4_lut_3_lut_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__58120\,
            in1 => \N__33816\,
            in2 => \_gnd_net_\,
            in3 => \N__39785\,
            lcout => \comm_spi.n23089\,
            ltout => \comm_spi.n23089_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12303_3_lut_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34455\,
            in2 => \N__34449\,
            in3 => \N__34446\,
            lcout => comm_rx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_12287_12288_set_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50892\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55938\,
            ce => 'H',
            sr => \N__37158\
        );

    \ADC_VDC.bit_cnt_3771__i0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34429\,
            in2 => \_gnd_net_\,
            in3 => \N__34404\,
            lcout => \ADC_VDC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \ADC_VDC.n19918\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34397\,
            in2 => \_gnd_net_\,
            in3 => \N__34377\,
            lcout => \ADC_VDC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19918\,
            carryout => \ADC_VDC.n19919\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34373\,
            in2 => \_gnd_net_\,
            in3 => \N__34341\,
            lcout => \ADC_VDC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19919\,
            carryout => \ADC_VDC.n19920\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34337\,
            in2 => \_gnd_net_\,
            in3 => \N__34308\,
            lcout => \ADC_VDC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19920\,
            carryout => \ADC_VDC.n19921\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34301\,
            in2 => \_gnd_net_\,
            in3 => \N__34278\,
            lcout => \ADC_VDC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19921\,
            carryout => \ADC_VDC.n19922\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34274\,
            in2 => \_gnd_net_\,
            in3 => \N__34257\,
            lcout => \ADC_VDC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19922\,
            carryout => \ADC_VDC.n19923\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i6_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34254\,
            in2 => \_gnd_net_\,
            in3 => \N__34239\,
            lcout => \ADC_VDC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19923\,
            carryout => \ADC_VDC.n19924\,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \ADC_VDC.bit_cnt_3771__i7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34752\,
            in2 => \_gnd_net_\,
            in3 => \N__34755\,
            lcout => \ADC_VDC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42221\,
            ce => \N__51075\,
            sr => \N__34737\
        );

    \i1_4_lut_adj_311_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__55346\,
            in1 => \N__37182\,
            in2 => \N__49392\,
            in3 => \N__35460\,
            lcout => n12662,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_150_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__37929\,
            in1 => \N__40683\,
            in2 => \N__35214\,
            in3 => \N__34879\,
            lcout => n21_adj_1594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_58_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39744\,
            in1 => \N__40002\,
            in2 => \N__40080\,
            in3 => \N__39966\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SecClk_292_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__34693\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34664\,
            lcout => \TEST_LED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50783\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34647\,
            in1 => \N__34629\,
            in2 => \N__34611\,
            in3 => \N__34593\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_198_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34572\,
            in1 => \N__34553\,
            in2 => \N__34539\,
            in3 => \N__34518\,
            lcout => n28_adj_1554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_146_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37863\,
            in1 => \N__43086\,
            in2 => \N__34487\,
            in3 => \N__42994\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19343_2_lut_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57186\,
            in2 => \_gnd_net_\,
            in3 => \N__34880\,
            lcout => n21703,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_93_2_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58066\,
            lcout => \comm_spi.data_tx_7__N_807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i12_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37196\,
            in1 => \N__35508\,
            in2 => \_gnd_net_\,
            in3 => \N__34881\,
            lcout => req_data_cnt_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i9_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35510\,
            in1 => \N__37445\,
            in2 => \_gnd_net_\,
            in3 => \N__42995\,
            lcout => req_data_cnt_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_148_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__37725\,
            in1 => \N__46527\,
            in2 => \N__35374\,
            in3 => \N__46567\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19520_4_lut_3_lut_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34804\,
            in1 => \N__53685\,
            in2 => \_gnd_net_\,
            in3 => \N__58067\,
            lcout => \comm_spi.n23095\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i2_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__34851\,
            in1 => \N__35509\,
            in2 => \N__35375\,
            in3 => \_gnd_net_\,
            lcout => req_data_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55943\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12325_12326_set_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34805\,
            in1 => \N__52631\,
            in2 => \_gnd_net_\,
            in3 => \N__57470\,
            lcout => \comm_spi.n14846\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58401\,
            ce => 'H',
            sr => \N__34788\
        );

    \i19332_2_lut_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57213\,
            in2 => \_gnd_net_\,
            in3 => \N__34776\,
            lcout => n21702,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19431_2_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35811\,
            in2 => \_gnd_net_\,
            in3 => \N__37035\,
            lcout => n14915,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35148\,
            in2 => \_gnd_net_\,
            in3 => \N__35130\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19746_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__35109\,
            in1 => \N__46402\,
            in2 => \N__35094\,
            in3 => \N__47729\,
            lcout => n22485,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18442_2_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37570\,
            in2 => \_gnd_net_\,
            in3 => \N__53997\,
            lcout => n11652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_3_i19_3_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35076\,
            in1 => \N__35045\,
            in2 => \_gnd_net_\,
            in3 => \N__57099\,
            lcout => n19_adj_1641,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i20_3_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57098\,
            in1 => \N__35025\,
            in2 => \_gnd_net_\,
            in3 => \N__34998\,
            lcout => n20_adj_1674,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_287_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__55207\,
            in1 => \N__55544\,
            in2 => \N__35280\,
            in3 => \N__54803\,
            lcout => n16821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i16_3_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__57101\,
            in1 => \_gnd_net_\,
            in2 => \N__35309\,
            in3 => \N__34971\,
            lcout => n16_adj_1664,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i20_3_lut_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34918\,
            in1 => \N__34902\,
            in2 => \_gnd_net_\,
            in3 => \N__57100\,
            lcout => n20_adj_1667,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_263_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011111"
        )
    port map (
            in0 => \N__54517\,
            in1 => \N__48237\,
            in2 => \N__54788\,
            in3 => \N__55298\,
            lcout => OPEN,
            ltout => \n12082_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_189_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__35279\,
            in1 => \N__48341\,
            in2 => \N__35256\,
            in3 => \N__55562\,
            lcout => n12089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i6_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__50952\,
            in1 => \N__37496\,
            in2 => \N__53235\,
            in3 => \N__48851\,
            lcout => comm_cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15463_2_lut_3_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45302\,
            in1 => \N__54710\,
            in2 => \_gnd_net_\,
            in3 => \N__54518\,
            lcout => n14_adj_1573,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_101_2_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50455\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58065\,
            lcout => \comm_spi.data_tx_7__N_817\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i24_3_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35736\,
            in1 => \N__57163\,
            in2 => \_gnd_net_\,
            in3 => \N__35210\,
            lcout => n24_adj_1686,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_300_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__54706\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55297\,
            lcout => n12442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i7_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37497\,
            in1 => \N__50953\,
            in2 => \N__48598\,
            in3 => \N__49993\,
            lcout => comm_cmd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55958\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__47675\,
            in1 => \N__35187\,
            in2 => \N__35175\,
            in3 => \N__46465\,
            lcout => OPEN,
            ltout => \n22641_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22641_bdd_4_lut_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__38238\,
            in1 => \N__35442\,
            in2 => \N__35430\,
            in3 => \N__47676\,
            lcout => n22644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i26_3_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35427\,
            in1 => \N__57195\,
            in2 => \_gnd_net_\,
            in3 => \N__37717\,
            lcout => OPEN,
            ltout => \n26_adj_1647_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19673_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__46466\,
            in1 => \N__42570\,
            in2 => \N__35403\,
            in3 => \N__47677\,
            lcout => OPEN,
            ltout => \n22383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22383_bdd_4_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47678\,
            in1 => \N__35400\,
            in2 => \N__35379\,
            in3 => \N__35376\,
            lcout => OPEN,
            ltout => \n22386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1568256_i1_3_lut_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__47233\,
            in1 => \N__35352\,
            in2 => \N__35346\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n30_adj_1648_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__50158\,
            in1 => \_gnd_net_\,
            in2 => \N__35343\,
            in3 => \N__54499\,
            lcout => comm_buf_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55967\,
            ce => \N__45195\,
            sr => \N__44002\
        );

    \i2_3_lut_adj_266_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__47232\,
            in1 => \N__46290\,
            in2 => \_gnd_net_\,
            in3 => \N__47674\,
            lcout => n66,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_154_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__44194\,
            in1 => \N__37690\,
            in2 => \N__35340\,
            in3 => \N__44140\,
            lcout => n18_adj_1644,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i13_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__35299\,
            in1 => \N__49311\,
            in2 => \N__52276\,
            in3 => \N__41644\,
            lcout => buf_dds0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_267_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__35643\,
            in1 => \N__48259\,
            in2 => \_gnd_net_\,
            in3 => \N__57146\,
            lcout => n20011,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i14_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__35629\,
            in1 => \N__49537\,
            in2 => \N__46910\,
            in3 => \N__46764\,
            lcout => buf_dds1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i7_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__46890\,
            in1 => \N__36568\,
            in2 => \N__44078\,
            in3 => \N__46765\,
            lcout => buf_dds1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i1_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__46763\,
            in1 => \N__53510\,
            in2 => \N__35602\,
            in3 => \N__46894\,
            lcout => buf_dds1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i1_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__44141\,
            in1 => \_gnd_net_\,
            in2 => \N__36166\,
            in3 => \N__35555\,
            lcout => req_data_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55978\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i1_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__53436\,
            in1 => \N__41989\,
            in2 => \N__49361\,
            in3 => \N__42937\,
            lcout => \DDS_RNG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_271_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__48266\,
            in1 => \N__49272\,
            in2 => \N__35478\,
            in3 => \N__55455\,
            lcout => n12144,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_4_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__46377\,
            in1 => \N__47643\,
            in2 => \N__57209\,
            in3 => \N__53988\,
            lcout => n7_adj_1650,
            ltout => \n7_adj_1650_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_283_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__54738\,
            in1 => \N__54487\,
            in2 => \N__35463\,
            in3 => \N__35456\,
            lcout => n10756,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i3_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41988\,
            in1 => \N__45326\,
            in2 => \N__49355\,
            in3 => \N__36215\,
            lcout => \SELIRNG1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15465_2_lut_3_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__54740\,
            in1 => \N__42710\,
            in2 => \_gnd_net_\,
            in3 => \N__54489\,
            lcout => n14_adj_1546,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15468_2_lut_3_lut_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__54488\,
            in1 => \N__53511\,
            in2 => \_gnd_net_\,
            in3 => \N__54739\,
            lcout => n14_adj_1549,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__55436\,
            in1 => \N__49209\,
            in2 => \N__38034\,
            in3 => \N__36128\,
            lcout => \data_index_9_N_212_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_78_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36546\,
            in1 => \N__43534\,
            in2 => \N__36846\,
            in3 => \N__43672\,
            lcout => n17_adj_1553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i5_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__52277\,
            in1 => \N__49215\,
            in2 => \N__35989\,
            in3 => \N__41990\,
            lcout => \AMPV_POW\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_256_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__55563\,
            in1 => \N__36513\,
            in2 => \N__49317\,
            in3 => \N__55438\,
            lcout => n11611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55435\,
            in1 => \N__49208\,
            in2 => \N__36237\,
            in3 => \N__38078\,
            lcout => \data_index_9_N_212_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19459_2_lut_3_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35880\,
            in1 => \N__35807\,
            in2 => \_gnd_net_\,
            in3 => \N__35710\,
            lcout => n21226,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i2_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__45718\,
            in1 => \N__49214\,
            in2 => \N__45869\,
            in3 => \N__41991\,
            lcout => \SELIRNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_268_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__49210\,
            in1 => \N__36512\,
            in2 => \_gnd_net_\,
            in3 => \N__55437\,
            lcout => n12596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i22_3_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36301\,
            in1 => \N__36501\,
            in2 => \_gnd_net_\,
            in3 => \N__47733\,
            lcout => n22_adj_1617,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15466_2_lut_3_lut_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__54553\,
            in1 => \N__45282\,
            in2 => \_gnd_net_\,
            in3 => \N__54826\,
            lcout => n14_adj_1547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6344_3_lut_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42708\,
            in1 => \N__38182\,
            in2 => \_gnd_net_\,
            in3 => \N__41101\,
            lcout => n8_adj_1564,
            ltout => \n8_adj_1564_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49132\,
            in1 => \N__55439\,
            in2 => \N__36441\,
            in3 => \N__38195\,
            lcout => \data_index_9_N_212_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i1_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__36302\,
            in1 => \N__38749\,
            in2 => \N__36351\,
            in3 => \N__38601\,
            lcout => buf_adcdata_iac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i16_3_lut_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36288\,
            in1 => \N__36258\,
            in2 => \_gnd_net_\,
            in3 => \N__57239\,
            lcout => n16_adj_1671,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6354_3_lut_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45281\,
            in1 => \N__38096\,
            in2 => \_gnd_net_\,
            in3 => \N__41100\,
            lcout => n8_adj_1566,
            ltout => \n8_adj_1566_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i3_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49133\,
            in1 => \N__55440\,
            in2 => \N__36636\,
            in3 => \N__38079\,
            lcout => data_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i7_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__38789\,
            in1 => \N__36633\,
            in2 => \N__44491\,
            in3 => \N__44629\,
            lcout => \SIG_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56036\,
            ce => \N__43903\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.i23_4_lut_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000010101"
        )
    port map (
            in0 => \N__44445\,
            in1 => \N__43926\,
            in2 => \N__44753\,
            in3 => \N__44628\,
            lcout => \SIG_DDS.n9_adj_1434\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19478_4_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111110"
        )
    port map (
            in0 => \N__44626\,
            in1 => \N__44744\,
            in2 => \N__43936\,
            in3 => \N__44444\,
            lcout => \SIG_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19199_2_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36612\,
            in2 => \_gnd_net_\,
            in3 => \N__44627\,
            lcout => \SIG_DDS.n21744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i16_3_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36569\,
            in1 => \N__38788\,
            in2 => \_gnd_net_\,
            in3 => \N__57238\,
            lcout => n16_adj_1620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i0_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37772\,
            in2 => \N__36545\,
            in3 => \_gnd_net_\,
            lcout => acadc_skipcnt_0,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => n19789,
            clk => \INVacadc_skipcnt_i0_i0C_net\,
            ce => \N__37043\,
            sr => \N__36525\
        );

    \add_73_2_THRU_CRY_0_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58702\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => n19789,
            carryout => \n19789_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58706\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19789_THRU_CRY_0_THRU_CO\,
            carryout => \n19789_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_2_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58703\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19789_THRU_CRY_1_THRU_CO\,
            carryout => \n19789_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_3_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58707\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19789_THRU_CRY_2_THRU_CO\,
            carryout => \n19789_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_4_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58704\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19789_THRU_CRY_3_THRU_CO\,
            carryout => \n19789_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_5_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58708\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19789_THRU_CRY_4_THRU_CO\,
            carryout => \n19789_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_6_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58705\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19789_THRU_CRY_5_THRU_CO\,
            carryout => \n19789_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i1_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36719\,
            in2 => \_gnd_net_\,
            in3 => \N__36705\,
            lcout => acadc_skipcnt_1,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => n19790,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i2_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36698\,
            in2 => \_gnd_net_\,
            in3 => \N__36684\,
            lcout => acadc_skipcnt_2,
            ltout => OPEN,
            carryin => n19790,
            carryout => n19791,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i3_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36680\,
            in2 => \_gnd_net_\,
            in3 => \N__36663\,
            lcout => acadc_skipcnt_3,
            ltout => OPEN,
            carryin => n19791,
            carryout => n19792,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i4_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36653\,
            in2 => \_gnd_net_\,
            in3 => \N__36639\,
            lcout => acadc_skipcnt_4,
            ltout => OPEN,
            carryin => n19792,
            carryout => n19793,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i5_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36863\,
            in2 => \_gnd_net_\,
            in3 => \N__36849\,
            lcout => acadc_skipcnt_5,
            ltout => OPEN,
            carryin => n19793,
            carryout => n19794,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i6_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36842\,
            in2 => \_gnd_net_\,
            in3 => \N__36828\,
            lcout => acadc_skipcnt_6,
            ltout => OPEN,
            carryin => n19794,
            carryout => n19795,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i7_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36818\,
            in2 => \_gnd_net_\,
            in3 => \N__36804\,
            lcout => acadc_skipcnt_7,
            ltout => OPEN,
            carryin => n19795,
            carryout => n19796,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i8_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36797\,
            in2 => \_gnd_net_\,
            in3 => \N__36783\,
            lcout => acadc_skipcnt_8,
            ltout => OPEN,
            carryin => n19796,
            carryout => n19797,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__37042\,
            sr => \N__36999\
        );

    \acadc_skipcnt_i0_i9_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36776\,
            in2 => \_gnd_net_\,
            in3 => \N__36762\,
            lcout => acadc_skipcnt_9,
            ltout => OPEN,
            carryin => \bfn_13_20_0_\,
            carryout => n19798,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \acadc_skipcnt_i0_i10_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50663\,
            in2 => \_gnd_net_\,
            in3 => \N__36759\,
            lcout => acadc_skipcnt_10,
            ltout => OPEN,
            carryin => n19798,
            carryout => n19799,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \acadc_skipcnt_i0_i11_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36746\,
            in2 => \_gnd_net_\,
            in3 => \N__36732\,
            lcout => acadc_skipcnt_11,
            ltout => OPEN,
            carryin => n19799,
            carryout => n19800,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \acadc_skipcnt_i0_i12_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50621\,
            in2 => \_gnd_net_\,
            in3 => \N__36729\,
            lcout => acadc_skipcnt_12,
            ltout => OPEN,
            carryin => n19800,
            carryout => n19801,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \acadc_skipcnt_i0_i13_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37109\,
            in2 => \_gnd_net_\,
            in3 => \N__37095\,
            lcout => acadc_skipcnt_13,
            ltout => OPEN,
            carryin => n19801,
            carryout => n19802,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \acadc_skipcnt_i0_i14_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37085\,
            in2 => \_gnd_net_\,
            in3 => \N__37071\,
            lcout => acadc_skipcnt_14,
            ltout => OPEN,
            carryin => n19802,
            carryout => n19803,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \acadc_skipcnt_i0_i15_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37058\,
            in2 => \_gnd_net_\,
            in3 => \N__37068\,
            lcout => acadc_skipcnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__37044\,
            sr => \N__36998\
        );

    \comm_spi.imiso_83_12297_12298_reset_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39813\,
            in1 => \N__39797\,
            in2 => \_gnd_net_\,
            in3 => \N__44331\,
            lcout => \comm_spi.n14819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12297_12298_resetC_net\,
            ce => 'H',
            sr => \N__42888\
        );

    \comm_spi.data_tx_i7_12294_12295_reset_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36972\,
            in1 => \N__36954\,
            in2 => \_gnd_net_\,
            in3 => \N__36933\,
            lcout => \comm_spi.n14816\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58356\,
            ce => 'H',
            sr => \N__42887\
        );

    \comm_spi.data_tx_i7_12294_12295_set_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36971\,
            in1 => \N__36950\,
            in2 => \_gnd_net_\,
            in3 => \N__36929\,
            lcout => \comm_spi.n14815\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58257\,
            ce => 'H',
            sr => \N__42836\
        );

    \ADC_VDC.genclk.t_clk_24_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56586\,
            lcout => \VDC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t_clk_24C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39758\,
            in1 => \N__39692\,
            in2 => \N__40038\,
            in3 => \N__39707\,
            lcout => n33,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12289_3_lut_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36904\,
            in1 => \N__36891\,
            in2 => \_gnd_net_\,
            in3 => \N__45025\,
            lcout => \comm_spi.imosi\,
            ltout => \comm_spi.imosi_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_86_2_lut_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37173\,
            in3 => \N__58059\,
            lcout => \comm_spi.DOUT_7__N_786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_88_2_lut_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50891\,
            in2 => \_gnd_net_\,
            in3 => \N__58058\,
            lcout => \comm_spi.imosi_N_792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__39722\,
            in1 => \N__39677\,
            in2 => \N__40113\,
            in3 => \N__40163\,
            lcout => n30_adj_1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40358\,
            in1 => \N__40343\,
            in2 => \N__40131\,
            in3 => \N__40094\,
            lcout => OPEN,
            ltout => \n12_adj_1542_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__39980\,
            in1 => \N__40211\,
            in2 => \N__37149\,
            in3 => \N__40227\,
            lcout => OPEN,
            ltout => \n19986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__39944\,
            in1 => \N__40016\,
            in2 => \N__37146\,
            in3 => \N__37143\,
            lcout => OPEN,
            ltout => \n34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18_4_lut_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37119\,
            in1 => \N__37137\,
            in2 => \N__37131\,
            in3 => \N__37128\,
            lcout => n49,
            ltout => \n49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \wdtick_flag_289_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37122\,
            in3 => \N__44815\,
            lcout => wdtick_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50784\,
            ce => 'H',
            sr => \N__42151\
        );

    \i13_4_lut_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40178\,
            in1 => \N__40193\,
            in2 => \N__40149\,
            in3 => \N__40056\,
            lcout => n32,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.bit_cnt_3767__i3_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__37296\,
            in1 => \N__42791\,
            in2 => \N__37281\,
            in3 => \N__37314\,
            lcout => \comm_spi.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__58165\
        );

    \comm_spi.bit_cnt_3767__i2_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__37313\,
            in1 => \N__37277\,
            in2 => \_gnd_net_\,
            in3 => \N__37295\,
            lcout => \comm_spi.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__58165\
        );

    \comm_spi.bit_cnt_3767__i1_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37312\,
            lcout => \comm_spi.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__58165\
        );

    \comm_spi.bit_cnt_3767__i0_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37275\,
            lcout => \comm_spi.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i3C_net\,
            ce => 'H',
            sr => \N__58165\
        );

    \comm_cmd_1__bdd_4_lut_19721_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__37335\,
            in1 => \N__46462\,
            in2 => \N__37323\,
            in3 => \N__47697\,
            lcout => n22461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i2_3_lut_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__37311\,
            in1 => \N__37294\,
            in2 => \_gnd_net_\,
            in3 => \N__37274\,
            lcout => \comm_spi.n17254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15452_2_lut_3_lut_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__50414\,
            in1 => \N__54506\,
            in2 => \N__54853\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_1579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15462_2_lut_3_lut_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__54504\,
            in1 => \N__54796\,
            in2 => \_gnd_net_\,
            in3 => \N__47786\,
            lcout => n14_adj_1572,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__46461\,
            in1 => \N__47696\,
            in2 => \N__57262\,
            in3 => \N__53969\,
            lcout => n4_adj_1637,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15469_2_lut_3_lut_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__54503\,
            in1 => \N__54795\,
            in2 => \_gnd_net_\,
            in3 => \N__42517\,
            lcout => n14_adj_1544,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15470_2_lut_3_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54505\,
            in2 => \N__54852\,
            in3 => \N__53423\,
            lcout => n14_adj_1575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19687_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__47698\,
            in1 => \N__37431\,
            in2 => \N__37422\,
            in3 => \N__46463\,
            lcout => OPEN,
            ltout => \n22413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22413_bdd_4_lut_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__37413\,
            in1 => \N__37407\,
            in2 => \N__37398\,
            in3 => \N__47699\,
            lcout => n22416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19847_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__46464\,
            in1 => \N__41754\,
            in2 => \N__37395\,
            in3 => \N__47700\,
            lcout => OPEN,
            ltout => \n22569_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22569_bdd_4_lut_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47701\,
            in1 => \N__37380\,
            in2 => \N__37365\,
            in3 => \N__37362\,
            lcout => OPEN,
            ltout => \n22572_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1565844_i1_3_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37356\,
            in2 => \N__37350\,
            in3 => \N__47267\,
            lcout => OPEN,
            ltout => \n30_adj_1669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i5_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53292\,
            in2 => \N__37347\,
            in3 => \N__54510\,
            lcout => comm_buf_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55959\,
            ce => \N__43325\,
            sr => \N__43249\
        );

    \comm_buf_0__i7_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__48572\,
            in1 => \N__54509\,
            in2 => \_gnd_net_\,
            in3 => \N__37344\,
            lcout => comm_buf_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55968\,
            ce => \N__43338\,
            sr => \N__43275\
        );

    \comm_buf_0__i6_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54507\,
            in1 => \N__53195\,
            in2 => \_gnd_net_\,
            in3 => \N__37629\,
            lcout => comm_buf_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55968\,
            ce => \N__43338\,
            sr => \N__43275\
        );

    \comm_buf_0__i3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__49856\,
            in1 => \N__54508\,
            in2 => \_gnd_net_\,
            in3 => \N__37614\,
            lcout => comm_buf_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55968\,
            ce => \N__43338\,
            sr => \N__43275\
        );

    \i22_4_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100001010"
        )
    port map (
            in0 => \N__52884\,
            in1 => \N__46038\,
            in2 => \N__54005\,
            in3 => \N__54737\,
            lcout => OPEN,
            ltout => \n8_adj_1689_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i2_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__52797\,
            in1 => \N__37545\,
            in2 => \N__37602\,
            in3 => \N__54494\,
            lcout => comm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55979\,
            ce => \N__37596\,
            sr => \N__55478\
        );

    \i1_4_lut_adj_285_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100111000"
        )
    port map (
            in0 => \N__52883\,
            in1 => \N__54685\,
            in2 => \N__54552\,
            in3 => \N__52799\,
            lcout => OPEN,
            ltout => \n26_adj_1595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19442_2_lut_3_lut_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55183\,
            in2 => \N__37599\,
            in3 => \N__53982\,
            lcout => n18_adj_1615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19360_4_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__53981\,
            in1 => \N__52798\,
            in2 => \N__54810\,
            in3 => \N__37590\,
            lcout => n21714,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i22_4_lut_4_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001000100"
        )
    port map (
            in0 => \N__54498\,
            in1 => \N__53980\,
            in2 => \N__52803\,
            in3 => \N__52882\,
            lcout => OPEN,
            ltout => \n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_241_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__55182\,
            in1 => \N__54684\,
            in2 => \N__37539\,
            in3 => \N__55553\,
            lcout => n12107,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_44_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__54683\,
            in1 => \N__55181\,
            in2 => \_gnd_net_\,
            in3 => \N__54490\,
            lcout => n21147,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_cntvec_i0_i0_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43840\,
            in2 => \N__37784\,
            in3 => \_gnd_net_\,
            lcout => data_cntvec_0,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => n19774,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44195\,
            in2 => \_gnd_net_\,
            in3 => \N__37728\,
            lcout => data_cntvec_1,
            ltout => OPEN,
            carryin => n19774,
            carryout => n19775,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i2_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37721\,
            in2 => \_gnd_net_\,
            in3 => \N__37701\,
            lcout => data_cntvec_2,
            ltout => OPEN,
            carryin => n19775,
            carryout => n19776,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i3_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41219\,
            in2 => \_gnd_net_\,
            in3 => \N__37698\,
            lcout => data_cntvec_3,
            ltout => OPEN,
            carryin => n19776,
            carryout => n19777,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i4_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37691\,
            in2 => \_gnd_net_\,
            in3 => \N__37671\,
            lcout => data_cntvec_4,
            ltout => OPEN,
            carryin => n19777,
            carryout => n19778,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i5_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37660\,
            in2 => \_gnd_net_\,
            in3 => \N__37638\,
            lcout => data_cntvec_5,
            ltout => OPEN,
            carryin => n19778,
            carryout => n19779,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i6_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43436\,
            in2 => \_gnd_net_\,
            in3 => \N__37635\,
            lcout => data_cntvec_6,
            ltout => OPEN,
            carryin => n19779,
            carryout => n19780,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i7_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46519\,
            in2 => \_gnd_net_\,
            in3 => \N__37632\,
            lcout => data_cntvec_7,
            ltout => OPEN,
            carryin => n19780,
            carryout => n19781,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__37842\,
            sr => \N__38151\
        );

    \data_cntvec_i0_i8_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40901\,
            in2 => \_gnd_net_\,
            in3 => \N__37971\,
            lcout => data_cntvec_8,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => n19782,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i9_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43078\,
            in2 => \_gnd_net_\,
            in3 => \N__37968\,
            lcout => data_cntvec_9,
            ltout => OPEN,
            carryin => n19782,
            carryout => n19783,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i10_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40678\,
            in2 => \_gnd_net_\,
            in3 => \N__37965\,
            lcout => data_cntvec_10,
            ltout => OPEN,
            carryin => n19783,
            carryout => n19784,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i11_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37954\,
            in2 => \_gnd_net_\,
            in3 => \N__37932\,
            lcout => data_cntvec_11,
            ltout => OPEN,
            carryin => n19784,
            carryout => n19785,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i12_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37925\,
            in2 => \_gnd_net_\,
            in3 => \N__37911\,
            lcout => data_cntvec_12,
            ltout => OPEN,
            carryin => n19785,
            carryout => n19786,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i13_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37904\,
            in2 => \_gnd_net_\,
            in3 => \N__37890\,
            lcout => data_cntvec_13,
            ltout => OPEN,
            carryin => n19786,
            carryout => n19787,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i14_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37883\,
            in2 => \_gnd_net_\,
            in3 => \N__37869\,
            lcout => data_cntvec_14,
            ltout => OPEN,
            carryin => n19787,
            carryout => n19788,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \data_cntvec_i0_i15_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37859\,
            in2 => \_gnd_net_\,
            in3 => \N__37866\,
            lcout => data_cntvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__37844\,
            sr => \N__38150\
        );

    \add_125_2_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41141\,
            in1 => \N__41140\,
            in2 => \N__38927\,
            in3 => \N__38106\,
            lcout => n7_adj_1539,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => n19804,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_3_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39357\,
            in1 => \N__39356\,
            in2 => \N__38931\,
            in3 => \N__38103\,
            lcout => n7_adj_1569,
            ltout => OPEN,
            carryin => n19804,
            carryout => n19805,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39222\,
            in1 => \N__39221\,
            in2 => \N__38928\,
            in3 => \N__38100\,
            lcout => n7_adj_1567,
            ltout => OPEN,
            carryin => n19805,
            carryout => n19806,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_5_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38097\,
            in1 => \N__38095\,
            in2 => \N__38932\,
            in3 => \N__38067\,
            lcout => n7_adj_1565,
            ltout => OPEN,
            carryin => n19806,
            carryout => n19807,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_6_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38184\,
            in1 => \N__38183\,
            in2 => \N__38929\,
            in3 => \N__38064\,
            lcout => n7_adj_1563,
            ltout => OPEN,
            carryin => n19807,
            carryout => n19808,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_7_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39057\,
            in1 => \N__39056\,
            in2 => \N__38933\,
            in3 => \N__38061\,
            lcout => n17703,
            ltout => OPEN,
            carryin => n19808,
            carryout => n19809,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_8_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38058\,
            in1 => \N__38057\,
            in2 => \N__38930\,
            in3 => \N__38013\,
            lcout => n7_adj_1561,
            ltout => OPEN,
            carryin => n19809,
            carryout => n19810,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_9_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38010\,
            in1 => \N__38009\,
            in2 => \N__38934\,
            in3 => \N__37977\,
            lcout => n7_adj_1559,
            ltout => OPEN,
            carryin => n19810,
            carryout => n19811,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_10_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__39177\,
            in1 => \N__39176\,
            in2 => \N__38944\,
            in3 => \N__37974\,
            lcout => n7_adj_1557,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => n19812,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_11_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38962\,
            in1 => \N__38963\,
            in2 => \N__38945\,
            in3 => \N__38859\,
            lcout => n7_adj_1555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i30_3_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__38856\,
            in1 => \N__38835\,
            in2 => \_gnd_net_\,
            in3 => \N__47271\,
            lcout => n30_adj_1618,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds1_305_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000001100100"
        )
    port map (
            in0 => \N__49061\,
            in1 => \N__55459\,
            in2 => \N__38810\,
            in3 => \N__46938\,
            lcout => trig_dds1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15204_3_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50422\,
            in1 => \N__39055\,
            in2 => \_gnd_net_\,
            in3 => \N__41102\,
            lcout => n17705,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i6_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49059\,
            in1 => \N__41456\,
            in2 => \N__49495\,
            in3 => \N__41614\,
            lcout => buf_dds0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i7_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49060\,
            in1 => \N__38790\,
            in2 => \N__44082\,
            in3 => \N__41615\,
            lcout => buf_dds0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i10_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__38773\,
            in1 => \N__38570\,
            in2 => \N__38236\,
            in3 => \N__38263\,
            lcout => buf_adcdata_iac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i4_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__38205\,
            in1 => \N__55294\,
            in2 => \N__49258\,
            in3 => \N__38199\,
            lcout => data_index_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds0_304_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__55292\,
            in1 => \N__49127\,
            in2 => \N__43944\,
            in3 => \N__38163\,
            lcout => trig_dds0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19663_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__39460\,
            in1 => \N__57212\,
            in2 => \N__39150\,
            in3 => \N__46467\,
            lcout => OPEN,
            ltout => \n22389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22389_bdd_4_lut_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__46468\,
            in1 => \N__39111\,
            in2 => \N__39084\,
            in3 => \N__39077\,
            lcout => n22392,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i9_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49126\,
            in1 => \N__41900\,
            in2 => \N__41922\,
            in3 => \N__55295\,
            lcout => data_index_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i5_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__55293\,
            in1 => \N__41439\,
            in2 => \N__41424\,
            in3 => \N__49131\,
            lcout => data_index_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56053\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.SCLK_27_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001000110001"
        )
    port map (
            in0 => \N__44409\,
            in1 => \N__44670\,
            in2 => \N__39026\,
            in3 => \N__44752\,
            lcout => \DDS_SCK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.MOSI_31_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__39009\,
            in1 => \N__44408\,
            in2 => \_gnd_net_\,
            in3 => \N__38975\,
            lcout => \DDS_MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i1_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__49124\,
            in1 => \N__39336\,
            in2 => \N__55479\,
            in3 => \N__39327\,
            lcout => data_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6294_3_lut_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__53437\,
            in1 => \N__38964\,
            in2 => \_gnd_net_\,
            in3 => \N__41119\,
            lcout => n8_adj_1556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6364_3_lut_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41120\,
            in1 => \N__45465\,
            in2 => \_gnd_net_\,
            in3 => \N__39214\,
            lcout => n8_adj_1568,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i1_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__53438\,
            in1 => \N__39662\,
            in2 => \N__39563\,
            in3 => \N__49125\,
            lcout => \buf_cfgRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i1_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49123\,
            in1 => \N__39543\,
            in2 => \N__45635\,
            in3 => \N__39461\,
            lcout => \IAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__39197\,
            in1 => \N__55472\,
            in2 => \N__49242\,
            in3 => \N__39188\,
            lcout => \data_index_9_N_212_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6304_3_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41121\,
            in1 => \N__45616\,
            in2 => \_gnd_net_\,
            in3 => \N__39169\,
            lcout => n8_adj_1558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6374_3_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__53499\,
            in1 => \N__39355\,
            in2 => \_gnd_net_\,
            in3 => \N__41122\,
            lcout => n8_adj_1570,
            ltout => \n8_adj_1570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49103\,
            in1 => \N__55471\,
            in2 => \N__39330\,
            in3 => \N__39326\,
            lcout => \data_index_9_N_212_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i2_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55473\,
            in1 => \N__49108\,
            in2 => \N__39930\,
            in3 => \N__39915\,
            lcout => data_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i8_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__39198\,
            in1 => \N__55474\,
            in2 => \N__49243\,
            in3 => \N__39189\,
            lcout => data_index_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55470\,
            in1 => \N__49104\,
            in2 => \N__39929\,
            in3 => \N__39914\,
            lcout => \data_index_9_N_212_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imiso_83_12297_12298_set_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39812\,
            in1 => \N__39798\,
            in2 => \_gnd_net_\,
            in3 => \N__44323\,
            lcout => \comm_spi.n14818\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12297_12298_setC_net\,
            ce => 'H',
            sr => \N__42837\
        );

    \comm_spi.RESET_I_0_87_2_lut_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39786\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58158\,
            lcout => \comm_spi.DOUT_7__N_787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \wdtick_cnt_3763_3764__i1_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40321\,
            in1 => \N__39759\,
            in2 => \_gnd_net_\,
            in3 => \N__39747\,
            lcout => wdtick_cnt_0,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => n19932,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i2_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40313\,
            in1 => \N__39740\,
            in2 => \_gnd_net_\,
            in3 => \N__39726\,
            lcout => wdtick_cnt_1,
            ltout => OPEN,
            carryin => n19932,
            carryout => n19933,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i3_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40322\,
            in1 => \N__39723\,
            in2 => \_gnd_net_\,
            in3 => \N__39711\,
            lcout => wdtick_cnt_2,
            ltout => OPEN,
            carryin => n19933,
            carryout => n19934,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i4_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40314\,
            in1 => \N__39708\,
            in2 => \_gnd_net_\,
            in3 => \N__39696\,
            lcout => wdtick_cnt_3,
            ltout => OPEN,
            carryin => n19934,
            carryout => n19935,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i5_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40323\,
            in1 => \N__39693\,
            in2 => \_gnd_net_\,
            in3 => \N__39681\,
            lcout => wdtick_cnt_4,
            ltout => OPEN,
            carryin => n19935,
            carryout => n19936,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i6_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40315\,
            in1 => \N__39678\,
            in2 => \_gnd_net_\,
            in3 => \N__39666\,
            lcout => wdtick_cnt_5,
            ltout => OPEN,
            carryin => n19936,
            carryout => n19937,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i7_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__40073\,
            in2 => \_gnd_net_\,
            in3 => \N__40059\,
            lcout => wdtick_cnt_6,
            ltout => OPEN,
            carryin => n19937,
            carryout => n19938,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i8_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40316\,
            in1 => \N__40055\,
            in2 => \_gnd_net_\,
            in3 => \N__40041\,
            lcout => wdtick_cnt_7,
            ltout => OPEN,
            carryin => n19938,
            carryout => n19939,
            clk => \N__50785\,
            ce => \N__42635\,
            sr => \N__42153\
        );

    \wdtick_cnt_3763_3764__i9_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40308\,
            in1 => \N__40034\,
            in2 => \_gnd_net_\,
            in3 => \N__40020\,
            lcout => wdtick_cnt_8,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => n19940,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i10_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40326\,
            in1 => \N__40017\,
            in2 => \_gnd_net_\,
            in3 => \N__40005\,
            lcout => wdtick_cnt_9,
            ltout => OPEN,
            carryin => n19940,
            carryout => n19941,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i11_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40305\,
            in1 => \N__39998\,
            in2 => \_gnd_net_\,
            in3 => \N__39984\,
            lcout => wdtick_cnt_10,
            ltout => OPEN,
            carryin => n19941,
            carryout => n19942,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i12_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40327\,
            in1 => \N__39981\,
            in2 => \_gnd_net_\,
            in3 => \N__39969\,
            lcout => wdtick_cnt_11,
            ltout => OPEN,
            carryin => n19942,
            carryout => n19943,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i13_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40306\,
            in1 => \N__39962\,
            in2 => \_gnd_net_\,
            in3 => \N__39948\,
            lcout => wdtick_cnt_12,
            ltout => OPEN,
            carryin => n19943,
            carryout => n19944,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i14_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40328\,
            in1 => \N__39945\,
            in2 => \_gnd_net_\,
            in3 => \N__39933\,
            lcout => wdtick_cnt_13,
            ltout => OPEN,
            carryin => n19944,
            carryout => n19945,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i15_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40307\,
            in1 => \N__40212\,
            in2 => \_gnd_net_\,
            in3 => \N__40197\,
            lcout => wdtick_cnt_14,
            ltout => OPEN,
            carryin => n19945,
            carryout => n19946,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i16_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40329\,
            in1 => \N__40194\,
            in2 => \_gnd_net_\,
            in3 => \N__40182\,
            lcout => wdtick_cnt_15,
            ltout => OPEN,
            carryin => n19946,
            carryout => n19947,
            clk => \N__50787\,
            ce => \N__42631\,
            sr => \N__42147\
        );

    \wdtick_cnt_3763_3764__i17_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40317\,
            in1 => \N__40179\,
            in2 => \_gnd_net_\,
            in3 => \N__40167\,
            lcout => wdtick_cnt_16,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => n19948,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i18_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40309\,
            in1 => \N__40164\,
            in2 => \_gnd_net_\,
            in3 => \N__40152\,
            lcout => wdtick_cnt_17,
            ltout => OPEN,
            carryin => n19948,
            carryout => n19949,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i19_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40318\,
            in1 => \N__40148\,
            in2 => \_gnd_net_\,
            in3 => \N__40134\,
            lcout => wdtick_cnt_18,
            ltout => OPEN,
            carryin => n19949,
            carryout => n19950,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i20_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40310\,
            in1 => \N__40130\,
            in2 => \_gnd_net_\,
            in3 => \N__40116\,
            lcout => wdtick_cnt_19,
            ltout => OPEN,
            carryin => n19950,
            carryout => n19951,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i21_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40319\,
            in1 => \N__40112\,
            in2 => \_gnd_net_\,
            in3 => \N__40098\,
            lcout => wdtick_cnt_20,
            ltout => OPEN,
            carryin => n19951,
            carryout => n19952,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i22_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40311\,
            in1 => \N__40095\,
            in2 => \_gnd_net_\,
            in3 => \N__40083\,
            lcout => wdtick_cnt_21,
            ltout => OPEN,
            carryin => n19952,
            carryout => n19953,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i23_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40320\,
            in1 => \N__40359\,
            in2 => \_gnd_net_\,
            in3 => \N__40347\,
            lcout => wdtick_cnt_22,
            ltout => OPEN,
            carryin => n19953,
            carryout => n19954,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i24_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__40312\,
            in1 => \N__40344\,
            in2 => \_gnd_net_\,
            in3 => \N__40332\,
            lcout => wdtick_cnt_23,
            ltout => OPEN,
            carryin => n19954,
            carryout => n19955,
            clk => \N__50789\,
            ce => \N__42630\,
            sr => \N__42143\
        );

    \wdtick_cnt_3763_3764__i25_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__40226\,
            in1 => \N__40325\,
            in2 => \_gnd_net_\,
            in3 => \N__40230\,
            lcout => wdtick_cnt_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50790\,
            ce => \N__42636\,
            sr => \N__42152\
        );

    \comm_spi.data_rx_i7_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__53160\,
            in1 => \N__42781\,
            in2 => \_gnd_net_\,
            in3 => \N__42746\,
            lcout => comm_rx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \comm_spi.data_rx_i6_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__42745\,
            in1 => \N__53291\,
            in2 => \N__42797\,
            in3 => \_gnd_net_\,
            lcout => comm_rx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \comm_spi.data_rx_i5_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__53584\,
            in1 => \N__42780\,
            in2 => \_gnd_net_\,
            in3 => \N__42744\,
            lcout => comm_rx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \comm_spi.data_rx_i4_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__42743\,
            in1 => \N__49810\,
            in2 => \N__42796\,
            in3 => \_gnd_net_\,
            lcout => comm_rx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \comm_spi.data_rx_i3_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__50094\,
            in1 => \N__42779\,
            in2 => \_gnd_net_\,
            in3 => \N__42742\,
            lcout => comm_rx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \comm_spi.data_rx_i2_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__42741\,
            in1 => \_gnd_net_\,
            in2 => \N__42795\,
            in3 => \N__49659\,
            lcout => comm_rx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \comm_spi.data_rx_i1_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__48677\,
            in1 => \N__42778\,
            in2 => \_gnd_net_\,
            in3 => \N__42740\,
            lcout => comm_rx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58402\,
            ce => 'H',
            sr => \N__58145\
        );

    \clk_RTD_287_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40473\,
            in1 => \N__45000\,
            in2 => \_gnd_net_\,
            in3 => \N__44976\,
            lcout => \clk_RTD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19121_2_lut_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__53965\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48188\,
            lcout => n21588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19054_2_lut_3_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__46036\,
            in1 => \N__52762\,
            in2 => \_gnd_net_\,
            in3 => \N__53964\,
            lcout => n21586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12442_2_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43305\,
            lcout => n14958,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15473_2_lut_3_lut_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__54754\,
            in1 => \N__45620\,
            in2 => \_gnd_net_\,
            in3 => \N__54367\,
            lcout => n14_adj_1550,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18549_4_lut_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__42471\,
            in1 => \N__52382\,
            in2 => \N__53070\,
            in3 => \N__43559\,
            lcout => n21276,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_250_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__54753\,
            in1 => \N__54366\,
            in2 => \_gnd_net_\,
            in3 => \N__55067\,
            lcout => n12433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22461_bdd_4_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__40422\,
            in1 => \N__40413\,
            in2 => \N__40401\,
            in3 => \N__47530\,
            lcout => n22464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19172_2_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40383\,
            in2 => \_gnd_net_\,
            in3 => \N__57179\,
            lcout => OPEN,
            ltout => \n21556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19770_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__42168\,
            in1 => \N__46471\,
            in2 => \N__40779\,
            in3 => \N__47529\,
            lcout => n22521,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22521_bdd_4_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__40776\,
            in1 => \N__40764\,
            in2 => \N__41478\,
            in3 => \N__47531\,
            lcout => OPEN,
            ltout => \n22524_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1565241_i1_3_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40758\,
            in2 => \N__40752\,
            in3 => \N__47163\,
            lcout => OPEN,
            ltout => \n30_adj_1676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i4_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__53600\,
            in1 => \_gnd_net_\,
            in2 => \N__40749\,
            in3 => \N__54401\,
            lcout => comm_buf_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55980\,
            ce => \N__43326\,
            sr => \N__43250\
        );

    \n22485_bdd_4_lut_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__40746\,
            in1 => \N__47691\,
            in2 => \N__40731\,
            in3 => \N__40716\,
            lcout => n22488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i26_3_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40704\,
            in1 => \N__57114\,
            in2 => \_gnd_net_\,
            in3 => \N__40682\,
            lcout => OPEN,
            ltout => \n26_adj_1687_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19716_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__52590\,
            in1 => \N__47692\,
            in2 => \N__40656\,
            in3 => \N__46485\,
            lcout => OPEN,
            ltout => \n22455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22455_bdd_4_lut_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47693\,
            in1 => \N__45699\,
            in2 => \N__40653\,
            in3 => \N__40650\,
            lcout => OPEN,
            ltout => \n22458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1564035_i1_3_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40632\,
            in2 => \N__40626\,
            in3 => \N__47268\,
            lcout => OPEN,
            ltout => \n30_adj_1688_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i2_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__50108\,
            in1 => \_gnd_net_\,
            in2 => \N__40932\,
            in3 => \N__54402\,
            lcout => comm_buf_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55993\,
            ce => \N__43336\,
            sr => \N__43264\
        );

    \mux_128_Mux_0_i26_3_lut_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40929\,
            in1 => \N__57109\,
            in2 => \_gnd_net_\,
            in3 => \N__40897\,
            lcout => OPEN,
            ltout => \n26_adj_1533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18519_4_lut_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__57110\,
            in1 => \N__40881\,
            in2 => \N__40866\,
            in3 => \N__46409\,
            lcout => OPEN,
            ltout => \n21246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19828_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__47250\,
            in1 => \N__40863\,
            in2 => \N__40854\,
            in3 => \N__47710\,
            lcout => OPEN,
            ltout => \n22581_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22581_bdd_4_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__40851\,
            in1 => \N__40839\,
            in2 => \N__40824\,
            in3 => \N__47251\,
            lcout => OPEN,
            ltout => \n22584_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i0_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54400\,
            in1 => \_gnd_net_\,
            in2 => \N__40821\,
            in3 => \N__48676\,
            lcout => comm_buf_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56007\,
            ce => \N__43337\,
            sr => \N__43263\
        );

    \i19282_4_lut_4_lut_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111011110011"
        )
    port map (
            in0 => \N__47709\,
            in1 => \N__46408\,
            in2 => \N__57217\,
            in3 => \N__47249\,
            lcout => n21479,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i3_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54556\,
            in1 => \N__49860\,
            in2 => \_gnd_net_\,
            in3 => \N__41250\,
            lcout => comm_buf_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56023\,
            ce => \N__45199\,
            sr => \N__44009\
        );

    \comm_cmd_1__bdd_4_lut_19862_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__47663\,
            in1 => \N__40818\,
            in2 => \N__40794\,
            in3 => \N__46479\,
            lcout => OPEN,
            ltout => \n22623_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22623_bdd_4_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__41304\,
            in1 => \N__41265\,
            in2 => \N__41256\,
            in3 => \N__47664\,
            lcout => OPEN,
            ltout => \n22626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1568859_i1_3_lut_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47255\,
            in2 => \N__41253\,
            in3 => \N__41148\,
            lcout => n30_adj_1643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_3_i26_3_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41244\,
            in1 => \N__57128\,
            in2 => \_gnd_net_\,
            in3 => \N__41215\,
            lcout => OPEN,
            ltout => \n26_adj_1642_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19692_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__47661\,
            in1 => \N__56601\,
            in2 => \N__41199\,
            in3 => \N__46478\,
            lcout => OPEN,
            ltout => \n22425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22425_bdd_4_lut_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__41196\,
            in1 => \N__47662\,
            in2 => \N__41172\,
            in3 => \N__41169\,
            lcout => n22428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i0_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__41052\,
            in1 => \N__41046\,
            in2 => \N__49331\,
            in3 => \N__55288\,
            lcout => data_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4379_3_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45669\,
            in1 => \N__41142\,
            in2 => \_gnd_net_\,
            in3 => \N__41123\,
            lcout => n8_adj_1540,
            ltout => \n8_adj_1540_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__49234\,
            in1 => \N__41045\,
            in2 => \N__41037\,
            in3 => \N__55287\,
            lcout => \data_index_9_N_212_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i4_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__47774\,
            in1 => \N__49235\,
            in2 => \N__42009\,
            in3 => \N__41497\,
            lcout => \VDC_RNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i0_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__41723\,
            in1 => \N__45670\,
            in2 => \N__46917\,
            in3 => \N__46745\,
            lcout => buf_dds1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_0_i16_3_lut_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57113\,
            in1 => \N__41530\,
            in2 => \_gnd_net_\,
            in3 => \N__41722\,
            lcout => OPEN,
            ltout => \n16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18530_3_lut_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46376\,
            in2 => \N__41709\,
            in3 => \N__41705\,
            lcout => n21257,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i0_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__43194\,
            in1 => \N__41531\,
            in2 => \_gnd_net_\,
            in3 => \N__41637\,
            lcout => buf_dds0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i23_3_lut_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57111\,
            in2 => \N__41501\,
            in3 => \N__50649\,
            lcout => n23_adj_1675,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i16_3_lut_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46958\,
            in1 => \N__41455\,
            in2 => \_gnd_net_\,
            in3 => \N__57112\,
            lcout => n16_adj_1624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4272_2_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54827\,
            in2 => \_gnd_net_\,
            in3 => \N__54380\,
            lcout => n9342,
            ltout => \n9342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15206_4_lut_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__55286\,
            in1 => \N__41438\,
            in2 => \N__41427\,
            in3 => \N__41417\,
            lcout => \data_index_9_N_212_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18635_3_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46477\,
            in1 => \N__42050\,
            in2 => \_gnd_net_\,
            in3 => \N__42021\,
            lcout => n21362,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i6_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49062\,
            in1 => \N__42008\,
            in2 => \N__49585\,
            in3 => \N__50710\,
            lcout => buf_control_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.CS_28_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__44669\,
            in1 => \N__44726\,
            in2 => \_gnd_net_\,
            in3 => \N__44388\,
            lcout => \DDS_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56080\,
            ce => \N__41934\,
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__41915\,
            in1 => \N__49112\,
            in2 => \N__55463\,
            in3 => \N__41904\,
            lcout => \data_index_9_N_212_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.MISO_48_12291_12292_reset_LC_16_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41799\,
            in1 => \N__41783\,
            in2 => \_gnd_net_\,
            in3 => \N__44313\,
            lcout => \comm_spi.n14813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12291_12292_resetC_net\,
            ce => 'H',
            sr => \N__42880\
        );

    \comm_spi.MISO_48_12291_12292_set_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41798\,
            in1 => \N__41787\,
            in2 => \_gnd_net_\,
            in3 => \N__44312\,
            lcout => \comm_spi.n14812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12291_12292_setC_net\,
            ce => 'H',
            sr => \N__42829\
        );

    \i19344_2_lut_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41769\,
            in2 => \_gnd_net_\,
            in3 => \N__57272\,
            lcout => n21672,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19397_2_lut_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__51753\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51493\,
            lcout => OPEN,
            ltout => \ADC_VDC.n22124_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.SCLK_46_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__42446\,
            in1 => \N__44262\,
            in2 => \N__41739\,
            in3 => \N__51208\,
            lcout => \VDC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__42363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19347_2_lut_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42183\,
            in2 => \_gnd_net_\,
            in3 => \N__57270\,
            lcout => n21557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \flagcntwd_303_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__53979\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54486\,
            lcout => flagcntwd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55945\,
            ce => \N__42099\,
            sr => \N__42083\
        );

    \i18460_2_lut_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54379\,
            in2 => \_gnd_net_\,
            in3 => \N__53978\,
            lcout => OPEN,
            ltout => \n21187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_277_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__55238\,
            in1 => \N__54862\,
            in2 => \N__42102\,
            in3 => \N__55572\,
            lcout => n11605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_186_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__54859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55235\,
            lcout => n80,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_56_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__55236\,
            in1 => \_gnd_net_\,
            in2 => \N__54502\,
            in3 => \N__54861\,
            lcout => n20578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_243_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__54860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53977\,
            lcout => OPEN,
            ltout => \n11576_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_289_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__55237\,
            in1 => \N__54485\,
            in2 => \N__42072\,
            in3 => \N__55571\,
            lcout => n12148,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_45_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__54858\,
            in1 => \N__54375\,
            in2 => \_gnd_net_\,
            in3 => \N__55234\,
            lcout => n21143,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i4_12317_12318_set_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56504\,
            in1 => \N__56487\,
            in2 => \_gnd_net_\,
            in3 => \N__57378\,
            lcout => \comm_spi.n14838\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58337\,
            ce => 'H',
            sr => \N__56421\
        );

    \i12470_2_lut_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55251\,
            in2 => \_gnd_net_\,
            in3 => \N__45059\,
            lcout => n14986,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12477_2_lut_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__48293\,
            in1 => \_gnd_net_\,
            in2 => \N__55358\,
            in3 => \_gnd_net_\,
            lcout => n14993,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9391_1_lut_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44822\,
            lcout => n11910,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15273_2_lut_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44992\,
            in2 => \_gnd_net_\,
            in3 => \N__44967\,
            lcout => n17773,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19029_2_lut_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__57271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42588\,
            lcout => n21385,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22539_bdd_4_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__43215\,
            in1 => \N__44071\,
            in2 => \N__42550\,
            in3 => \N__52447\,
            lcout => OPEN,
            ltout => \n22542_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i7_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__52555\,
            in1 => \N__42483\,
            in2 => \N__42474\,
            in3 => \_gnd_net_\,
            lcout => comm_tx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55960\,
            ce => \N__50341\,
            sr => \N__50261\
        );

    \mux_137_Mux_7_i4_3_lut_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48048\,
            in1 => \N__44907\,
            in2 => \_gnd_net_\,
            in3 => \N__53073\,
            lcout => n4_adj_1580,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19490_4_lut_3_lut_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__44311\,
            in1 => \N__42847\,
            in2 => \N__58156\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_100_2_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__42852\,
            in3 => \N__58108\,
            lcout => \comm_spi.data_tx_7__N_814\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_92_2_lut_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__58109\,
            in1 => \N__42851\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_806\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_valid_85_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__42801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42750\,
            lcout => comm_data_vld,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.data_valid_85C_net\,
            ce => 'H',
            sr => \N__58122\
        );

    \comm_index_0__bdd_4_lut_19794_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__53047\,
            in1 => \N__49890\,
            in2 => \N__45975\,
            in3 => \N__52379\,
            lcout => OPEN,
            ltout => \n22551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22551_bdd_4_lut_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52380\,
            in1 => \N__47759\,
            in2 => \N__42717\,
            in3 => \N__42709\,
            lcout => n22554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_4_i4_3_lut_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53048\,
            in1 => \N__47985\,
            in2 => \_gnd_net_\,
            in3 => \N__44856\,
            lcout => OPEN,
            ltout => \n4_adj_1582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18558_4_lut_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__52381\,
            in1 => \N__53556\,
            in2 => \N__42648\,
            in3 => \N__53049\,
            lcout => OPEN,
            ltout => \n21285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i4_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__52523\,
            in1 => \_gnd_net_\,
            in2 => \N__42645\,
            in3 => \N__42642\,
            lcout => comm_tx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55981\,
            ce => \N__50334\,
            sr => \N__50243\
        );

    \i19295_2_lut_3_lut_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__52378\,
            in1 => \N__52522\,
            in2 => \_gnd_net_\,
            in3 => \N__49932\,
            lcout => OPEN,
            ltout => \n21474_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_290_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110011"
        )
    port map (
            in0 => \N__53046\,
            in1 => \N__54374\,
            in2 => \N__43113\,
            in3 => \N__48241\,
            lcout => OPEN,
            ltout => \n12_adj_1596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_291_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48411\,
            in2 => \N__43110\,
            in3 => \N__48749\,
            lcout => n12184,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_1_i26_3_lut_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43107\,
            in1 => \N__57162\,
            in2 => \_gnd_net_\,
            in3 => \N__43085\,
            lcout => OPEN,
            ltout => \n26_adj_1694_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18633_4_lut_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__43059\,
            in1 => \N__57180\,
            in2 => \N__43050\,
            in3 => \N__46472\,
            lcout => n21360,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19852_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__46473\,
            in1 => \N__43047\,
            in2 => \N__57258\,
            in3 => \N__43002\,
            lcout => OPEN,
            ltout => \n22617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22617_bdd_4_lut_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__42981\,
            in1 => \N__42953\,
            in2 => \N__42918\,
            in3 => \N__46474\,
            lcout => OPEN,
            ltout => \n22620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18634_3_lut_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47517\,
            in1 => \_gnd_net_\,
            in2 => \N__42915\,
            in3 => \N__42912\,
            lcout => OPEN,
            ltout => \n21361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1563432_i1_3_lut_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42906\,
            in2 => \N__42891\,
            in3 => \N__47154\,
            lcout => OPEN,
            ltout => \n30_adj_1695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i1_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54484\,
            in1 => \_gnd_net_\,
            in2 => \N__43341\,
            in3 => \N__49678\,
            lcout => comm_buf_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55994\,
            ce => \N__43324\,
            sr => \N__43274\
        );

    \i41_4_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100100100000"
        )
    port map (
            in0 => \N__46470\,
            in1 => \N__47153\,
            in2 => \N__57249\,
            in3 => \N__47516\,
            lcout => n24_adj_1639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19784_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__45507\,
            in1 => \N__52445\,
            in2 => \N__48510\,
            in3 => \N__53066\,
            lcout => n22539,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15538_2_lut_3_lut_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45677\,
            in1 => \N__54777\,
            in2 => \_gnd_net_\,
            in3 => \N__54438\,
            lcout => n14_adj_1541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_4_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001000"
        )
    port map (
            in0 => \N__54437\,
            in1 => \N__55247\,
            in2 => \N__54842\,
            in3 => \N__53962\,
            lcout => n12541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i30_3_lut_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47254\,
            in1 => \N__43152\,
            in2 => \_gnd_net_\,
            in3 => \N__43137\,
            lcout => n30_adj_1531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_3_i7_4_lut_4_lut_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111100110"
        )
    port map (
            in0 => \N__54439\,
            in1 => \N__54787\,
            in2 => \N__43125\,
            in3 => \N__53963\,
            lcout => n18070,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12449_2_lut_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__45170\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55249\,
            lcout => n14965,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12456_2_lut_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55250\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45902\,
            lcout => n14972,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i7_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__55248\,
            in1 => \N__48588\,
            in2 => \N__43560\,
            in3 => \N__53142\,
            lcout => comm_buf_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56008\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22515_bdd_4_lut_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011000010"
        )
    port map (
            in0 => \N__43542\,
            in1 => \N__43410\,
            in2 => \N__47728\,
            in3 => \N__43518\,
            lcout => n22518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19804_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__43497\,
            in1 => \N__46484\,
            in2 => \N__43488\,
            in3 => \N__47712\,
            lcout => n22527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i26_3_lut_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43461\,
            in1 => \N__57250\,
            in2 => \_gnd_net_\,
            in3 => \N__43432\,
            lcout => OPEN,
            ltout => \n26_adj_1626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19765_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__53244\,
            in1 => \N__46483\,
            in2 => \N__43413\,
            in3 => \N__47711\,
            lcout => n22515,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22527_bdd_4_lut_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__47716\,
            in1 => \N__43404\,
            in2 => \N__43388\,
            in3 => \N__43359\,
            lcout => OPEN,
            ltout => \n22530_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1570668_i1_3_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47256\,
            in2 => \N__43353\,
            in3 => \N__43350\,
            lcout => OPEN,
            ltout => \n30_adj_1627_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i6_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53217\,
            in2 => \N__43344\,
            in3 => \N__54542\,
            lcout => comm_buf_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56024\,
            ce => \N__45209\,
            sr => \N__43962\
        );

    \mux_129_Mux_0_i26_3_lut_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43869\,
            in1 => \N__57130\,
            in2 => \_gnd_net_\,
            in3 => \N__43845\,
            lcout => OPEN,
            ltout => \n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18534_4_lut_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__46482\,
            in1 => \N__43818\,
            in2 => \N__43803\,
            in3 => \N__57131\,
            lcout => OPEN,
            ltout => \n21261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19814_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__43626\,
            in1 => \N__47196\,
            in2 => \N__43800\,
            in3 => \N__47717\,
            lcout => OPEN,
            ltout => \n22563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22563_bdd_4_lut_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__43683\,
            in1 => \N__47257\,
            in2 => \N__43797\,
            in3 => \N__43794\,
            lcout => OPEN,
            ltout => \n22566_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i0_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48697\,
            in2 => \N__43785\,
            in3 => \N__54543\,
            lcout => comm_buf_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56039\,
            ce => \N__45194\,
            sr => \N__44001\
        );

    \mux_129_Mux_0_i19_3_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__57129\,
            in1 => \N__43782\,
            in2 => \N__43757\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18531_3_lut_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__43710\,
            in1 => \_gnd_net_\,
            in2 => \N__43686\,
            in3 => \N__46481\,
            lcout => n21258,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18533_3_lut_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46480\,
            in1 => \N__43677\,
            in2 => \_gnd_net_\,
            in3 => \N__43656\,
            lcout => n21260,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22431_bdd_4_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__47722\,
            in1 => \N__43613\,
            in2 => \N__43587\,
            in3 => \N__43575\,
            lcout => n22434,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i26_3_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44217\,
            in1 => \N__57251\,
            in2 => \_gnd_net_\,
            in3 => \N__44199\,
            lcout => OPEN,
            ltout => \n26_adj_1653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19755_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__46476\,
            in1 => \N__57291\,
            in2 => \N__44175\,
            in3 => \N__47723\,
            lcout => OPEN,
            ltout => \n22497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22497_bdd_4_lut_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47724\,
            in1 => \N__44172\,
            in2 => \N__44151\,
            in3 => \N__44148\,
            lcout => OPEN,
            ltout => \n22500_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1567653_i1_3_lut_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44127\,
            in2 => \N__44121\,
            in3 => \N__47253\,
            lcout => OPEN,
            ltout => \n30_adj_1654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i1_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54541\,
            in2 => \N__44118\,
            in3 => \N__49722\,
            lcout => comm_buf_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56055\,
            ce => \N__45211\,
            sr => \N__44014\
        );

    \i1_2_lut_4_lut_adj_230_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__46475\,
            in1 => \N__47252\,
            in2 => \N__44115\,
            in3 => \N__47721\,
            lcout => n68,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i7_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54567\,
            in1 => \N__48599\,
            in2 => \_gnd_net_\,
            in3 => \N__46971\,
            lcout => comm_buf_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56067\,
            ce => \N__45210\,
            sr => \N__44013\
        );

    \SIG_DDS.i19394_4_lut_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100110"
        )
    port map (
            in0 => \N__44657\,
            in1 => \N__44748\,
            in2 => \N__43943\,
            in3 => \N__44376\,
            lcout => \SIG_DDS.n12895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15221_2_lut_2_lut_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__44829\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44799\,
            lcout => \CONT_SD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i1_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44754\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44668\,
            lcout => dds_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56087\,
            ce => \N__44543\,
            sr => \N__44503\
        );

    \comm_spi.i12293_3_lut_LC_17_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44343\,
            in1 => \N__44337\,
            in2 => \_gnd_net_\,
            in3 => \N__44330\,
            lcout => \ICE_SPI_MISO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19395_4_lut_4_lut_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111001"
        )
    port map (
            in0 => \N__51492\,
            in1 => \N__51895\,
            in2 => \N__51761\,
            in3 => \N__51213\,
            lcout => \ADC_VDC.n11895\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19480_4_lut_3_lut_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44256\,
            in1 => \N__48140\,
            in2 => \_gnd_net_\,
            in3 => \N__58159\,
            lcout => \comm_spi.n23086\,
            ltout => \comm_spi.n23086_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12285_3_lut_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__46653\,
            in1 => \N__44247\,
            in2 => \N__44250\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.iclk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12283_12284_set_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48141\,
            lcout => \comm_spi.n14804\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55946\,
            ce => 'H',
            sr => \N__46647\
        );

    \i19131_4_lut_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__44241\,
            in1 => \N__47270\,
            in2 => \N__44235\,
            in3 => \N__47642\,
            lcout => n21481,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19510_4_lut_3_lut_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__56503\,
            in1 => \N__56140\,
            in2 => \_gnd_net_\,
            in3 => \N__57988\,
            lcout => \comm_spi.n23101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19485_4_lut_3_lut_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45016\,
            in1 => \N__50869\,
            in2 => \_gnd_net_\,
            in3 => \N__57987\,
            lcout => \comm_spi.n23092\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_cnt_3761_3762__i2_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__44969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44993\,
            lcout => clk_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50791\,
            ce => 'H',
            sr => \N__44949\
        );

    \clk_cnt_3761_3762__i1_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44968\,
            lcout => clk_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__50791\,
            ce => 'H',
            sr => \N__44949\
        );

    \comm_buf_4__i0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44940\,
            in1 => \N__54335\,
            in2 => \_gnd_net_\,
            in3 => \N__48703\,
            lcout => comm_buf_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i7_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54334\,
            in1 => \_gnd_net_\,
            in2 => \N__48596\,
            in3 => \N__44922\,
            lcout => comm_buf_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i6_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53227\,
            in1 => \N__44901\,
            in2 => \_gnd_net_\,
            in3 => \N__54338\,
            lcout => comm_buf_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i5_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54333\,
            in1 => \N__53331\,
            in2 => \_gnd_net_\,
            in3 => \N__44889\,
            lcout => comm_buf_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i4_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53619\,
            in1 => \N__44874\,
            in2 => \_gnd_net_\,
            in3 => \N__54337\,
            lcout => comm_buf_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i3_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54332\,
            in1 => \N__49867\,
            in2 => \_gnd_net_\,
            in3 => \N__44847\,
            lcout => comm_buf_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i2_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50145\,
            in1 => \N__45126\,
            in2 => \_gnd_net_\,
            in3 => \N__54336\,
            lcout => comm_buf_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \comm_buf_4__i1_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54331\,
            in1 => \N__49717\,
            in2 => \_gnd_net_\,
            in3 => \N__45108\,
            lcout => comm_buf_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55970\,
            ce => \N__45060\,
            sr => \N__45090\
        );

    \i18541_4_lut_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__52151\,
            in1 => \N__45075\,
            in2 => \N__45069\,
            in3 => \N__54841\,
            lcout => OPEN,
            ltout => \n21268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i0_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49374\,
            in2 => \N__45078\,
            in3 => \N__55066\,
            lcout => comm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55982\,
            ce => \N__48453\,
            sr => \_gnd_net_\
        );

    \i19367_3_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__50003\,
            in1 => \N__46037\,
            in2 => \_gnd_net_\,
            in3 => \N__54191\,
            lcout => n22094,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18539_3_lut_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011101"
        )
    port map (
            in0 => \N__54192\,
            in1 => \N__52782\,
            in2 => \_gnd_net_\,
            in3 => \N__53869\,
            lcout => n21266,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_301_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__48764\,
            in1 => \N__53071\,
            in2 => \N__45390\,
            in3 => \N__45039\,
            lcout => n12407,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_304_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__52783\,
            in1 => \N__50002\,
            in2 => \N__52855\,
            in3 => \N__53868\,
            lcout => n21085,
            ltout => \n21085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_262_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__52446\,
            in1 => \_gnd_net_\,
            in2 => \N__45042\,
            in3 => \N__52553\,
            lcout => n19188,
            ltout => \n19188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_309_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__53072\,
            in1 => \N__45388\,
            in2 => \N__45360\,
            in3 => \N__48765\,
            lcout => n12431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__52990\,
            in1 => \N__45948\,
            in2 => \N__49776\,
            in3 => \N__52409\,
            lcout => OPEN,
            ltout => \n22557_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22557_bdd_4_lut_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52410\,
            in1 => \N__45334\,
            in2 => \N__45285\,
            in3 => \N__45280\,
            lcout => n22560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_3_i4_3_lut_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__52991\,
            in1 => \_gnd_net_\,
            in2 => \N__47961\,
            in3 => \N__45252\,
            lcout => OPEN,
            ltout => \n4_adj_1583_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18561_4_lut_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__52411\,
            in1 => \N__46620\,
            in2 => \N__45243\,
            in3 => \N__52992\,
            lcout => OPEN,
            ltout => \n21288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i3_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45240\,
            in2 => \N__45234\,
            in3 => \N__52521\,
            lcout => comm_tx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55995\,
            ce => \N__50333\,
            sr => \N__50254\
        );

    \i19129_3_lut_4_lut_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__52520\,
            in1 => \N__52989\,
            in2 => \N__52439\,
            in3 => \N__49931\,
            lcout => OPEN,
            ltout => \n21477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i48_4_lut_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__45231\,
            in1 => \N__54440\,
            in2 => \N__45219\,
            in3 => \N__48257\,
            lcout => OPEN,
            ltout => \n44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_294_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48409\,
            in2 => \N__45216\,
            in3 => \N__48742\,
            lcout => n12260,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_2_i1_3_lut_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45829\,
            in1 => \N__45475\,
            in2 => \_gnd_net_\,
            in3 => \N__53065\,
            lcout => OPEN,
            ltout => \n1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i2_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__52560\,
            in1 => \N__45420\,
            in2 => \N__45423\,
            in3 => \N__45396\,
            lcout => comm_tx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56009\,
            ce => \N__50355\,
            sr => \N__50265\
        );

    \i19154_2_lut_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__50072\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53062\,
            lcout => n21528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_2_i2_3_lut_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53064\,
            in1 => \_gnd_net_\,
            in2 => \N__49755\,
            in3 => \N__45927\,
            lcout => n2_adj_1584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_2_i4_3_lut_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47937\,
            in1 => \N__45414\,
            in2 => \_gnd_net_\,
            in3 => \N__53063\,
            lcout => OPEN,
            ltout => \n4_adj_1585_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__52559\,
            in1 => \N__45405\,
            in2 => \N__45399\,
            in3 => \N__52444\,
            lcout => n22491,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_281_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__52443\,
            in1 => \N__52558\,
            in2 => \_gnd_net_\,
            in3 => \N__49943\,
            lcout => OPEN,
            ltout => \n19193_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_299_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__53061\,
            in1 => \N__45389\,
            in2 => \N__45363\,
            in3 => \N__48763\,
            lcout => n12353,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45687\,
            in1 => \N__45549\,
            in2 => \_gnd_net_\,
            in3 => \N__52557\,
            lcout => comm_tx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56025\,
            ce => \N__50305\,
            sr => \N__50231\
        );

    \i18546_4_lut_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__52434\,
            in1 => \N__50037\,
            in2 => \N__46641\,
            in3 => \N__53052\,
            lcout => n21273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19779_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__53051\,
            in1 => \N__45525\,
            in2 => \N__48624\,
            in3 => \N__52432\,
            lcout => OPEN,
            ltout => \n22533_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22533_bdd_4_lut_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__52433\,
            in1 => \N__45681\,
            in2 => \N__45651\,
            in3 => \N__45621\,
            lcout => n22536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19137_3_lut_4_lut_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__52556\,
            in1 => \N__53050\,
            in2 => \N__52448\,
            in3 => \N__49942\,
            lcout => OPEN,
            ltout => \n21497_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i39_4_lut_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__45543\,
            in1 => \N__54525\,
            in2 => \N__45537\,
            in3 => \N__48258\,
            lcout => OPEN,
            ltout => \n34_adj_1649_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_296_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__48750\,
            in1 => \_gnd_net_\,
            in2 => \N__45534\,
            in3 => \N__48410\,
            lcout => n12314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i0_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48699\,
            in1 => \N__45531\,
            in2 => \_gnd_net_\,
            in3 => \N__54548\,
            lcout => comm_buf_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i7_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54547\,
            in1 => \N__48595\,
            in2 => \_gnd_net_\,
            in3 => \N__45519\,
            lcout => comm_buf_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i6_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45501\,
            in1 => \N__54551\,
            in2 => \_gnd_net_\,
            in3 => \N__53218\,
            lcout => comm_buf_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i5_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54546\,
            in1 => \_gnd_net_\,
            in2 => \N__53345\,
            in3 => \N__46005\,
            lcout => comm_buf_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i4_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45990\,
            in1 => \N__53649\,
            in2 => \_gnd_net_\,
            in3 => \N__54550\,
            lcout => comm_buf_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i3_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54545\,
            in1 => \N__49868\,
            in2 => \_gnd_net_\,
            in3 => \N__45963\,
            lcout => comm_buf_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i2_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50165\,
            in1 => \N__45939\,
            in2 => \_gnd_net_\,
            in3 => \N__54549\,
            lcout => comm_buf_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \comm_buf_2__i1_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54544\,
            in1 => \N__49723\,
            in2 => \_gnd_net_\,
            in3 => \N__45918\,
            lcout => comm_buf_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56040\,
            ce => \N__45906\,
            sr => \N__45891\
        );

    \i1_2_lut_3_lut_adj_57_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__52090\,
            in1 => \N__54847\,
            in2 => \_gnd_net_\,
            in3 => \N__55270\,
            lcout => n16824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i10_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49310\,
            in1 => \N__47920\,
            in2 => \N__45864\,
            in3 => \N__50607\,
            lcout => \acadc_skipCount_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56056\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19161_2_lut_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45768\,
            in2 => \_gnd_net_\,
            in3 => \N__57210\,
            lcout => n21543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_2_i23_3_lut_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57211\,
            in1 => \N__45728\,
            in2 => \_gnd_net_\,
            in3 => \N__50606\,
            lcout => n23_adj_1685,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i0_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__55271\,
            in1 => \N__48698\,
            in2 => \N__46640\,
            in3 => \N__53128\,
            lcout => comm_buf_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56056\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i3_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__53129\,
            in1 => \N__46616\,
            in2 => \N__55388\,
            in3 => \N__49877\,
            lcout => comm_buf_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56056\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18641_3_lut_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46372\,
            in1 => \N__46602\,
            in2 => \_gnd_net_\,
            in3 => \N__46578\,
            lcout => n21368,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i26_3_lut_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46551\,
            in1 => \N__57252\,
            in2 => \_gnd_net_\,
            in3 => \N__46526\,
            lcout => OPEN,
            ltout => \n26_adj_1622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18642_4_lut_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__57253\,
            in1 => \N__46500\,
            in2 => \N__46488\,
            in3 => \N__46373\,
            lcout => n21369,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i0_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101000110110"
        )
    port map (
            in0 => \N__46374\,
            in1 => \N__47195\,
            in2 => \N__47708\,
            in3 => \N__57257\,
            lcout => comm_length_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56068\,
            ce => \N__52095\,
            sr => \N__46059\
        );

    \comm_length_i1_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101101011111101"
        )
    port map (
            in0 => \N__47194\,
            in1 => \N__47638\,
            in2 => \N__57273\,
            in3 => \N__46375\,
            lcout => comm_length_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56068\,
            ce => \N__52095\,
            sr => \N__46059\
        );

    \i2_3_lut_adj_298_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__46047\,
            in1 => \N__52449\,
            in2 => \_gnd_net_\,
            in3 => \N__48429\,
            lcout => n5_adj_1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i12_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__49309\,
            in1 => \N__47925\,
            in2 => \N__47815\,
            in3 => \N__50648\,
            lcout => \acadc_skipCount_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__47262\,
            in1 => \N__47637\,
            in2 => \N__47316\,
            in3 => \N__47307\,
            lcout => OPEN,
            ltout => \n22599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22599_bdd_4_lut_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__47301\,
            in1 => \N__47292\,
            in2 => \N__47274\,
            in3 => \N__47263\,
            lcout => n22602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i6_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__46957\,
            in1 => \N__46810\,
            in2 => \N__49487\,
            in3 => \N__46696\,
            lcout => buf_dds1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_245_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__55268\,
            in1 => \N__53775\,
            in2 => \N__46934\,
            in3 => \N__55574\,
            lcout => n12048,
            ltout => \n12048_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001111"
        )
    port map (
            in0 => \N__54843\,
            in1 => \N__54534\,
            in2 => \N__46770\,
            in3 => \N__55269\,
            lcout => n16971,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_clear_301_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__54566\,
            in1 => \N__55387\,
            in2 => \_gnd_net_\,
            in3 => \N__53947\,
            lcout => comm_clear,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56088\,
            ce => \N__50580\,
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12283_12284_reset_LC_18_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48137\,
            lcout => \comm_spi.n14805\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55947\,
            ce => 'H',
            sr => \N__48090\
        );

    \comm_spi.RESET_I_0_90_2_lut_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__58054\,
            in1 => \N__48138\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.iclk_N_802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_91_2_lut_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58053\,
            in2 => \_gnd_net_\,
            in3 => \N__48139\,
            lcout => \comm_spi.iclk_N_803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_213_LC_18_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54874\,
            in2 => \_gnd_net_\,
            in3 => \N__55104\,
            lcout => n21110,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_5__i0_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48078\,
            in1 => \N__54197\,
            in2 => \_gnd_net_\,
            in3 => \N__48708\,
            lcout => comm_buf_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i7_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54196\,
            in1 => \_gnd_net_\,
            in2 => \N__48597\,
            in3 => \N__48066\,
            lcout => comm_buf_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i6_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53226\,
            in1 => \N__48036\,
            in2 => \_gnd_net_\,
            in3 => \N__54200\,
            lcout => comm_buf_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i5_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54195\,
            in1 => \N__53332\,
            in2 => \_gnd_net_\,
            in3 => \N__48021\,
            lcout => comm_buf_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i4_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53645\,
            in1 => \N__48003\,
            in2 => \_gnd_net_\,
            in3 => \N__54199\,
            lcout => comm_buf_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i3_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54194\,
            in1 => \N__49876\,
            in2 => \_gnd_net_\,
            in3 => \N__47973\,
            lcout => comm_buf_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i2_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47949\,
            in1 => \N__50146\,
            in2 => \_gnd_net_\,
            in3 => \N__54198\,
            lcout => comm_buf_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_buf_5__i1_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54193\,
            in1 => \_gnd_net_\,
            in2 => \N__48309\,
            in3 => \N__49721\,
            lcout => comm_buf_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55971\,
            ce => \N__48297\,
            sr => \N__48276\
        );

    \comm_state_1__bdd_4_lut_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__54891\,
            in1 => \N__54173\,
            in2 => \N__52152\,
            in3 => \N__48267\,
            lcout => n22611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__48162\,
            in1 => \N__52690\,
            in2 => \N__54339\,
            in3 => \N__53872\,
            lcout => OPEN,
            ltout => \n2_adj_1576_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22611_bdd_4_lut_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__54892\,
            in1 => \N__53946\,
            in2 => \N__48201\,
            in3 => \N__48198\,
            lcout => n22614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i227_2_lut_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52691\,
            in2 => \_gnd_net_\,
            in3 => \N__52881\,
            lcout => n1348,
            ltout => \n1348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__53873\,
            in1 => \N__48192\,
            in2 => \N__48168\,
            in3 => \N__54177\,
            lcout => n8_adj_1577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__54172\,
            in1 => \N__53870\,
            in2 => \N__48408\,
            in3 => \N__52044\,
            lcout => OPEN,
            ltout => \n21139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_302_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__53871\,
            in1 => \N__55564\,
            in2 => \N__48165\,
            in3 => \N__48161\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i1_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__55120\,
            in1 => \N__48153\,
            in2 => \N__49375\,
            in3 => \N__48147\,
            lcout => comm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55983\,
            ce => \N__52113\,
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_303_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__48417\,
            in1 => \N__48358\,
            in2 => \N__52796\,
            in3 => \N__48462\,
            lcout => n21013,
            ltout => \n21013_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__48359\,
            in1 => \N__52038\,
            in2 => \N__48456\,
            in3 => \N__48315\,
            lcout => n21035,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_312_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001111111011"
        )
    port map (
            in0 => \N__52863\,
            in1 => \N__54179\,
            in2 => \N__52795\,
            in3 => \N__53923\,
            lcout => n4_adj_1589,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_297_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__52513\,
            in1 => \N__52938\,
            in2 => \N__48444\,
            in3 => \N__52055\,
            lcout => n4_adj_1623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15288_2_lut_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54178\,
            in2 => \_gnd_net_\,
            in3 => \N__53922\,
            lcout => n3,
            ltout => \n3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_4_lut_adj_305_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__52781\,
            in1 => \N__48407\,
            in2 => \N__48363\,
            in3 => \N__52862\,
            lcout => OPEN,
            ltout => \n20095_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_46_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__48360\,
            in1 => \N__48330\,
            in2 => \N__48324\,
            in3 => \N__48321\,
            lcout => n21033,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_314_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__52150\,
            in1 => \N__48792\,
            in2 => \_gnd_net_\,
            in3 => \N__52861\,
            lcout => n11619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__55537\,
            in1 => \N__55028\,
            in2 => \N__53986\,
            in3 => \N__54840\,
            lcout => n11600,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i3_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011101"
        )
    port map (
            in0 => \N__55029\,
            in1 => \N__49401\,
            in2 => \N__49386\,
            in3 => \N__48891\,
            lcout => comm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56010\,
            ce => \N__48879\,
            sr => \_gnd_net_\
        );

    \i18492_3_lut_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__48870\,
            in1 => \N__48858\,
            in2 => \_gnd_net_\,
            in3 => \N__48831\,
            lcout => OPEN,
            ltout => \n21219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_308_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__48807\,
            in1 => \N__48791\,
            in2 => \N__48768\,
            in3 => \N__48741\,
            lcout => n21089,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_49_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__55536\,
            in1 => \N__54839\,
            in2 => \_gnd_net_\,
            in3 => \N__55027\,
            lcout => n21043,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i0_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__48720\,
            in1 => \N__54433\,
            in2 => \_gnd_net_\,
            in3 => \N__48707\,
            lcout => comm_buf_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i7_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54432\,
            in1 => \N__48615\,
            in2 => \_gnd_net_\,
            in3 => \N__48600\,
            lcout => comm_buf_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i6_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53225\,
            in1 => \N__48492\,
            in2 => \_gnd_net_\,
            in3 => \N__54436\,
            lcout => comm_buf_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i5_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__54431\,
            in1 => \_gnd_net_\,
            in2 => \N__53344\,
            in3 => \N__48477\,
            lcout => comm_buf_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53636\,
            in1 => \N__49905\,
            in2 => \_gnd_net_\,
            in3 => \N__54435\,
            lcout => comm_buf_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i3_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54430\,
            in1 => \N__49875\,
            in2 => \_gnd_net_\,
            in3 => \N__49788\,
            lcout => comm_buf_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i2_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50156\,
            in1 => \N__49767\,
            in2 => \_gnd_net_\,
            in3 => \N__54434\,
            lcout => comm_buf_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \comm_buf_3__i1_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54429\,
            in1 => \N__49704\,
            in2 => \_gnd_net_\,
            in3 => \N__49632\,
            lcout => comm_buf_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => \N__49428\,
            sr => \N__49413\
        );

    \mux_137_Mux_6_i4_3_lut_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53031\,
            in1 => \N__49623\,
            in2 => \_gnd_net_\,
            in3 => \N__49614\,
            lcout => n4_adj_1581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19789_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__49602\,
            in1 => \N__52394\,
            in2 => \N__49596\,
            in3 => \N__53032\,
            lcout => OPEN,
            ltout => \n22545_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22545_bdd_4_lut_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52395\,
            in1 => \N__49557\,
            in2 => \N__49500\,
            in3 => \N__49486\,
            lcout => n22548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12463_2_lut_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55164\,
            in2 => \_gnd_net_\,
            in3 => \N__49424\,
            lcout => n14979,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i2_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__55165\,
            in1 => \N__50073\,
            in2 => \N__50169\,
            in3 => \N__53126\,
            lcout => comm_buf_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56041\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_0_i4_3_lut_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50061\,
            in1 => \N__50049\,
            in2 => \_gnd_net_\,
            in3 => \N__53030\,
            lcout => n4_adj_1457,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_1_i4_3_lut_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53033\,
            in1 => \N__50031\,
            in2 => \_gnd_net_\,
            in3 => \N__50019\,
            lcout => n4_adj_1588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12491_3_lut_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__50321\,
            in1 => \N__55163\,
            in2 => \_gnd_net_\,
            in3 => \N__50007\,
            lcout => n15007,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19086_2_lut_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49977\,
            in2 => \_gnd_net_\,
            in3 => \N__53067\,
            lcout => OPEN,
            ltout => \n21433_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19741_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__52436\,
            in1 => \N__49959\,
            in2 => \N__49953\,
            in3 => \N__52562\,
            lcout => OPEN,
            ltout => \n22419_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i1_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52563\,
            in1 => \N__53358\,
            in2 => \N__49950\,
            in3 => \N__53517\,
            lcout => comm_tx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56057\,
            ce => \N__50354\,
            sr => \N__50227\
        );

    \i2_2_lut_3_lut_adj_284_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__52435\,
            in1 => \N__52561\,
            in2 => \_gnd_net_\,
            in3 => \N__49947\,
            lcout => OPEN,
            ltout => \n7_adj_1458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_232_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__52890\,
            in1 => \N__55573\,
            in2 => \N__49908\,
            in3 => \N__55108\,
            lcout => n12477,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18555_4_lut_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__52438\,
            in1 => \N__50487\,
            in2 => \N__53088\,
            in3 => \N__53068\,
            lcout => OPEN,
            ltout => \n21282_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i6_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52566\,
            in2 => \N__50478\,
            in3 => \N__50475\,
            lcout => comm_tx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56069\,
            ce => \N__50342\,
            sr => \N__50250\
        );

    \i15197_3_lut_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__52564\,
            in1 => \N__50433\,
            in2 => \_gnd_net_\,
            in3 => \N__50423\,
            lcout => OPEN,
            ltout => \n17698_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18543_4_lut_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__50370\,
            in1 => \N__52565\,
            in2 => \N__50361\,
            in3 => \N__52437\,
            lcout => OPEN,
            ltout => \n21270_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i5_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52182\,
            in2 => \N__50358\,
            in3 => \N__53069\,
            lcout => comm_tx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56069\,
            ce => \N__50342\,
            sr => \N__50250\
        );

    \i6_4_lut_adj_274_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50567\,
            in1 => \N__51005\,
            in2 => \N__50535\,
            in3 => \N__50181\,
            lcout => n20996,
            ltout => \n20996_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15361_2_lut_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__51020\,
            in1 => \_gnd_net_\,
            in2 => \N__50184\,
            in3 => \_gnd_net_\,
            lcout => n10_adj_1528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_273_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__50501\,
            in1 => \N__50516\,
            in2 => \N__50553\,
            in3 => \N__51044\,
            lcout => n12_adj_1663,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclk_294_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__50729\,
            in1 => \_gnd_net_\,
            in2 => \N__51024\,
            in3 => \N__50175\,
            lcout => dds0_mclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclk_294C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_16MHz_I_0_3_lut_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__50811\,
            in1 => \N__50730\,
            in2 => \_gnd_net_\,
            in3 => \N__50721\,
            lcout => \DDS_MCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_65_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__50670\,
            in1 => \N__50644\,
            in2 => \N__50628\,
            in3 => \N__50605\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_272_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__54342\,
            in1 => \N__55272\,
            in2 => \_gnd_net_\,
            in3 => \N__53987\,
            lcout => n11590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i0_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50568\,
            in2 => \_gnd_net_\,
            in3 => \N__50556\,
            lcout => dds0_mclkcnt_0,
            ltout => OPEN,
            carryin => \bfn_18_16_0_\,
            carryout => n19925,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i1_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50552\,
            in2 => \_gnd_net_\,
            in3 => \N__50538\,
            lcout => dds0_mclkcnt_1,
            ltout => OPEN,
            carryin => n19925,
            carryout => n19926,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i2_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50534\,
            in2 => \_gnd_net_\,
            in3 => \N__50520\,
            lcout => dds0_mclkcnt_2,
            ltout => OPEN,
            carryin => n19926,
            carryout => n19927,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i3_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50517\,
            in2 => \_gnd_net_\,
            in3 => \N__50505\,
            lcout => dds0_mclkcnt_3,
            ltout => OPEN,
            carryin => n19927,
            carryout => n19928,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i4_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50502\,
            in2 => \_gnd_net_\,
            in3 => \N__50490\,
            lcout => dds0_mclkcnt_4,
            ltout => OPEN,
            carryin => n19928,
            carryout => n19929,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i5_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51045\,
            in2 => \_gnd_net_\,
            in3 => \N__51033\,
            lcout => dds0_mclkcnt_5,
            ltout => OPEN,
            carryin => n19929,
            carryout => n19930,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i6_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51030\,
            in2 => \_gnd_net_\,
            in3 => \N__51012\,
            lcout => dds0_mclkcnt_6,
            ltout => OPEN,
            carryin => n19930,
            carryout => n19931,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i7_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51006\,
            in2 => \_gnd_net_\,
            in3 => \N__51009\,
            lcout => dds0_mclkcnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12205_2_lut_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54516\,
            in2 => \_gnd_net_\,
            in3 => \N__55233\,
            lcout => n14716,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_12313_12314_set_LC_19_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__57417\,
            in1 => \N__57441\,
            in2 => \_gnd_net_\,
            in3 => \N__57399\,
            lcout => \comm_spi.n14834\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58328\,
            ce => 'H',
            sr => \N__50820\
        );

    \comm_spi.RESET_I_0_89_2_lut_LC_19_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50875\,
            in2 => \_gnd_net_\,
            in3 => \N__58051\,
            lcout => \comm_spi.imosi_N_793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_96_2_lut_LC_19_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__58052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56154\,
            lcout => \comm_spi.data_tx_7__N_810\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i1_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__56230\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56574\,
            lcout => \ADC_VDC.genclk.div_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i1C_net\,
            ce => \N__53691\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19403_2_lut_LC_19_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__56229\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56573\,
            lcout => \ADC_VDC.genclk.n11900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_26_LC_19_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__52005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51903\,
            lcout => OPEN,
            ltout => \ADC_VDC.n52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16282_4_lut_LC_19_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100011011100"
        )
    port map (
            in0 => \N__51760\,
            in1 => \N__51479\,
            in2 => \N__51216\,
            in3 => \N__51204\,
            lcout => \ADC_VDC.n11905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0off_i0_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56340\,
            in2 => \_gnd_net_\,
            in3 => \N__51063\,
            lcout => \ADC_VDC.genclk.t0off_0\,
            ltout => OPEN,
            carryin => \bfn_19_7_0_\,
            carryout => \ADC_VDC.genclk.n19888\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i1_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56370\,
            in2 => \N__58743\,
            in3 => \N__51060\,
            lcout => \ADC_VDC.genclk.t0off_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19888\,
            carryout => \ADC_VDC.genclk.n19889\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i2_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58656\,
            in2 => \N__53742\,
            in3 => \N__51057\,
            lcout => \ADC_VDC.genclk.t0off_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19889\,
            carryout => \ADC_VDC.genclk.n19890\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56279\,
            in2 => \N__58744\,
            in3 => \N__51054\,
            lcout => \ADC_VDC.genclk.t0off_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19890\,
            carryout => \ADC_VDC.genclk.n19891\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i4_LC_19_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58660\,
            in2 => \N__56358\,
            in3 => \N__51051\,
            lcout => \ADC_VDC.genclk.t0off_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19891\,
            carryout => \ADC_VDC.genclk.n19892\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i5_LC_19_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56264\,
            in2 => \N__58745\,
            in3 => \N__51048\,
            lcout => \ADC_VDC.genclk.t0off_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19892\,
            carryout => \ADC_VDC.genclk.n19893\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i6_LC_19_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58664\,
            in2 => \N__56385\,
            in3 => \N__52032\,
            lcout => \ADC_VDC.genclk.t0off_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19893\,
            carryout => \ADC_VDC.genclk.n19894\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i7_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53726\,
            in2 => \N__58746\,
            in3 => \N__52029\,
            lcout => \ADC_VDC.genclk.t0off_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19894\,
            carryout => \ADC_VDC.genclk.n19895\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__52169\,
            sr => \N__58977\
        );

    \ADC_VDC.genclk.t0off_i8_LC_19_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56250\,
            in2 => \N__58718\,
            in3 => \N__52026\,
            lcout => \ADC_VDC.genclk.t0off_8\,
            ltout => OPEN,
            carryin => \bfn_19_8_0_\,
            carryout => \ADC_VDC.genclk.n19896\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i9_LC_19_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58626\,
            in2 => \N__56184\,
            in3 => \N__52023\,
            lcout => \ADC_VDC.genclk.t0off_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19896\,
            carryout => \ADC_VDC.genclk.n19897\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i10_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53711\,
            in2 => \N__58715\,
            in3 => \N__52020\,
            lcout => \ADC_VDC.genclk.t0off_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19897\,
            carryout => \ADC_VDC.genclk.n19898\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i11_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58614\,
            in2 => \N__56541\,
            in3 => \N__52017\,
            lcout => \ADC_VDC.genclk.t0off_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19898\,
            carryout => \ADC_VDC.genclk.n19899\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i12_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53756\,
            in2 => \N__58716\,
            in3 => \N__52014\,
            lcout => \ADC_VDC.genclk.t0off_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19899\,
            carryout => \ADC_VDC.genclk.n19900\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i13_LC_19_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58618\,
            in2 => \N__56298\,
            in3 => \N__52011\,
            lcout => \ADC_VDC.genclk.t0off_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19900\,
            carryout => \ADC_VDC.genclk.n19901\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i14_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56199\,
            in2 => \N__58717\,
            in3 => \N__52008\,
            lcout => \ADC_VDC.genclk.t0off_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19901\,
            carryout => \ADC_VDC.genclk.n19902\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \ADC_VDC.genclk.t0off_i15_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__56168\,
            in1 => \N__58622\,
            in2 => \_gnd_net_\,
            in3 => \N__52173\,
            lcout => \ADC_VDC.genclk.t0off_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__52170\,
            sr => \N__58972\
        );

    \i19104_2_lut_3_lut_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__52763\,
            in1 => \N__54183\,
            in2 => \_gnd_net_\,
            in3 => \N__52857\,
            lcout => n21453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_306_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52767\,
            in2 => \_gnd_net_\,
            in3 => \N__53919\,
            lcout => n14350,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19264_4_lut_4_lut_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000010000"
        )
    port map (
            in0 => \N__54875\,
            in1 => \N__54184\,
            in2 => \N__52793\,
            in3 => \N__52858\,
            lcout => OPEN,
            ltout => \n21454_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19433_4_lut_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__52122\,
            in1 => \N__55065\,
            in2 => \N__52116\,
            in3 => \N__53921\,
            lcout => n14_adj_1638,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i2_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52107\,
            in1 => \N__52056\,
            in2 => \_gnd_net_\,
            in3 => \N__52094\,
            lcout => comm_length_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3881_2_lut_3_lut_LC_19_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__52860\,
            in1 => \N__52769\,
            in2 => \_gnd_net_\,
            in3 => \N__52986\,
            lcout => n6401,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4211_2_lut_LC_19_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__52770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52856\,
            lcout => n6541,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_4_lut_LC_19_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111101111"
        )
    port map (
            in0 => \N__52859\,
            in1 => \N__52768\,
            in2 => \N__54340\,
            in3 => \N__53920\,
            lcout => n21154,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i1_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__52987\,
            in1 => \N__52376\,
            in2 => \N__52794\,
            in3 => \N__52880\,
            lcout => comm_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56027\,
            ce => \N__54903\,
            sr => \N__52647\
        );

    \comm_index_i0_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__52879\,
            in1 => \N__52771\,
            in2 => \_gnd_net_\,
            in3 => \N__52988\,
            lcout => comm_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56027\,
            ce => \N__54903\,
            sr => \N__52647\
        );

    \comm_index_i2_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__52653\,
            in1 => \N__52377\,
            in2 => \_gnd_net_\,
            in3 => \N__52512\,
            lcout => comm_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56027\,
            ce => \N__54903\,
            sr => \N__52647\
        );

    \comm_spi.data_tx_i5_12321_12322_set_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__57492\,
            in1 => \N__57537\,
            in2 => \_gnd_net_\,
            in3 => \N__57515\,
            lcout => \comm_spi.n14842\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58392\,
            ce => 'H',
            sr => \N__53655\
        );

    \i19106_2_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52602\,
            in2 => \_gnd_net_\,
            in3 => \N__57267\,
            lcout => n21460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_102_2_lut_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__53674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58126\,
            lcout => \comm_spi.data_tx_7__N_820\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19515_4_lut_3_lut_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__56448\,
            in1 => \_gnd_net_\,
            in2 => \N__58160\,
            in3 => \N__57535\,
            lcout => \comm_spi.n23098\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_2__bdd_4_lut_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__52578\,
            in1 => \N__52392\,
            in2 => \N__52554\,
            in3 => \N__53267\,
            lcout => OPEN,
            ltout => \n22503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22503_bdd_4_lut_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__52393\,
            in1 => \N__52278\,
            in2 => \N__52200\,
            in3 => \N__52197\,
            lcout => n22506,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_94_2_lut_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58127\,
            lcout => \comm_spi.data_tx_7__N_808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i4_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__53552\,
            in1 => \N__53620\,
            in2 => \N__55285\,
            in3 => \N__53130\,
            lcout => comm_buf_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56058\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_1_i2_3_lut_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53538\,
            in1 => \N__53529\,
            in2 => \_gnd_net_\,
            in3 => \N__53042\,
            lcout => n2_adj_1587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_1_i1_3_lut_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53503\,
            in1 => \N__53424\,
            in2 => \_gnd_net_\,
            in3 => \N__53029\,
            lcout => n1_adj_1586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i5_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__53268\,
            in1 => \N__55180\,
            in2 => \N__53349\,
            in3 => \N__53127\,
            lcout => comm_buf_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19164_2_lut_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53256\,
            in2 => \_gnd_net_\,
            in3 => \N__57266\,
            lcout => n21547,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i6_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__53087\,
            in1 => \N__55281\,
            in2 => \N__53234\,
            in3 => \N__53131\,
            lcout => comm_buf_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53028\,
            in2 => \N__54894\,
            in3 => \N__54417\,
            lcout => n8_adj_1456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_104_2_lut_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__56147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58113\,
            lcout => \comm_spi.data_tx_7__N_826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_response_302_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001101010000"
        )
    port map (
            in0 => \N__54004\,
            in1 => \N__54887\,
            in2 => \N__54515\,
            in3 => \N__55280\,
            lcout => \ICE_GPMI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56089\,
            ce => \N__55599\,
            sr => \_gnd_net_\
        );

    \i17_3_lut_3_lut_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__54886\,
            in1 => \N__54410\,
            in2 => \_gnd_net_\,
            in3 => \N__54003\,
            lcout => OPEN,
            ltout => \n10_adj_1619_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_288_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55578\,
            in2 => \N__55482\,
            in3 => \N__55279\,
            lcout => n12079,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_227_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__54885\,
            in1 => \N__54409\,
            in2 => \_gnd_net_\,
            in3 => \N__54002\,
            lcout => n10804,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_LC_20_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__53760\,
            in1 => \N__53741\,
            in2 => \N__53727\,
            in3 => \N__53712\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19142_4_lut_LC_20_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56526\,
            in1 => \N__56238\,
            in2 => \N__53697\,
            in3 => \N__56328\,
            lcout => \ADC_VDC.genclk.n21598\,
            ltout => \ADC_VDC.genclk.n21598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19468_2_lut_4_lut_LC_20_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101111111111"
        )
    port map (
            in0 => \N__56578\,
            in1 => \N__56319\,
            in2 => \N__53694\,
            in3 => \N__56231\,
            lcout => \ADC_VDC.genclk.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19033_4_lut_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__56381\,
            in1 => \N__56369\,
            in2 => \N__56357\,
            in3 => \N__56339\,
            lcout => \ADC_VDC.genclk.n21600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_adj_25_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57677\,
            in1 => \N__57816\,
            in2 => \N__57567\,
            in3 => \N__57858\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n27_adj_1449_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19193_4_lut_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56205\,
            in1 => \N__56517\,
            in2 => \N__56322\,
            in3 => \N__56304\,
            lcout => \ADC_VDC.genclk.n21597\,
            ltout => \ADC_VDC.genclk.n21597_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i0_LC_20_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__56572\,
            in1 => \N__56313\,
            in2 => \N__56307\,
            in3 => \N__56232\,
            lcout => \ADC_VDC.genclk.div_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19022_4_lut_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__57587\,
            in1 => \N__57714\,
            in2 => \N__57636\,
            in3 => \N__57696\,
            lcout => \ADC_VDC.genclk.n21603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56297\,
            in1 => \N__56280\,
            in2 => \N__56265\,
            in3 => \N__56249\,
            lcout => \ADC_VDC.genclk.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19414_2_lut_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56228\,
            in2 => \_gnd_net_\,
            in3 => \N__56571\,
            lcout => \ADC_VDC.genclk.n14894\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_adj_23_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57774\,
            in1 => \N__57878\,
            in2 => \N__57753\,
            in3 => \N__57836\,
            lcout => \ADC_VDC.genclk.n28_adj_1447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56198\,
            in1 => \N__56180\,
            in2 => \N__56169\,
            in3 => \N__56537\,
            lcout => \ADC_VDC.genclk.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_adj_24_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57794\,
            in1 => \N__57897\,
            in2 => \N__57612\,
            in3 => \N__57657\,
            lcout => \ADC_VDC.genclk.n26_adj_1448\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i4_12317_12318_reset_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56511\,
            in1 => \N__56486\,
            in2 => \_gnd_net_\,
            in3 => \N__57371\,
            lcout => \comm_spi.n14839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58384\,
            ce => 'H',
            sr => \N__56466\
        );

    \comm_spi.data_tx_i2_12309_12310_set_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58800\,
            in1 => \N__58860\,
            in2 => \_gnd_net_\,
            in3 => \N__58910\,
            lcout => \comm_spi.n14830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58406\,
            ce => 'H',
            sr => \N__56457\
        );

    \comm_spi.RESET_I_0_103_2_lut_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56446\,
            in2 => \_gnd_net_\,
            in3 => \N__58131\,
            lcout => \comm_spi.data_tx_7__N_823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_97_2_lut_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__56402\,
            in1 => \_gnd_net_\,
            in2 => \N__58162\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_811\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_105_2_lut_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56401\,
            in2 => \_gnd_net_\,
            in3 => \N__58132\,
            lcout => \comm_spi.data_tx_7__N_829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_95_2_lut_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__56447\,
            in1 => \_gnd_net_\,
            in2 => \N__58161\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_809\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19505_4_lut_3_lut_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__57430\,
            in1 => \N__56403\,
            in2 => \_gnd_net_\,
            in3 => \N__58139\,
            lcout => \comm_spi.n23104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i2_12309_12310_reset_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58796\,
            in1 => \N__58856\,
            in2 => \_gnd_net_\,
            in3 => \N__58914\,
            lcout => \comm_spi.n14831\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58367\,
            ce => 'H',
            sr => \N__57546\
        );

    \comm_spi.data_tx_i5_12321_12322_reset_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57536\,
            in1 => \N__57519\,
            in2 => \_gnd_net_\,
            in3 => \N__57491\,
            lcout => \comm_spi.n14843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58407\,
            ce => 'H',
            sr => \N__57450\
        );

    \comm_spi.data_tx_i3_12313_12314_reset_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57437\,
            in1 => \N__57413\,
            in2 => \_gnd_net_\,
            in3 => \N__57395\,
            lcout => \comm_spi.n14835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58412\,
            ce => 'H',
            sr => \N__57354\
        );

    \i19378_2_lut_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57342\,
            in2 => \_gnd_net_\,
            in3 => \N__57127\,
            lcout => n21456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19099_2_lut_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57324\,
            in2 => \_gnd_net_\,
            in3 => \N__57264\,
            lcout => n21447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19145_2_lut_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__57300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57265\,
            lcout => n21512,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19302_2_lut_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57279\,
            in2 => \_gnd_net_\,
            in3 => \N__57263\,
            lcout => n21434,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12279_12280_reset_LC_22_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58721\,
            lcout => \comm_spi.n14801\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58371\,
            ce => 'H',
            sr => \N__58926\
        );

    \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_22_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56582\,
            lcout => \ADC_VDC.genclk.div_state_1__N_1432\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0on_i0_LC_22_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57713\,
            in2 => \_gnd_net_\,
            in3 => \N__57699\,
            lcout => \ADC_VDC.genclk.t0on_0\,
            ltout => OPEN,
            carryin => \bfn_22_7_0_\,
            carryout => \ADC_VDC.genclk.n19903\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i1_LC_22_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57695\,
            in2 => \N__58751\,
            in3 => \N__57681\,
            lcout => \ADC_VDC.genclk.t0on_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19903\,
            carryout => \ADC_VDC.genclk.n19904\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i2_LC_22_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58687\,
            in2 => \N__57678\,
            in3 => \N__57660\,
            lcout => \ADC_VDC.genclk.t0on_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19904\,
            carryout => \ADC_VDC.genclk.n19905\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i3_LC_22_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57653\,
            in2 => \N__58752\,
            in3 => \N__57639\,
            lcout => \ADC_VDC.genclk.t0on_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19905\,
            carryout => \ADC_VDC.genclk.n19906\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i4_LC_22_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58691\,
            in2 => \N__57635\,
            in3 => \N__57615\,
            lcout => \ADC_VDC.genclk.t0on_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19906\,
            carryout => \ADC_VDC.genclk.n19907\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i5_LC_22_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57605\,
            in2 => \N__58753\,
            in3 => \N__57591\,
            lcout => \ADC_VDC.genclk.t0on_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19907\,
            carryout => \ADC_VDC.genclk.n19908\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i6_LC_22_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58695\,
            in2 => \N__57588\,
            in3 => \N__57570\,
            lcout => \ADC_VDC.genclk.t0on_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19908\,
            carryout => \ADC_VDC.genclk.n19909\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i7_LC_22_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57563\,
            in2 => \N__58754\,
            in3 => \N__57549\,
            lcout => \ADC_VDC.genclk.t0on_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19909\,
            carryout => \ADC_VDC.genclk.n19910\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__57735\,
            sr => \N__58973\
        );

    \ADC_VDC.genclk.t0on_i8_LC_22_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57896\,
            in2 => \N__58750\,
            in3 => \N__57882\,
            lcout => \ADC_VDC.genclk.t0on_8\,
            ltout => OPEN,
            carryin => \bfn_22_8_0_\,
            carryout => \ADC_VDC.genclk.n19911\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i9_LC_22_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58683\,
            in2 => \N__57879\,
            in3 => \N__57861\,
            lcout => \ADC_VDC.genclk.t0on_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19911\,
            carryout => \ADC_VDC.genclk.n19912\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i10_LC_22_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57854\,
            in2 => \N__58747\,
            in3 => \N__57840\,
            lcout => \ADC_VDC.genclk.t0on_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19912\,
            carryout => \ADC_VDC.genclk.n19913\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i11_LC_22_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58671\,
            in2 => \N__57837\,
            in3 => \N__57819\,
            lcout => \ADC_VDC.genclk.t0on_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19913\,
            carryout => \ADC_VDC.genclk.n19914\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i12_LC_22_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57812\,
            in2 => \N__58748\,
            in3 => \N__57798\,
            lcout => \ADC_VDC.genclk.t0on_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19914\,
            carryout => \ADC_VDC.genclk.n19915\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i13_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58675\,
            in2 => \N__57795\,
            in3 => \N__57777\,
            lcout => \ADC_VDC.genclk.t0on_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19915\,
            carryout => \ADC_VDC.genclk.n19916\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i14_LC_22_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57773\,
            in2 => \N__58749\,
            in3 => \N__57759\,
            lcout => \ADC_VDC.genclk.t0on_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19916\,
            carryout => \ADC_VDC.genclk.n19917\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \ADC_VDC.genclk.t0on_i15_LC_22_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__57749\,
            in1 => \N__58679\,
            in2 => \_gnd_net_\,
            in3 => \N__57756\,
            lcout => \ADC_VDC.genclk.t0on_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__57734\,
            sr => \N__58968\
        );

    \comm_spi.RESET_I_0_2_lut_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__58163\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58193\,
            lcout => \comm_spi.data_tx_7__N_835\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19530_4_lut_3_lut_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__58194\,
            in1 => \N__58891\,
            in2 => \_gnd_net_\,
            in3 => \N__58164\,
            lcout => \comm_spi.n23110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i1_12305_12306_reset_LC_22_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58892\,
            in1 => \N__58431\,
            in2 => \_gnd_net_\,
            in3 => \N__58874\,
            lcout => \comm_spi.n14827\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58408\,
            ce => 'H',
            sr => \N__58830\
        );

    \comm_spi.data_tx_i1_12305_12306_set_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__58896\,
            in1 => \N__58430\,
            in2 => \_gnd_net_\,
            in3 => \N__58875\,
            lcout => \comm_spi.n14826\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58399\,
            ce => 'H',
            sr => \N__58839\
        );

    \comm_spi.RESET_I_0_98_2_lut_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__58817\,
            in1 => \_gnd_net_\,
            in2 => \N__58166\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_812\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_106_2_lut_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58816\,
            in2 => \_gnd_net_\,
            in3 => \N__58149\,
            lcout => \comm_spi.data_tx_7__N_832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19495_4_lut_3_lut_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__58818\,
            in1 => \_gnd_net_\,
            in2 => \N__58167\,
            in3 => \N__58789\,
            lcout => \comm_spi.n23107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12279_12280_set_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58765\,
            lcout => \comm_spi.n14800\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__58413\,
            ce => 'H',
            sr => \N__57903\
        );

    \comm_spi.RESET_I_0_99_2_lut_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__58192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58157\,
            lcout => \comm_spi.data_tx_7__N_813\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
