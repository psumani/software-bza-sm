zim_pll_inst: zim_pll
port map(
          REFERENCECLK => ,
          PLLOUTCOREA => ,
          PLLOUTCOREB => ,
          PLLOUTGLOBALA => ,
          PLLOUTGLOBALB => ,
          RESET => 
        );
