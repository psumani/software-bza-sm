// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 28 2024 17:12:41

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "zim" view "INTERFACE"

module zim (
    VAC_DRDY,
    IAC_FLT1,
    DDS_SCK,
    ICE_IOR_166,
    ICE_IOR_119,
    DDS_MOSI,
    VAC_MISO,
    DDS_MOSI1,
    ICE_IOR_146,
    VDC_CLK,
    ICE_IOT_222,
    IAC_CS,
    ICE_IOL_18B,
    ICE_IOL_13A,
    ICE_IOB_81,
    VAC_OSR1,
    IAC_MOSI,
    DDS_CS1,
    ICE_IOL_4B,
    ICE_IOB_94,
    VAC_CS,
    VAC_CLK,
    ICE_SPI_CE0,
    ICE_IOR_167,
    ICE_IOR_118,
    RTD_SDO,
    IAC_OSR0,
    VDC_SCLK,
    VAC_FLT1,
    ICE_SPI_MOSI,
    ICE_IOR_165,
    ICE_IOR_147,
    ICE_IOL_14A,
    ICE_IOL_13B,
    ICE_IOB_91,
    ICE_GPMO_0,
    DDS_RNG_0,
    VDC_RNG0,
    ICE_SPI_SCLK,
    ICE_IOR_152,
    ICE_IOL_12A,
    RTD_DRDY,
    ICE_SPI_MISO,
    ICE_IOT_177,
    ICE_IOR_141,
    ICE_IOB_102,
    ICE_GPMO_2,
    ICE_GPMI_0,
    IAC_MISO,
    VAC_OSR0,
    VAC_MOSI,
    TEST_LED,
    ICE_IOR_148,
    STAT_COMM,
    ICE_SYSCLK,
    ICE_IOR_161,
    ICE_IOB_95,
    ICE_IOB_82,
    ICE_IOB_104,
    IAC_CLK,
    DDS_CS,
    SELIRNG0,
    RTD_SDI,
    ICE_IOT_221,
    ICE_IOT_197,
    DDS_MCLK,
    RTD_SCLK,
    RTD_CS,
    ICE_IOR_137,
    IAC_OSR1,
    VAC_FLT0,
    ICE_IOR_144,
    ICE_IOR_128,
    ICE_GPMO_1,
    IAC_SCLK,
    EIS_SYNCCLK,
    ICE_IOR_139,
    ICE_IOL_4A,
    VAC_SCLK,
    THERMOSTAT,
    ICE_IOR_164,
    ICE_IOB_103,
    OUT_SYNCCLK,
    AMPV_POW,
    VDC_SDO,
    ICE_IOT_174,
    ICE_IOR_140,
    ICE_IOB_96,
    CONT_SD,
    AC_ADC_SYNC,
    SELIRNG1,
    ICE_IOL_12B,
    ICE_IOR_160,
    ICE_IOR_136,
    DDS_MCLK1,
    ICE_IOT_198,
    ICE_IOT_173,
    IAC_DRDY,
    ICE_IOT_178,
    ICE_IOR_138,
    ICE_IOR_120,
    IAC_FLT0,
    DDS_SCK1);

    input VAC_DRDY;
    output IAC_FLT1;
    output DDS_SCK;
    input ICE_IOR_166;
    input ICE_IOR_119;
    output DDS_MOSI;
    input VAC_MISO;
    output DDS_MOSI1;
    input ICE_IOR_146;
    output VDC_CLK;
    input ICE_IOT_222;
    output IAC_CS;
    input ICE_IOL_18B;
    input ICE_IOL_13A;
    input ICE_IOB_81;
    output VAC_OSR1;
    output IAC_MOSI;
    output DDS_CS1;
    input ICE_IOL_4B;
    input ICE_IOB_94;
    output VAC_CS;
    output VAC_CLK;
    input ICE_SPI_CE0;
    input ICE_IOR_167;
    input ICE_IOR_118;
    input RTD_SDO;
    output IAC_OSR0;
    output VDC_SCLK;
    output VAC_FLT1;
    input ICE_SPI_MOSI;
    input ICE_IOR_165;
    input ICE_IOR_147;
    input ICE_IOL_14A;
    input ICE_IOL_13B;
    input ICE_IOB_91;
    input ICE_GPMO_0;
    output DDS_RNG_0;
    output VDC_RNG0;
    input ICE_SPI_SCLK;
    input ICE_IOR_152;
    input ICE_IOL_12A;
    input RTD_DRDY;
    output ICE_SPI_MISO;
    input ICE_IOT_177;
    input ICE_IOR_141;
    input ICE_IOB_102;
    input ICE_GPMO_2;
    output ICE_GPMI_0;
    input IAC_MISO;
    output VAC_OSR0;
    output VAC_MOSI;
    output TEST_LED;
    input ICE_IOR_148;
    output STAT_COMM;
    input ICE_SYSCLK;
    input ICE_IOR_161;
    input ICE_IOB_95;
    input ICE_IOB_82;
    input ICE_IOB_104;
    output IAC_CLK;
    output DDS_CS;
    output SELIRNG0;
    output RTD_SDI;
    input ICE_IOT_221;
    input ICE_IOT_197;
    output DDS_MCLK;
    output RTD_SCLK;
    output RTD_CS;
    input ICE_IOR_137;
    output IAC_OSR1;
    output VAC_FLT0;
    input ICE_IOR_144;
    input ICE_IOR_128;
    input ICE_GPMO_1;
    output IAC_SCLK;
    input EIS_SYNCCLK;
    input ICE_IOR_139;
    input ICE_IOL_4A;
    output VAC_SCLK;
    input THERMOSTAT;
    input ICE_IOR_164;
    input ICE_IOB_103;
    output OUT_SYNCCLK;
    output AMPV_POW;
    input VDC_SDO;
    input ICE_IOT_174;
    input ICE_IOR_140;
    input ICE_IOB_96;
    output CONT_SD;
    output AC_ADC_SYNC;
    output SELIRNG1;
    input ICE_IOL_12B;
    input ICE_IOR_160;
    input ICE_IOR_136;
    output DDS_MCLK1;
    input ICE_IOT_198;
    input ICE_IOT_173;
    input IAC_DRDY;
    input ICE_IOT_178;
    input ICE_IOR_138;
    input ICE_IOR_120;
    output IAC_FLT0;
    output DDS_SCK1;

    wire N__59184;
    wire N__59183;
    wire N__59182;
    wire N__59175;
    wire N__59174;
    wire N__59173;
    wire N__59166;
    wire N__59165;
    wire N__59164;
    wire N__59157;
    wire N__59156;
    wire N__59155;
    wire N__59148;
    wire N__59147;
    wire N__59146;
    wire N__59139;
    wire N__59138;
    wire N__59137;
    wire N__59130;
    wire N__59129;
    wire N__59128;
    wire N__59121;
    wire N__59120;
    wire N__59119;
    wire N__59112;
    wire N__59111;
    wire N__59110;
    wire N__59103;
    wire N__59102;
    wire N__59101;
    wire N__59094;
    wire N__59093;
    wire N__59092;
    wire N__59085;
    wire N__59084;
    wire N__59083;
    wire N__59076;
    wire N__59075;
    wire N__59074;
    wire N__59067;
    wire N__59066;
    wire N__59065;
    wire N__59058;
    wire N__59057;
    wire N__59056;
    wire N__59049;
    wire N__59048;
    wire N__59047;
    wire N__59040;
    wire N__59039;
    wire N__59038;
    wire N__59031;
    wire N__59030;
    wire N__59029;
    wire N__59022;
    wire N__59021;
    wire N__59020;
    wire N__59013;
    wire N__59012;
    wire N__59011;
    wire N__59004;
    wire N__59003;
    wire N__59002;
    wire N__58995;
    wire N__58994;
    wire N__58993;
    wire N__58986;
    wire N__58985;
    wire N__58984;
    wire N__58977;
    wire N__58976;
    wire N__58975;
    wire N__58968;
    wire N__58967;
    wire N__58966;
    wire N__58959;
    wire N__58958;
    wire N__58957;
    wire N__58950;
    wire N__58949;
    wire N__58948;
    wire N__58941;
    wire N__58940;
    wire N__58939;
    wire N__58932;
    wire N__58931;
    wire N__58930;
    wire N__58923;
    wire N__58922;
    wire N__58921;
    wire N__58914;
    wire N__58913;
    wire N__58912;
    wire N__58905;
    wire N__58904;
    wire N__58903;
    wire N__58896;
    wire N__58895;
    wire N__58894;
    wire N__58887;
    wire N__58886;
    wire N__58885;
    wire N__58878;
    wire N__58877;
    wire N__58876;
    wire N__58869;
    wire N__58868;
    wire N__58867;
    wire N__58860;
    wire N__58859;
    wire N__58858;
    wire N__58851;
    wire N__58850;
    wire N__58849;
    wire N__58842;
    wire N__58841;
    wire N__58840;
    wire N__58833;
    wire N__58832;
    wire N__58831;
    wire N__58824;
    wire N__58823;
    wire N__58822;
    wire N__58815;
    wire N__58814;
    wire N__58813;
    wire N__58806;
    wire N__58805;
    wire N__58804;
    wire N__58797;
    wire N__58796;
    wire N__58795;
    wire N__58788;
    wire N__58787;
    wire N__58786;
    wire N__58779;
    wire N__58778;
    wire N__58777;
    wire N__58770;
    wire N__58769;
    wire N__58768;
    wire N__58761;
    wire N__58760;
    wire N__58759;
    wire N__58752;
    wire N__58751;
    wire N__58750;
    wire N__58743;
    wire N__58742;
    wire N__58741;
    wire N__58734;
    wire N__58733;
    wire N__58732;
    wire N__58725;
    wire N__58724;
    wire N__58723;
    wire N__58716;
    wire N__58715;
    wire N__58714;
    wire N__58707;
    wire N__58706;
    wire N__58705;
    wire N__58698;
    wire N__58697;
    wire N__58696;
    wire N__58689;
    wire N__58688;
    wire N__58687;
    wire N__58680;
    wire N__58679;
    wire N__58678;
    wire N__58671;
    wire N__58670;
    wire N__58669;
    wire N__58662;
    wire N__58661;
    wire N__58660;
    wire N__58653;
    wire N__58652;
    wire N__58651;
    wire N__58644;
    wire N__58643;
    wire N__58642;
    wire N__58635;
    wire N__58634;
    wire N__58633;
    wire N__58626;
    wire N__58625;
    wire N__58624;
    wire N__58617;
    wire N__58616;
    wire N__58615;
    wire N__58608;
    wire N__58607;
    wire N__58606;
    wire N__58599;
    wire N__58598;
    wire N__58597;
    wire N__58590;
    wire N__58589;
    wire N__58588;
    wire N__58581;
    wire N__58580;
    wire N__58579;
    wire N__58572;
    wire N__58571;
    wire N__58570;
    wire N__58563;
    wire N__58562;
    wire N__58561;
    wire N__58554;
    wire N__58553;
    wire N__58552;
    wire N__58545;
    wire N__58544;
    wire N__58543;
    wire N__58536;
    wire N__58535;
    wire N__58534;
    wire N__58527;
    wire N__58526;
    wire N__58525;
    wire N__58518;
    wire N__58517;
    wire N__58516;
    wire N__58509;
    wire N__58508;
    wire N__58507;
    wire N__58500;
    wire N__58499;
    wire N__58498;
    wire N__58491;
    wire N__58490;
    wire N__58489;
    wire N__58482;
    wire N__58481;
    wire N__58480;
    wire N__58473;
    wire N__58472;
    wire N__58471;
    wire N__58464;
    wire N__58463;
    wire N__58462;
    wire N__58455;
    wire N__58454;
    wire N__58453;
    wire N__58446;
    wire N__58445;
    wire N__58444;
    wire N__58437;
    wire N__58436;
    wire N__58435;
    wire N__58428;
    wire N__58427;
    wire N__58426;
    wire N__58419;
    wire N__58418;
    wire N__58417;
    wire N__58410;
    wire N__58409;
    wire N__58408;
    wire N__58401;
    wire N__58400;
    wire N__58399;
    wire N__58392;
    wire N__58391;
    wire N__58390;
    wire N__58383;
    wire N__58382;
    wire N__58381;
    wire N__58374;
    wire N__58373;
    wire N__58372;
    wire N__58365;
    wire N__58364;
    wire N__58363;
    wire N__58356;
    wire N__58355;
    wire N__58354;
    wire N__58347;
    wire N__58346;
    wire N__58345;
    wire N__58338;
    wire N__58337;
    wire N__58336;
    wire N__58329;
    wire N__58328;
    wire N__58327;
    wire N__58320;
    wire N__58319;
    wire N__58318;
    wire N__58311;
    wire N__58310;
    wire N__58309;
    wire N__58302;
    wire N__58301;
    wire N__58300;
    wire N__58293;
    wire N__58292;
    wire N__58291;
    wire N__58284;
    wire N__58283;
    wire N__58282;
    wire N__58275;
    wire N__58274;
    wire N__58273;
    wire N__58266;
    wire N__58265;
    wire N__58264;
    wire N__58247;
    wire N__58244;
    wire N__58241;
    wire N__58238;
    wire N__58237;
    wire N__58234;
    wire N__58231;
    wire N__58228;
    wire N__58225;
    wire N__58224;
    wire N__58221;
    wire N__58218;
    wire N__58215;
    wire N__58208;
    wire N__58207;
    wire N__58204;
    wire N__58201;
    wire N__58198;
    wire N__58193;
    wire N__58192;
    wire N__58189;
    wire N__58186;
    wire N__58181;
    wire N__58178;
    wire N__58177;
    wire N__58174;
    wire N__58171;
    wire N__58166;
    wire N__58163;
    wire N__58160;
    wire N__58157;
    wire N__58154;
    wire N__58153;
    wire N__58152;
    wire N__58149;
    wire N__58146;
    wire N__58143;
    wire N__58136;
    wire N__58135;
    wire N__58132;
    wire N__58129;
    wire N__58128;
    wire N__58125;
    wire N__58122;
    wire N__58119;
    wire N__58116;
    wire N__58113;
    wire N__58110;
    wire N__58103;
    wire N__58100;
    wire N__58097;
    wire N__58094;
    wire N__58091;
    wire N__58088;
    wire N__58085;
    wire N__58084;
    wire N__58081;
    wire N__58078;
    wire N__58073;
    wire N__58070;
    wire N__58067;
    wire N__58064;
    wire N__58061;
    wire N__58058;
    wire N__58055;
    wire N__58054;
    wire N__58051;
    wire N__58048;
    wire N__58045;
    wire N__58042;
    wire N__58041;
    wire N__58038;
    wire N__58035;
    wire N__58032;
    wire N__58031;
    wire N__58030;
    wire N__58025;
    wire N__58022;
    wire N__58019;
    wire N__58016;
    wire N__58013;
    wire N__58006;
    wire N__58001;
    wire N__57998;
    wire N__57995;
    wire N__57992;
    wire N__57989;
    wire N__57986;
    wire N__57983;
    wire N__57982;
    wire N__57981;
    wire N__57980;
    wire N__57979;
    wire N__57978;
    wire N__57977;
    wire N__57976;
    wire N__57975;
    wire N__57974;
    wire N__57973;
    wire N__57972;
    wire N__57971;
    wire N__57970;
    wire N__57969;
    wire N__57968;
    wire N__57967;
    wire N__57966;
    wire N__57965;
    wire N__57964;
    wire N__57963;
    wire N__57962;
    wire N__57961;
    wire N__57960;
    wire N__57959;
    wire N__57958;
    wire N__57957;
    wire N__57956;
    wire N__57955;
    wire N__57954;
    wire N__57953;
    wire N__57952;
    wire N__57951;
    wire N__57950;
    wire N__57949;
    wire N__57948;
    wire N__57947;
    wire N__57946;
    wire N__57945;
    wire N__57944;
    wire N__57943;
    wire N__57942;
    wire N__57941;
    wire N__57940;
    wire N__57939;
    wire N__57938;
    wire N__57937;
    wire N__57936;
    wire N__57935;
    wire N__57934;
    wire N__57933;
    wire N__57932;
    wire N__57931;
    wire N__57930;
    wire N__57929;
    wire N__57928;
    wire N__57927;
    wire N__57926;
    wire N__57925;
    wire N__57924;
    wire N__57923;
    wire N__57922;
    wire N__57921;
    wire N__57920;
    wire N__57919;
    wire N__57918;
    wire N__57917;
    wire N__57916;
    wire N__57915;
    wire N__57914;
    wire N__57913;
    wire N__57912;
    wire N__57911;
    wire N__57910;
    wire N__57909;
    wire N__57908;
    wire N__57907;
    wire N__57906;
    wire N__57905;
    wire N__57904;
    wire N__57903;
    wire N__57902;
    wire N__57901;
    wire N__57900;
    wire N__57899;
    wire N__57898;
    wire N__57897;
    wire N__57896;
    wire N__57895;
    wire N__57894;
    wire N__57893;
    wire N__57892;
    wire N__57891;
    wire N__57890;
    wire N__57889;
    wire N__57888;
    wire N__57887;
    wire N__57886;
    wire N__57885;
    wire N__57884;
    wire N__57883;
    wire N__57882;
    wire N__57881;
    wire N__57880;
    wire N__57879;
    wire N__57878;
    wire N__57877;
    wire N__57876;
    wire N__57875;
    wire N__57874;
    wire N__57873;
    wire N__57872;
    wire N__57871;
    wire N__57870;
    wire N__57869;
    wire N__57868;
    wire N__57867;
    wire N__57866;
    wire N__57865;
    wire N__57864;
    wire N__57863;
    wire N__57862;
    wire N__57861;
    wire N__57860;
    wire N__57859;
    wire N__57858;
    wire N__57857;
    wire N__57856;
    wire N__57855;
    wire N__57854;
    wire N__57853;
    wire N__57852;
    wire N__57851;
    wire N__57850;
    wire N__57849;
    wire N__57848;
    wire N__57847;
    wire N__57846;
    wire N__57845;
    wire N__57844;
    wire N__57843;
    wire N__57842;
    wire N__57841;
    wire N__57840;
    wire N__57839;
    wire N__57838;
    wire N__57837;
    wire N__57836;
    wire N__57835;
    wire N__57834;
    wire N__57833;
    wire N__57832;
    wire N__57831;
    wire N__57830;
    wire N__57829;
    wire N__57828;
    wire N__57827;
    wire N__57826;
    wire N__57825;
    wire N__57824;
    wire N__57823;
    wire N__57822;
    wire N__57821;
    wire N__57820;
    wire N__57819;
    wire N__57818;
    wire N__57817;
    wire N__57816;
    wire N__57815;
    wire N__57814;
    wire N__57813;
    wire N__57812;
    wire N__57811;
    wire N__57810;
    wire N__57809;
    wire N__57808;
    wire N__57807;
    wire N__57806;
    wire N__57805;
    wire N__57804;
    wire N__57443;
    wire N__57440;
    wire N__57437;
    wire N__57434;
    wire N__57431;
    wire N__57428;
    wire N__57425;
    wire N__57424;
    wire N__57423;
    wire N__57422;
    wire N__57419;
    wire N__57418;
    wire N__57415;
    wire N__57414;
    wire N__57411;
    wire N__57410;
    wire N__57395;
    wire N__57394;
    wire N__57393;
    wire N__57392;
    wire N__57391;
    wire N__57390;
    wire N__57389;
    wire N__57388;
    wire N__57385;
    wire N__57384;
    wire N__57383;
    wire N__57382;
    wire N__57381;
    wire N__57380;
    wire N__57379;
    wire N__57376;
    wire N__57375;
    wire N__57374;
    wire N__57373;
    wire N__57370;
    wire N__57369;
    wire N__57366;
    wire N__57365;
    wire N__57362;
    wire N__57361;
    wire N__57358;
    wire N__57357;
    wire N__57354;
    wire N__57353;
    wire N__57350;
    wire N__57347;
    wire N__57346;
    wire N__57343;
    wire N__57342;
    wire N__57339;
    wire N__57338;
    wire N__57335;
    wire N__57334;
    wire N__57331;
    wire N__57328;
    wire N__57327;
    wire N__57326;
    wire N__57325;
    wire N__57324;
    wire N__57321;
    wire N__57320;
    wire N__57319;
    wire N__57318;
    wire N__57301;
    wire N__57286;
    wire N__57283;
    wire N__57266;
    wire N__57263;
    wire N__57260;
    wire N__57259;
    wire N__57256;
    wire N__57255;
    wire N__57252;
    wire N__57251;
    wire N__57248;
    wire N__57245;
    wire N__57242;
    wire N__57239;
    wire N__57238;
    wire N__57237;
    wire N__57236;
    wire N__57233;
    wire N__57232;
    wire N__57227;
    wire N__57222;
    wire N__57219;
    wire N__57204;
    wire N__57197;
    wire N__57194;
    wire N__57191;
    wire N__57188;
    wire N__57187;
    wire N__57186;
    wire N__57185;
    wire N__57182;
    wire N__57179;
    wire N__57174;
    wire N__57171;
    wire N__57168;
    wire N__57167;
    wire N__57158;
    wire N__57155;
    wire N__57152;
    wire N__57149;
    wire N__57148;
    wire N__57147;
    wire N__57144;
    wire N__57141;
    wire N__57138;
    wire N__57133;
    wire N__57130;
    wire N__57121;
    wire N__57118;
    wire N__57115;
    wire N__57112;
    wire N__57109;
    wire N__57106;
    wire N__57103;
    wire N__57100;
    wire N__57093;
    wire N__57080;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57070;
    wire N__57067;
    wire N__57062;
    wire N__57059;
    wire N__57058;
    wire N__57055;
    wire N__57052;
    wire N__57051;
    wire N__57050;
    wire N__57049;
    wire N__57044;
    wire N__57041;
    wire N__57040;
    wire N__57037;
    wire N__57036;
    wire N__57035;
    wire N__57032;
    wire N__57027;
    wire N__57024;
    wire N__57021;
    wire N__57018;
    wire N__57017;
    wire N__57016;
    wire N__57013;
    wire N__57012;
    wire N__57009;
    wire N__57004;
    wire N__56999;
    wire N__56998;
    wire N__56997;
    wire N__56996;
    wire N__56995;
    wire N__56992;
    wire N__56991;
    wire N__56988;
    wire N__56987;
    wire N__56984;
    wire N__56983;
    wire N__56980;
    wire N__56975;
    wire N__56972;
    wire N__56969;
    wire N__56966;
    wire N__56963;
    wire N__56960;
    wire N__56957;
    wire N__56954;
    wire N__56951;
    wire N__56948;
    wire N__56945;
    wire N__56942;
    wire N__56939;
    wire N__56936;
    wire N__56931;
    wire N__56926;
    wire N__56919;
    wire N__56918;
    wire N__56917;
    wire N__56912;
    wire N__56911;
    wire N__56910;
    wire N__56907;
    wire N__56904;
    wire N__56899;
    wire N__56892;
    wire N__56889;
    wire N__56886;
    wire N__56883;
    wire N__56880;
    wire N__56877;
    wire N__56858;
    wire N__56855;
    wire N__56854;
    wire N__56853;
    wire N__56852;
    wire N__56849;
    wire N__56846;
    wire N__56845;
    wire N__56844;
    wire N__56843;
    wire N__56842;
    wire N__56841;
    wire N__56838;
    wire N__56837;
    wire N__56836;
    wire N__56835;
    wire N__56834;
    wire N__56833;
    wire N__56832;
    wire N__56829;
    wire N__56824;
    wire N__56823;
    wire N__56818;
    wire N__56817;
    wire N__56816;
    wire N__56811;
    wire N__56810;
    wire N__56809;
    wire N__56808;
    wire N__56807;
    wire N__56804;
    wire N__56795;
    wire N__56792;
    wire N__56787;
    wire N__56784;
    wire N__56781;
    wire N__56778;
    wire N__56777;
    wire N__56776;
    wire N__56775;
    wire N__56772;
    wire N__56767;
    wire N__56764;
    wire N__56761;
    wire N__56760;
    wire N__56755;
    wire N__56752;
    wire N__56751;
    wire N__56750;
    wire N__56749;
    wire N__56748;
    wire N__56747;
    wire N__56746;
    wire N__56745;
    wire N__56744;
    wire N__56743;
    wire N__56742;
    wire N__56737;
    wire N__56732;
    wire N__56727;
    wire N__56724;
    wire N__56719;
    wire N__56716;
    wire N__56713;
    wire N__56706;
    wire N__56703;
    wire N__56698;
    wire N__56695;
    wire N__56684;
    wire N__56675;
    wire N__56672;
    wire N__56667;
    wire N__56662;
    wire N__56655;
    wire N__56650;
    wire N__56633;
    wire N__56632;
    wire N__56629;
    wire N__56628;
    wire N__56625;
    wire N__56622;
    wire N__56619;
    wire N__56616;
    wire N__56611;
    wire N__56608;
    wire N__56605;
    wire N__56600;
    wire N__56597;
    wire N__56594;
    wire N__56591;
    wire N__56588;
    wire N__56585;
    wire N__56584;
    wire N__56581;
    wire N__56578;
    wire N__56577;
    wire N__56572;
    wire N__56569;
    wire N__56564;
    wire N__56563;
    wire N__56560;
    wire N__56557;
    wire N__56554;
    wire N__56549;
    wire N__56546;
    wire N__56543;
    wire N__56542;
    wire N__56539;
    wire N__56536;
    wire N__56535;
    wire N__56530;
    wire N__56527;
    wire N__56524;
    wire N__56521;
    wire N__56516;
    wire N__56513;
    wire N__56510;
    wire N__56507;
    wire N__56506;
    wire N__56505;
    wire N__56502;
    wire N__56499;
    wire N__56496;
    wire N__56489;
    wire N__56488;
    wire N__56487;
    wire N__56484;
    wire N__56481;
    wire N__56478;
    wire N__56475;
    wire N__56470;
    wire N__56467;
    wire N__56464;
    wire N__56459;
    wire N__56456;
    wire N__56455;
    wire N__56452;
    wire N__56449;
    wire N__56444;
    wire N__56441;
    wire N__56438;
    wire N__56435;
    wire N__56432;
    wire N__56429;
    wire N__56426;
    wire N__56425;
    wire N__56422;
    wire N__56419;
    wire N__56414;
    wire N__56411;
    wire N__56408;
    wire N__56405;
    wire N__56402;
    wire N__56399;
    wire N__56396;
    wire N__56395;
    wire N__56394;
    wire N__56391;
    wire N__56388;
    wire N__56385;
    wire N__56378;
    wire N__56377;
    wire N__56374;
    wire N__56373;
    wire N__56372;
    wire N__56371;
    wire N__56370;
    wire N__56369;
    wire N__56368;
    wire N__56367;
    wire N__56364;
    wire N__56363;
    wire N__56362;
    wire N__56361;
    wire N__56360;
    wire N__56359;
    wire N__56358;
    wire N__56357;
    wire N__56348;
    wire N__56345;
    wire N__56342;
    wire N__56341;
    wire N__56340;
    wire N__56339;
    wire N__56338;
    wire N__56337;
    wire N__56336;
    wire N__56335;
    wire N__56334;
    wire N__56333;
    wire N__56332;
    wire N__56331;
    wire N__56330;
    wire N__56329;
    wire N__56326;
    wire N__56325;
    wire N__56324;
    wire N__56323;
    wire N__56322;
    wire N__56321;
    wire N__56320;
    wire N__56319;
    wire N__56318;
    wire N__56317;
    wire N__56314;
    wire N__56313;
    wire N__56310;
    wire N__56309;
    wire N__56306;
    wire N__56305;
    wire N__56304;
    wire N__56303;
    wire N__56302;
    wire N__56301;
    wire N__56300;
    wire N__56299;
    wire N__56298;
    wire N__56297;
    wire N__56296;
    wire N__56295;
    wire N__56292;
    wire N__56291;
    wire N__56288;
    wire N__56287;
    wire N__56286;
    wire N__56283;
    wire N__56282;
    wire N__56281;
    wire N__56278;
    wire N__56275;
    wire N__56272;
    wire N__56271;
    wire N__56270;
    wire N__56269;
    wire N__56268;
    wire N__56265;
    wire N__56264;
    wire N__56263;
    wire N__56260;
    wire N__56257;
    wire N__56254;
    wire N__56253;
    wire N__56252;
    wire N__56251;
    wire N__56250;
    wire N__56249;
    wire N__56248;
    wire N__56247;
    wire N__56246;
    wire N__56245;
    wire N__56244;
    wire N__56241;
    wire N__56238;
    wire N__56237;
    wire N__56236;
    wire N__56231;
    wire N__56226;
    wire N__56223;
    wire N__56216;
    wire N__56213;
    wire N__56210;
    wire N__56207;
    wire N__56204;
    wire N__56197;
    wire N__56188;
    wire N__56187;
    wire N__56186;
    wire N__56185;
    wire N__56184;
    wire N__56183;
    wire N__56182;
    wire N__56181;
    wire N__56180;
    wire N__56177;
    wire N__56174;
    wire N__56171;
    wire N__56168;
    wire N__56167;
    wire N__56166;
    wire N__56163;
    wire N__56160;
    wire N__56159;
    wire N__56154;
    wire N__56145;
    wire N__56144;
    wire N__56143;
    wire N__56140;
    wire N__56137;
    wire N__56132;
    wire N__56129;
    wire N__56126;
    wire N__56123;
    wire N__56120;
    wire N__56115;
    wire N__56112;
    wire N__56107;
    wire N__56106;
    wire N__56103;
    wire N__56100;
    wire N__56097;
    wire N__56094;
    wire N__56087;
    wire N__56084;
    wire N__56079;
    wire N__56074;
    wire N__56073;
    wire N__56072;
    wire N__56071;
    wire N__56068;
    wire N__56061;
    wire N__56056;
    wire N__56051;
    wire N__56046;
    wire N__56043;
    wire N__56040;
    wire N__56037;
    wire N__56032;
    wire N__56029;
    wire N__56020;
    wire N__56009;
    wire N__56008;
    wire N__56007;
    wire N__56006;
    wire N__55999;
    wire N__55996;
    wire N__55993;
    wire N__55988;
    wire N__55985;
    wire N__55978;
    wire N__55975;
    wire N__55970;
    wire N__55967;
    wire N__55964;
    wire N__55961;
    wire N__55956;
    wire N__55953;
    wire N__55950;
    wire N__55949;
    wire N__55948;
    wire N__55947;
    wire N__55946;
    wire N__55945;
    wire N__55944;
    wire N__55943;
    wire N__55940;
    wire N__55935;
    wire N__55932;
    wire N__55929;
    wire N__55924;
    wire N__55917;
    wire N__55914;
    wire N__55909;
    wire N__55900;
    wire N__55897;
    wire N__55894;
    wire N__55891;
    wire N__55886;
    wire N__55881;
    wire N__55876;
    wire N__55873;
    wire N__55864;
    wire N__55857;
    wire N__55850;
    wire N__55847;
    wire N__55842;
    wire N__55839;
    wire N__55836;
    wire N__55831;
    wire N__55818;
    wire N__55817;
    wire N__55816;
    wire N__55813;
    wire N__55810;
    wire N__55803;
    wire N__55798;
    wire N__55795;
    wire N__55788;
    wire N__55781;
    wire N__55770;
    wire N__55755;
    wire N__55740;
    wire N__55735;
    wire N__55712;
    wire N__55709;
    wire N__55706;
    wire N__55703;
    wire N__55700;
    wire N__55697;
    wire N__55694;
    wire N__55691;
    wire N__55688;
    wire N__55685;
    wire N__55684;
    wire N__55681;
    wire N__55678;
    wire N__55673;
    wire N__55670;
    wire N__55667;
    wire N__55664;
    wire N__55661;
    wire N__55658;
    wire N__55655;
    wire N__55654;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55644;
    wire N__55637;
    wire N__55636;
    wire N__55633;
    wire N__55630;
    wire N__55627;
    wire N__55624;
    wire N__55619;
    wire N__55618;
    wire N__55615;
    wire N__55612;
    wire N__55607;
    wire N__55604;
    wire N__55601;
    wire N__55598;
    wire N__55595;
    wire N__55592;
    wire N__55589;
    wire N__55586;
    wire N__55583;
    wire N__55580;
    wire N__55577;
    wire N__55574;
    wire N__55571;
    wire N__55568;
    wire N__55565;
    wire N__55562;
    wire N__55559;
    wire N__55556;
    wire N__55553;
    wire N__55550;
    wire N__55547;
    wire N__55544;
    wire N__55541;
    wire N__55538;
    wire N__55535;
    wire N__55534;
    wire N__55531;
    wire N__55528;
    wire N__55523;
    wire N__55520;
    wire N__55517;
    wire N__55514;
    wire N__55511;
    wire N__55510;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55497;
    wire N__55492;
    wire N__55489;
    wire N__55484;
    wire N__55481;
    wire N__55478;
    wire N__55477;
    wire N__55476;
    wire N__55473;
    wire N__55470;
    wire N__55469;
    wire N__55466;
    wire N__55465;
    wire N__55460;
    wire N__55457;
    wire N__55454;
    wire N__55451;
    wire N__55450;
    wire N__55445;
    wire N__55440;
    wire N__55437;
    wire N__55434;
    wire N__55427;
    wire N__55424;
    wire N__55423;
    wire N__55420;
    wire N__55417;
    wire N__55412;
    wire N__55411;
    wire N__55408;
    wire N__55405;
    wire N__55400;
    wire N__55397;
    wire N__55394;
    wire N__55393;
    wire N__55390;
    wire N__55387;
    wire N__55386;
    wire N__55381;
    wire N__55378;
    wire N__55373;
    wire N__55370;
    wire N__55367;
    wire N__55366;
    wire N__55363;
    wire N__55360;
    wire N__55357;
    wire N__55354;
    wire N__55349;
    wire N__55346;
    wire N__55343;
    wire N__55340;
    wire N__55339;
    wire N__55336;
    wire N__55333;
    wire N__55328;
    wire N__55325;
    wire N__55322;
    wire N__55319;
    wire N__55318;
    wire N__55315;
    wire N__55312;
    wire N__55311;
    wire N__55308;
    wire N__55305;
    wire N__55302;
    wire N__55299;
    wire N__55294;
    wire N__55291;
    wire N__55288;
    wire N__55283;
    wire N__55280;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55272;
    wire N__55267;
    wire N__55264;
    wire N__55259;
    wire N__55256;
    wire N__55253;
    wire N__55250;
    wire N__55247;
    wire N__55246;
    wire N__55241;
    wire N__55238;
    wire N__55237;
    wire N__55234;
    wire N__55231;
    wire N__55226;
    wire N__55223;
    wire N__55220;
    wire N__55219;
    wire N__55218;
    wire N__55215;
    wire N__55212;
    wire N__55209;
    wire N__55202;
    wire N__55201;
    wire N__55198;
    wire N__55195;
    wire N__55190;
    wire N__55187;
    wire N__55186;
    wire N__55183;
    wire N__55180;
    wire N__55175;
    wire N__55172;
    wire N__55169;
    wire N__55166;
    wire N__55163;
    wire N__55160;
    wire N__55157;
    wire N__55154;
    wire N__55153;
    wire N__55152;
    wire N__55149;
    wire N__55144;
    wire N__55141;
    wire N__55138;
    wire N__55135;
    wire N__55132;
    wire N__55127;
    wire N__55124;
    wire N__55123;
    wire N__55120;
    wire N__55117;
    wire N__55112;
    wire N__55109;
    wire N__55106;
    wire N__55103;
    wire N__55100;
    wire N__55097;
    wire N__55094;
    wire N__55091;
    wire N__55088;
    wire N__55085;
    wire N__55082;
    wire N__55079;
    wire N__55076;
    wire N__55073;
    wire N__55070;
    wire N__55069;
    wire N__55068;
    wire N__55065;
    wire N__55062;
    wire N__55059;
    wire N__55052;
    wire N__55049;
    wire N__55046;
    wire N__55043;
    wire N__55040;
    wire N__55039;
    wire N__55036;
    wire N__55033;
    wire N__55028;
    wire N__55027;
    wire N__55024;
    wire N__55021;
    wire N__55020;
    wire N__55017;
    wire N__55014;
    wire N__55011;
    wire N__55008;
    wire N__55003;
    wire N__55000;
    wire N__54997;
    wire N__54992;
    wire N__54989;
    wire N__54986;
    wire N__54983;
    wire N__54982;
    wire N__54981;
    wire N__54978;
    wire N__54977;
    wire N__54976;
    wire N__54975;
    wire N__54974;
    wire N__54973;
    wire N__54972;
    wire N__54971;
    wire N__54968;
    wire N__54967;
    wire N__54966;
    wire N__54965;
    wire N__54964;
    wire N__54963;
    wire N__54962;
    wire N__54961;
    wire N__54960;
    wire N__54955;
    wire N__54954;
    wire N__54953;
    wire N__54950;
    wire N__54949;
    wire N__54948;
    wire N__54947;
    wire N__54946;
    wire N__54945;
    wire N__54932;
    wire N__54929;
    wire N__54924;
    wire N__54923;
    wire N__54922;
    wire N__54917;
    wire N__54914;
    wire N__54913;
    wire N__54912;
    wire N__54911;
    wire N__54908;
    wire N__54907;
    wire N__54904;
    wire N__54903;
    wire N__54902;
    wire N__54901;
    wire N__54900;
    wire N__54899;
    wire N__54896;
    wire N__54895;
    wire N__54894;
    wire N__54893;
    wire N__54892;
    wire N__54891;
    wire N__54890;
    wire N__54889;
    wire N__54888;
    wire N__54887;
    wire N__54884;
    wire N__54879;
    wire N__54872;
    wire N__54871;
    wire N__54870;
    wire N__54869;
    wire N__54868;
    wire N__54867;
    wire N__54864;
    wire N__54859;
    wire N__54854;
    wire N__54851;
    wire N__54848;
    wire N__54847;
    wire N__54846;
    wire N__54843;
    wire N__54838;
    wire N__54837;
    wire N__54836;
    wire N__54833;
    wire N__54830;
    wire N__54829;
    wire N__54828;
    wire N__54825;
    wire N__54824;
    wire N__54823;
    wire N__54818;
    wire N__54811;
    wire N__54810;
    wire N__54809;
    wire N__54808;
    wire N__54807;
    wire N__54806;
    wire N__54805;
    wire N__54804;
    wire N__54803;
    wire N__54796;
    wire N__54785;
    wire N__54776;
    wire N__54773;
    wire N__54766;
    wire N__54765;
    wire N__54764;
    wire N__54763;
    wire N__54758;
    wire N__54751;
    wire N__54740;
    wire N__54737;
    wire N__54736;
    wire N__54735;
    wire N__54732;
    wire N__54727;
    wire N__54724;
    wire N__54723;
    wire N__54722;
    wire N__54719;
    wire N__54718;
    wire N__54717;
    wire N__54714;
    wire N__54711;
    wire N__54710;
    wire N__54709;
    wire N__54708;
    wire N__54707;
    wire N__54706;
    wire N__54705;
    wire N__54700;
    wire N__54697;
    wire N__54694;
    wire N__54691;
    wire N__54686;
    wire N__54677;
    wire N__54668;
    wire N__54661;
    wire N__54656;
    wire N__54655;
    wire N__54654;
    wire N__54649;
    wire N__54646;
    wire N__54641;
    wire N__54638;
    wire N__54637;
    wire N__54636;
    wire N__54635;
    wire N__54632;
    wire N__54629;
    wire N__54626;
    wire N__54621;
    wire N__54616;
    wire N__54613;
    wire N__54610;
    wire N__54605;
    wire N__54600;
    wire N__54593;
    wire N__54588;
    wire N__54585;
    wire N__54580;
    wire N__54577;
    wire N__54566;
    wire N__54563;
    wire N__54560;
    wire N__54559;
    wire N__54558;
    wire N__54555;
    wire N__54548;
    wire N__54545;
    wire N__54538;
    wire N__54537;
    wire N__54534;
    wire N__54531;
    wire N__54530;
    wire N__54529;
    wire N__54528;
    wire N__54525;
    wire N__54522;
    wire N__54507;
    wire N__54496;
    wire N__54493;
    wire N__54488;
    wire N__54479;
    wire N__54476;
    wire N__54471;
    wire N__54468;
    wire N__54463;
    wire N__54456;
    wire N__54453;
    wire N__54446;
    wire N__54431;
    wire N__54428;
    wire N__54425;
    wire N__54422;
    wire N__54419;
    wire N__54416;
    wire N__54413;
    wire N__54410;
    wire N__54407;
    wire N__54404;
    wire N__54401;
    wire N__54398;
    wire N__54395;
    wire N__54392;
    wire N__54389;
    wire N__54386;
    wire N__54383;
    wire N__54382;
    wire N__54381;
    wire N__54380;
    wire N__54379;
    wire N__54378;
    wire N__54375;
    wire N__54374;
    wire N__54373;
    wire N__54372;
    wire N__54371;
    wire N__54370;
    wire N__54369;
    wire N__54368;
    wire N__54367;
    wire N__54356;
    wire N__54353;
    wire N__54352;
    wire N__54351;
    wire N__54348;
    wire N__54347;
    wire N__54346;
    wire N__54345;
    wire N__54344;
    wire N__54343;
    wire N__54332;
    wire N__54331;
    wire N__54330;
    wire N__54329;
    wire N__54328;
    wire N__54327;
    wire N__54324;
    wire N__54321;
    wire N__54320;
    wire N__54319;
    wire N__54318;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54308;
    wire N__54303;
    wire N__54298;
    wire N__54291;
    wire N__54290;
    wire N__54289;
    wire N__54288;
    wire N__54287;
    wire N__54284;
    wire N__54273;
    wire N__54272;
    wire N__54271;
    wire N__54270;
    wire N__54269;
    wire N__54266;
    wire N__54257;
    wire N__54254;
    wire N__54249;
    wire N__54246;
    wire N__54239;
    wire N__54230;
    wire N__54225;
    wire N__54216;
    wire N__54207;
    wire N__54204;
    wire N__54191;
    wire N__54188;
    wire N__54185;
    wire N__54182;
    wire N__54179;
    wire N__54178;
    wire N__54177;
    wire N__54176;
    wire N__54175;
    wire N__54174;
    wire N__54173;
    wire N__54172;
    wire N__54171;
    wire N__54170;
    wire N__54169;
    wire N__54168;
    wire N__54167;
    wire N__54166;
    wire N__54165;
    wire N__54164;
    wire N__54151;
    wire N__54150;
    wire N__54149;
    wire N__54146;
    wire N__54145;
    wire N__54142;
    wire N__54141;
    wire N__54140;
    wire N__54139;
    wire N__54138;
    wire N__54137;
    wire N__54136;
    wire N__54133;
    wire N__54130;
    wire N__54129;
    wire N__54128;
    wire N__54125;
    wire N__54124;
    wire N__54113;
    wire N__54110;
    wire N__54107;
    wire N__54106;
    wire N__54095;
    wire N__54092;
    wire N__54091;
    wire N__54090;
    wire N__54089;
    wire N__54088;
    wire N__54087;
    wire N__54086;
    wire N__54085;
    wire N__54084;
    wire N__54083;
    wire N__54082;
    wire N__54081;
    wire N__54080;
    wire N__54079;
    wire N__54078;
    wire N__54077;
    wire N__54076;
    wire N__54075;
    wire N__54074;
    wire N__54073;
    wire N__54072;
    wire N__54071;
    wire N__54070;
    wire N__54069;
    wire N__54068;
    wire N__54067;
    wire N__54064;
    wire N__54057;
    wire N__54056;
    wire N__54055;
    wire N__54054;
    wire N__54053;
    wire N__54052;
    wire N__54051;
    wire N__54048;
    wire N__54045;
    wire N__54040;
    wire N__54037;
    wire N__54036;
    wire N__54035;
    wire N__54034;
    wire N__54033;
    wire N__54032;
    wire N__54031;
    wire N__54030;
    wire N__54029;
    wire N__54028;
    wire N__54027;
    wire N__54026;
    wire N__54023;
    wire N__54022;
    wire N__54015;
    wire N__54012;
    wire N__54009;
    wire N__54008;
    wire N__54007;
    wire N__54006;
    wire N__54005;
    wire N__53998;
    wire N__53997;
    wire N__53996;
    wire N__53995;
    wire N__53994;
    wire N__53991;
    wire N__53988;
    wire N__53985;
    wire N__53982;
    wire N__53965;
    wire N__53964;
    wire N__53963;
    wire N__53960;
    wire N__53959;
    wire N__53958;
    wire N__53957;
    wire N__53956;
    wire N__53955;
    wire N__53952;
    wire N__53951;
    wire N__53950;
    wire N__53947;
    wire N__53930;
    wire N__53925;
    wire N__53922;
    wire N__53921;
    wire N__53918;
    wire N__53917;
    wire N__53914;
    wire N__53911;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53895;
    wire N__53892;
    wire N__53885;
    wire N__53878;
    wire N__53875;
    wire N__53872;
    wire N__53869;
    wire N__53866;
    wire N__53863;
    wire N__53862;
    wire N__53859;
    wire N__53856;
    wire N__53851;
    wire N__53844;
    wire N__53843;
    wire N__53842;
    wire N__53839;
    wire N__53836;
    wire N__53829;
    wire N__53826;
    wire N__53817;
    wire N__53814;
    wire N__53813;
    wire N__53812;
    wire N__53807;
    wire N__53806;
    wire N__53805;
    wire N__53804;
    wire N__53801;
    wire N__53794;
    wire N__53789;
    wire N__53788;
    wire N__53787;
    wire N__53786;
    wire N__53783;
    wire N__53778;
    wire N__53775;
    wire N__53774;
    wire N__53773;
    wire N__53772;
    wire N__53771;
    wire N__53770;
    wire N__53765;
    wire N__53760;
    wire N__53757;
    wire N__53754;
    wire N__53741;
    wire N__53732;
    wire N__53729;
    wire N__53722;
    wire N__53719;
    wire N__53710;
    wire N__53705;
    wire N__53698;
    wire N__53691;
    wire N__53686;
    wire N__53683;
    wire N__53676;
    wire N__53669;
    wire N__53662;
    wire N__53655;
    wire N__53650;
    wire N__53643;
    wire N__53628;
    wire N__53621;
    wire N__53616;
    wire N__53591;
    wire N__53590;
    wire N__53589;
    wire N__53588;
    wire N__53587;
    wire N__53586;
    wire N__53583;
    wire N__53582;
    wire N__53581;
    wire N__53572;
    wire N__53569;
    wire N__53568;
    wire N__53567;
    wire N__53566;
    wire N__53565;
    wire N__53564;
    wire N__53563;
    wire N__53562;
    wire N__53561;
    wire N__53558;
    wire N__53555;
    wire N__53554;
    wire N__53553;
    wire N__53550;
    wire N__53549;
    wire N__53548;
    wire N__53545;
    wire N__53542;
    wire N__53539;
    wire N__53538;
    wire N__53537;
    wire N__53534;
    wire N__53531;
    wire N__53524;
    wire N__53521;
    wire N__53520;
    wire N__53519;
    wire N__53518;
    wire N__53517;
    wire N__53516;
    wire N__53513;
    wire N__53510;
    wire N__53507;
    wire N__53506;
    wire N__53505;
    wire N__53504;
    wire N__53503;
    wire N__53498;
    wire N__53497;
    wire N__53496;
    wire N__53495;
    wire N__53492;
    wire N__53489;
    wire N__53486;
    wire N__53479;
    wire N__53474;
    wire N__53471;
    wire N__53468;
    wire N__53467;
    wire N__53466;
    wire N__53465;
    wire N__53460;
    wire N__53455;
    wire N__53448;
    wire N__53443;
    wire N__53440;
    wire N__53435;
    wire N__53430;
    wire N__53427;
    wire N__53420;
    wire N__53417;
    wire N__53414;
    wire N__53411;
    wire N__53408;
    wire N__53405;
    wire N__53400;
    wire N__53393;
    wire N__53386;
    wire N__53383;
    wire N__53364;
    wire N__53351;
    wire N__53350;
    wire N__53347;
    wire N__53346;
    wire N__53341;
    wire N__53338;
    wire N__53333;
    wire N__53330;
    wire N__53327;
    wire N__53326;
    wire N__53325;
    wire N__53324;
    wire N__53321;
    wire N__53318;
    wire N__53313;
    wire N__53306;
    wire N__53303;
    wire N__53300;
    wire N__53297;
    wire N__53296;
    wire N__53295;
    wire N__53292;
    wire N__53289;
    wire N__53286;
    wire N__53279;
    wire N__53278;
    wire N__53277;
    wire N__53274;
    wire N__53271;
    wire N__53268;
    wire N__53265;
    wire N__53260;
    wire N__53255;
    wire N__53254;
    wire N__53251;
    wire N__53250;
    wire N__53247;
    wire N__53242;
    wire N__53237;
    wire N__53234;
    wire N__53231;
    wire N__53230;
    wire N__53229;
    wire N__53226;
    wire N__53223;
    wire N__53220;
    wire N__53217;
    wire N__53214;
    wire N__53207;
    wire N__53206;
    wire N__53201;
    wire N__53200;
    wire N__53199;
    wire N__53198;
    wire N__53195;
    wire N__53192;
    wire N__53189;
    wire N__53186;
    wire N__53185;
    wire N__53184;
    wire N__53183;
    wire N__53180;
    wire N__53179;
    wire N__53178;
    wire N__53177;
    wire N__53176;
    wire N__53175;
    wire N__53172;
    wire N__53167;
    wire N__53166;
    wire N__53163;
    wire N__53160;
    wire N__53157;
    wire N__53156;
    wire N__53153;
    wire N__53146;
    wire N__53143;
    wire N__53140;
    wire N__53135;
    wire N__53132;
    wire N__53131;
    wire N__53130;
    wire N__53129;
    wire N__53128;
    wire N__53127;
    wire N__53124;
    wire N__53121;
    wire N__53118;
    wire N__53117;
    wire N__53116;
    wire N__53113;
    wire N__53110;
    wire N__53105;
    wire N__53102;
    wire N__53097;
    wire N__53092;
    wire N__53085;
    wire N__53080;
    wire N__53077;
    wire N__53070;
    wire N__53069;
    wire N__53068;
    wire N__53063;
    wire N__53060;
    wire N__53053;
    wire N__53050;
    wire N__53047;
    wire N__53044;
    wire N__53039;
    wire N__53036;
    wire N__53033;
    wire N__53030;
    wire N__53021;
    wire N__53012;
    wire N__53011;
    wire N__53008;
    wire N__53007;
    wire N__53006;
    wire N__53005;
    wire N__53004;
    wire N__53003;
    wire N__53002;
    wire N__53001;
    wire N__53000;
    wire N__52999;
    wire N__52998;
    wire N__52997;
    wire N__52996;
    wire N__52995;
    wire N__52994;
    wire N__52993;
    wire N__52992;
    wire N__52991;
    wire N__52990;
    wire N__52989;
    wire N__52986;
    wire N__52983;
    wire N__52970;
    wire N__52967;
    wire N__52960;
    wire N__52959;
    wire N__52958;
    wire N__52955;
    wire N__52954;
    wire N__52953;
    wire N__52952;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52937;
    wire N__52936;
    wire N__52935;
    wire N__52934;
    wire N__52933;
    wire N__52930;
    wire N__52927;
    wire N__52924;
    wire N__52917;
    wire N__52916;
    wire N__52915;
    wire N__52912;
    wire N__52911;
    wire N__52908;
    wire N__52903;
    wire N__52900;
    wire N__52891;
    wire N__52886;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52878;
    wire N__52877;
    wire N__52876;
    wire N__52875;
    wire N__52866;
    wire N__52863;
    wire N__52858;
    wire N__52855;
    wire N__52854;
    wire N__52851;
    wire N__52850;
    wire N__52849;
    wire N__52848;
    wire N__52847;
    wire N__52846;
    wire N__52845;
    wire N__52844;
    wire N__52841;
    wire N__52838;
    wire N__52835;
    wire N__52832;
    wire N__52829;
    wire N__52820;
    wire N__52819;
    wire N__52806;
    wire N__52801;
    wire N__52796;
    wire N__52793;
    wire N__52788;
    wire N__52779;
    wire N__52774;
    wire N__52769;
    wire N__52764;
    wire N__52759;
    wire N__52758;
    wire N__52757;
    wire N__52756;
    wire N__52755;
    wire N__52754;
    wire N__52753;
    wire N__52752;
    wire N__52751;
    wire N__52750;
    wire N__52749;
    wire N__52748;
    wire N__52747;
    wire N__52746;
    wire N__52743;
    wire N__52740;
    wire N__52735;
    wire N__52722;
    wire N__52721;
    wire N__52720;
    wire N__52717;
    wire N__52710;
    wire N__52709;
    wire N__52708;
    wire N__52707;
    wire N__52706;
    wire N__52703;
    wire N__52696;
    wire N__52683;
    wire N__52680;
    wire N__52675;
    wire N__52672;
    wire N__52667;
    wire N__52662;
    wire N__52653;
    wire N__52634;
    wire N__52633;
    wire N__52630;
    wire N__52627;
    wire N__52626;
    wire N__52623;
    wire N__52618;
    wire N__52613;
    wire N__52610;
    wire N__52609;
    wire N__52606;
    wire N__52603;
    wire N__52602;
    wire N__52599;
    wire N__52596;
    wire N__52593;
    wire N__52588;
    wire N__52583;
    wire N__52580;
    wire N__52577;
    wire N__52574;
    wire N__52571;
    wire N__52568;
    wire N__52565;
    wire N__52562;
    wire N__52559;
    wire N__52556;
    wire N__52553;
    wire N__52550;
    wire N__52547;
    wire N__52544;
    wire N__52541;
    wire N__52538;
    wire N__52535;
    wire N__52532;
    wire N__52529;
    wire N__52526;
    wire N__52523;
    wire N__52520;
    wire N__52517;
    wire N__52514;
    wire N__52511;
    wire N__52508;
    wire N__52507;
    wire N__52506;
    wire N__52505;
    wire N__52500;
    wire N__52497;
    wire N__52494;
    wire N__52493;
    wire N__52490;
    wire N__52489;
    wire N__52486;
    wire N__52483;
    wire N__52480;
    wire N__52477;
    wire N__52474;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52460;
    wire N__52457;
    wire N__52454;
    wire N__52451;
    wire N__52448;
    wire N__52439;
    wire N__52438;
    wire N__52437;
    wire N__52436;
    wire N__52435;
    wire N__52434;
    wire N__52433;
    wire N__52432;
    wire N__52421;
    wire N__52420;
    wire N__52417;
    wire N__52416;
    wire N__52413;
    wire N__52412;
    wire N__52411;
    wire N__52410;
    wire N__52409;
    wire N__52408;
    wire N__52407;
    wire N__52406;
    wire N__52403;
    wire N__52400;
    wire N__52397;
    wire N__52394;
    wire N__52393;
    wire N__52392;
    wire N__52391;
    wire N__52390;
    wire N__52389;
    wire N__52388;
    wire N__52387;
    wire N__52384;
    wire N__52381;
    wire N__52380;
    wire N__52379;
    wire N__52378;
    wire N__52377;
    wire N__52376;
    wire N__52371;
    wire N__52370;
    wire N__52369;
    wire N__52368;
    wire N__52367;
    wire N__52366;
    wire N__52365;
    wire N__52364;
    wire N__52361;
    wire N__52356;
    wire N__52353;
    wire N__52350;
    wire N__52349;
    wire N__52348;
    wire N__52345;
    wire N__52342;
    wire N__52339;
    wire N__52336;
    wire N__52327;
    wire N__52326;
    wire N__52319;
    wire N__52314;
    wire N__52307;
    wire N__52306;
    wire N__52305;
    wire N__52304;
    wire N__52303;
    wire N__52302;
    wire N__52297;
    wire N__52294;
    wire N__52289;
    wire N__52286;
    wire N__52283;
    wire N__52280;
    wire N__52275;
    wire N__52270;
    wire N__52267;
    wire N__52260;
    wire N__52259;
    wire N__52254;
    wire N__52247;
    wire N__52244;
    wire N__52237;
    wire N__52232;
    wire N__52225;
    wire N__52216;
    wire N__52203;
    wire N__52200;
    wire N__52195;
    wire N__52190;
    wire N__52175;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52160;
    wire N__52157;
    wire N__52154;
    wire N__52153;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52143;
    wire N__52140;
    wire N__52137;
    wire N__52134;
    wire N__52131;
    wire N__52128;
    wire N__52121;
    wire N__52120;
    wire N__52117;
    wire N__52114;
    wire N__52109;
    wire N__52106;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52094;
    wire N__52091;
    wire N__52090;
    wire N__52089;
    wire N__52088;
    wire N__52087;
    wire N__52086;
    wire N__52085;
    wire N__52082;
    wire N__52079;
    wire N__52078;
    wire N__52077;
    wire N__52076;
    wire N__52075;
    wire N__52074;
    wire N__52073;
    wire N__52072;
    wire N__52071;
    wire N__52068;
    wire N__52065;
    wire N__52058;
    wire N__52053;
    wire N__52048;
    wire N__52047;
    wire N__52046;
    wire N__52043;
    wire N__52040;
    wire N__52031;
    wire N__52028;
    wire N__52023;
    wire N__52020;
    wire N__52017;
    wire N__52016;
    wire N__52015;
    wire N__52014;
    wire N__52009;
    wire N__52006;
    wire N__52005;
    wire N__52004;
    wire N__52003;
    wire N__52002;
    wire N__51999;
    wire N__51994;
    wire N__51991;
    wire N__51988;
    wire N__51985;
    wire N__51984;
    wire N__51983;
    wire N__51982;
    wire N__51981;
    wire N__51980;
    wire N__51979;
    wire N__51978;
    wire N__51977;
    wire N__51974;
    wire N__51969;
    wire N__51964;
    wire N__51959;
    wire N__51954;
    wire N__51947;
    wire N__51942;
    wire N__51937;
    wire N__51932;
    wire N__51923;
    wire N__51920;
    wire N__51915;
    wire N__51908;
    wire N__51905;
    wire N__51890;
    wire N__51889;
    wire N__51886;
    wire N__51885;
    wire N__51878;
    wire N__51875;
    wire N__51874;
    wire N__51873;
    wire N__51870;
    wire N__51867;
    wire N__51864;
    wire N__51861;
    wire N__51858;
    wire N__51855;
    wire N__51852;
    wire N__51845;
    wire N__51844;
    wire N__51843;
    wire N__51842;
    wire N__51841;
    wire N__51840;
    wire N__51839;
    wire N__51838;
    wire N__51835;
    wire N__51832;
    wire N__51829;
    wire N__51828;
    wire N__51827;
    wire N__51826;
    wire N__51825;
    wire N__51820;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51804;
    wire N__51801;
    wire N__51794;
    wire N__51789;
    wire N__51786;
    wire N__51783;
    wire N__51782;
    wire N__51777;
    wire N__51774;
    wire N__51767;
    wire N__51766;
    wire N__51763;
    wire N__51762;
    wire N__51759;
    wire N__51756;
    wire N__51753;
    wire N__51748;
    wire N__51747;
    wire N__51746;
    wire N__51745;
    wire N__51742;
    wire N__51741;
    wire N__51738;
    wire N__51735;
    wire N__51732;
    wire N__51729;
    wire N__51724;
    wire N__51717;
    wire N__51714;
    wire N__51703;
    wire N__51700;
    wire N__51697;
    wire N__51692;
    wire N__51691;
    wire N__51690;
    wire N__51689;
    wire N__51688;
    wire N__51683;
    wire N__51680;
    wire N__51677;
    wire N__51674;
    wire N__51673;
    wire N__51672;
    wire N__51671;
    wire N__51670;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51658;
    wire N__51653;
    wire N__51648;
    wire N__51647;
    wire N__51646;
    wire N__51643;
    wire N__51642;
    wire N__51639;
    wire N__51632;
    wire N__51629;
    wire N__51620;
    wire N__51611;
    wire N__51608;
    wire N__51605;
    wire N__51602;
    wire N__51599;
    wire N__51596;
    wire N__51593;
    wire N__51590;
    wire N__51589;
    wire N__51586;
    wire N__51585;
    wire N__51584;
    wire N__51581;
    wire N__51574;
    wire N__51573;
    wire N__51570;
    wire N__51569;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51552;
    wire N__51551;
    wire N__51550;
    wire N__51549;
    wire N__51546;
    wire N__51543;
    wire N__51542;
    wire N__51539;
    wire N__51536;
    wire N__51533;
    wire N__51530;
    wire N__51527;
    wire N__51522;
    wire N__51519;
    wire N__51516;
    wire N__51513;
    wire N__51508;
    wire N__51505;
    wire N__51498;
    wire N__51493;
    wire N__51482;
    wire N__51481;
    wire N__51478;
    wire N__51477;
    wire N__51476;
    wire N__51473;
    wire N__51470;
    wire N__51465;
    wire N__51462;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51446;
    wire N__51443;
    wire N__51442;
    wire N__51439;
    wire N__51436;
    wire N__51435;
    wire N__51432;
    wire N__51429;
    wire N__51426;
    wire N__51423;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51407;
    wire N__51406;
    wire N__51405;
    wire N__51402;
    wire N__51399;
    wire N__51398;
    wire N__51395;
    wire N__51394;
    wire N__51393;
    wire N__51390;
    wire N__51387;
    wire N__51384;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51362;
    wire N__51359;
    wire N__51356;
    wire N__51353;
    wire N__51350;
    wire N__51343;
    wire N__51342;
    wire N__51335;
    wire N__51330;
    wire N__51327;
    wire N__51320;
    wire N__51319;
    wire N__51314;
    wire N__51313;
    wire N__51312;
    wire N__51311;
    wire N__51308;
    wire N__51303;
    wire N__51300;
    wire N__51299;
    wire N__51298;
    wire N__51293;
    wire N__51290;
    wire N__51285;
    wire N__51284;
    wire N__51281;
    wire N__51276;
    wire N__51273;
    wire N__51266;
    wire N__51265;
    wire N__51262;
    wire N__51259;
    wire N__51254;
    wire N__51251;
    wire N__51248;
    wire N__51245;
    wire N__51242;
    wire N__51239;
    wire N__51236;
    wire N__51233;
    wire N__51230;
    wire N__51227;
    wire N__51224;
    wire N__51221;
    wire N__51218;
    wire N__51215;
    wire N__51212;
    wire N__51209;
    wire N__51208;
    wire N__51205;
    wire N__51202;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51187;
    wire N__51184;
    wire N__51183;
    wire N__51182;
    wire N__51181;
    wire N__51178;
    wire N__51175;
    wire N__51172;
    wire N__51169;
    wire N__51168;
    wire N__51165;
    wire N__51162;
    wire N__51157;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51124;
    wire N__51119;
    wire N__51118;
    wire N__51115;
    wire N__51112;
    wire N__51109;
    wire N__51106;
    wire N__51103;
    wire N__51100;
    wire N__51095;
    wire N__51094;
    wire N__51091;
    wire N__51088;
    wire N__51085;
    wire N__51082;
    wire N__51077;
    wire N__51076;
    wire N__51073;
    wire N__51070;
    wire N__51067;
    wire N__51064;
    wire N__51059;
    wire N__51056;
    wire N__51055;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51047;
    wire N__51044;
    wire N__51043;
    wire N__51042;
    wire N__51039;
    wire N__51036;
    wire N__51033;
    wire N__51032;
    wire N__51029;
    wire N__51026;
    wire N__51023;
    wire N__51018;
    wire N__51015;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51003;
    wire N__50996;
    wire N__50995;
    wire N__50994;
    wire N__50989;
    wire N__50984;
    wire N__50981;
    wire N__50978;
    wire N__50969;
    wire N__50968;
    wire N__50965;
    wire N__50960;
    wire N__50957;
    wire N__50954;
    wire N__50951;
    wire N__50948;
    wire N__50945;
    wire N__50942;
    wire N__50939;
    wire N__50936;
    wire N__50933;
    wire N__50932;
    wire N__50931;
    wire N__50930;
    wire N__50927;
    wire N__50926;
    wire N__50925;
    wire N__50922;
    wire N__50917;
    wire N__50914;
    wire N__50911;
    wire N__50908;
    wire N__50907;
    wire N__50906;
    wire N__50903;
    wire N__50898;
    wire N__50895;
    wire N__50892;
    wire N__50887;
    wire N__50886;
    wire N__50885;
    wire N__50882;
    wire N__50879;
    wire N__50872;
    wire N__50867;
    wire N__50858;
    wire N__50855;
    wire N__50854;
    wire N__50851;
    wire N__50850;
    wire N__50847;
    wire N__50844;
    wire N__50841;
    wire N__50834;
    wire N__50831;
    wire N__50828;
    wire N__50825;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50813;
    wire N__50810;
    wire N__50807;
    wire N__50804;
    wire N__50801;
    wire N__50798;
    wire N__50795;
    wire N__50792;
    wire N__50789;
    wire N__50786;
    wire N__50783;
    wire N__50782;
    wire N__50779;
    wire N__50778;
    wire N__50777;
    wire N__50776;
    wire N__50775;
    wire N__50772;
    wire N__50771;
    wire N__50768;
    wire N__50765;
    wire N__50762;
    wire N__50761;
    wire N__50758;
    wire N__50755;
    wire N__50752;
    wire N__50749;
    wire N__50742;
    wire N__50739;
    wire N__50736;
    wire N__50733;
    wire N__50728;
    wire N__50723;
    wire N__50720;
    wire N__50715;
    wire N__50712;
    wire N__50705;
    wire N__50702;
    wire N__50701;
    wire N__50698;
    wire N__50695;
    wire N__50692;
    wire N__50687;
    wire N__50686;
    wire N__50685;
    wire N__50684;
    wire N__50683;
    wire N__50682;
    wire N__50681;
    wire N__50680;
    wire N__50679;
    wire N__50678;
    wire N__50671;
    wire N__50670;
    wire N__50669;
    wire N__50668;
    wire N__50667;
    wire N__50666;
    wire N__50665;
    wire N__50664;
    wire N__50663;
    wire N__50662;
    wire N__50659;
    wire N__50652;
    wire N__50645;
    wire N__50642;
    wire N__50637;
    wire N__50636;
    wire N__50633;
    wire N__50632;
    wire N__50631;
    wire N__50626;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50604;
    wire N__50601;
    wire N__50598;
    wire N__50593;
    wire N__50590;
    wire N__50585;
    wire N__50580;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50558;
    wire N__50555;
    wire N__50554;
    wire N__50553;
    wire N__50552;
    wire N__50549;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50545;
    wire N__50544;
    wire N__50539;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50535;
    wire N__50534;
    wire N__50533;
    wire N__50532;
    wire N__50529;
    wire N__50526;
    wire N__50523;
    wire N__50518;
    wire N__50513;
    wire N__50510;
    wire N__50507;
    wire N__50506;
    wire N__50499;
    wire N__50496;
    wire N__50495;
    wire N__50494;
    wire N__50493;
    wire N__50488;
    wire N__50485;
    wire N__50484;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50478;
    wire N__50475;
    wire N__50466;
    wire N__50463;
    wire N__50458;
    wire N__50451;
    wire N__50448;
    wire N__50445;
    wire N__50436;
    wire N__50429;
    wire N__50414;
    wire N__50411;
    wire N__50408;
    wire N__50405;
    wire N__50402;
    wire N__50399;
    wire N__50396;
    wire N__50393;
    wire N__50390;
    wire N__50387;
    wire N__50384;
    wire N__50381;
    wire N__50380;
    wire N__50377;
    wire N__50374;
    wire N__50371;
    wire N__50366;
    wire N__50363;
    wire N__50362;
    wire N__50361;
    wire N__50360;
    wire N__50359;
    wire N__50358;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50350;
    wire N__50349;
    wire N__50346;
    wire N__50343;
    wire N__50340;
    wire N__50337;
    wire N__50334;
    wire N__50329;
    wire N__50324;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50296;
    wire N__50295;
    wire N__50278;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50255;
    wire N__50254;
    wire N__50251;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50243;
    wire N__50240;
    wire N__50237;
    wire N__50234;
    wire N__50233;
    wire N__50230;
    wire N__50225;
    wire N__50224;
    wire N__50223;
    wire N__50220;
    wire N__50213;
    wire N__50210;
    wire N__50205;
    wire N__50200;
    wire N__50197;
    wire N__50186;
    wire N__50185;
    wire N__50184;
    wire N__50183;
    wire N__50182;
    wire N__50181;
    wire N__50180;
    wire N__50179;
    wire N__50178;
    wire N__50177;
    wire N__50176;
    wire N__50173;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50139;
    wire N__50138;
    wire N__50137;
    wire N__50134;
    wire N__50133;
    wire N__50132;
    wire N__50131;
    wire N__50130;
    wire N__50127;
    wire N__50124;
    wire N__50121;
    wire N__50116;
    wire N__50099;
    wire N__50098;
    wire N__50095;
    wire N__50092;
    wire N__50087;
    wire N__50086;
    wire N__50085;
    wire N__50084;
    wire N__50083;
    wire N__50082;
    wire N__50077;
    wire N__50074;
    wire N__50071;
    wire N__50064;
    wire N__50057;
    wire N__50052;
    wire N__50039;
    wire N__50036;
    wire N__50033;
    wire N__50030;
    wire N__50027;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50014;
    wire N__50009;
    wire N__50006;
    wire N__50003;
    wire N__50002;
    wire N__49999;
    wire N__49998;
    wire N__49995;
    wire N__49992;
    wire N__49989;
    wire N__49986;
    wire N__49979;
    wire N__49978;
    wire N__49975;
    wire N__49972;
    wire N__49971;
    wire N__49968;
    wire N__49965;
    wire N__49962;
    wire N__49959;
    wire N__49952;
    wire N__49949;
    wire N__49946;
    wire N__49943;
    wire N__49940;
    wire N__49937;
    wire N__49934;
    wire N__49931;
    wire N__49928;
    wire N__49925;
    wire N__49924;
    wire N__49923;
    wire N__49922;
    wire N__49921;
    wire N__49920;
    wire N__49919;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49915;
    wire N__49914;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49905;
    wire N__49904;
    wire N__49901;
    wire N__49900;
    wire N__49899;
    wire N__49898;
    wire N__49897;
    wire N__49896;
    wire N__49895;
    wire N__49890;
    wire N__49887;
    wire N__49882;
    wire N__49879;
    wire N__49876;
    wire N__49875;
    wire N__49872;
    wire N__49871;
    wire N__49868;
    wire N__49861;
    wire N__49856;
    wire N__49849;
    wire N__49840;
    wire N__49839;
    wire N__49838;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49828;
    wire N__49827;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49823;
    wire N__49820;
    wire N__49815;
    wire N__49810;
    wire N__49803;
    wire N__49792;
    wire N__49785;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49768;
    wire N__49767;
    wire N__49762;
    wire N__49759;
    wire N__49758;
    wire N__49755;
    wire N__49754;
    wire N__49751;
    wire N__49750;
    wire N__49749;
    wire N__49746;
    wire N__49743;
    wire N__49740;
    wire N__49739;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49721;
    wire N__49720;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49708;
    wire N__49705;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49699;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49691;
    wire N__49688;
    wire N__49687;
    wire N__49686;
    wire N__49683;
    wire N__49682;
    wire N__49679;
    wire N__49674;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49664;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49652;
    wire N__49647;
    wire N__49642;
    wire N__49639;
    wire N__49638;
    wire N__49631;
    wire N__49630;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49626;
    wire N__49623;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49605;
    wire N__49602;
    wire N__49599;
    wire N__49596;
    wire N__49595;
    wire N__49594;
    wire N__49593;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49587;
    wire N__49576;
    wire N__49569;
    wire N__49562;
    wire N__49555;
    wire N__49548;
    wire N__49539;
    wire N__49536;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49509;
    wire N__49506;
    wire N__49497;
    wire N__49492;
    wire N__49489;
    wire N__49482;
    wire N__49473;
    wire N__49462;
    wire N__49457;
    wire N__49450;
    wire N__49449;
    wire N__49448;
    wire N__49445;
    wire N__49436;
    wire N__49433;
    wire N__49428;
    wire N__49423;
    wire N__49418;
    wire N__49407;
    wire N__49404;
    wire N__49401;
    wire N__49396;
    wire N__49389;
    wire N__49384;
    wire N__49373;
    wire N__49372;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49368;
    wire N__49367;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49359;
    wire N__49358;
    wire N__49357;
    wire N__49356;
    wire N__49345;
    wire N__49344;
    wire N__49343;
    wire N__49342;
    wire N__49339;
    wire N__49336;
    wire N__49333;
    wire N__49326;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49312;
    wire N__49309;
    wire N__49306;
    wire N__49303;
    wire N__49296;
    wire N__49283;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49275;
    wire N__49272;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49253;
    wire N__49250;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49237;
    wire N__49234;
    wire N__49229;
    wire N__49226;
    wire N__49225;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49205;
    wire N__49202;
    wire N__49199;
    wire N__49196;
    wire N__49193;
    wire N__49190;
    wire N__49187;
    wire N__49184;
    wire N__49181;
    wire N__49180;
    wire N__49177;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49162;
    wire N__49157;
    wire N__49154;
    wire N__49153;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49117;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49107;
    wire N__49106;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49101;
    wire N__49100;
    wire N__49099;
    wire N__49098;
    wire N__49095;
    wire N__49092;
    wire N__49089;
    wire N__49086;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49074;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49059;
    wire N__49058;
    wire N__49057;
    wire N__49056;
    wire N__49055;
    wire N__49054;
    wire N__49053;
    wire N__49052;
    wire N__49051;
    wire N__49050;
    wire N__49049;
    wire N__49046;
    wire N__49039;
    wire N__49030;
    wire N__49021;
    wire N__49014;
    wire N__49013;
    wire N__49012;
    wire N__49011;
    wire N__49010;
    wire N__49007;
    wire N__49004;
    wire N__49003;
    wire N__49000;
    wire N__48999;
    wire N__48998;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48984;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48966;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48954;
    wire N__48953;
    wire N__48952;
    wire N__48951;
    wire N__48946;
    wire N__48941;
    wire N__48938;
    wire N__48935;
    wire N__48928;
    wire N__48919;
    wire N__48916;
    wire N__48911;
    wire N__48906;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48887;
    wire N__48880;
    wire N__48877;
    wire N__48876;
    wire N__48875;
    wire N__48874;
    wire N__48873;
    wire N__48870;
    wire N__48865;
    wire N__48860;
    wire N__48857;
    wire N__48856;
    wire N__48853;
    wire N__48846;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48826;
    wire N__48817;
    wire N__48816;
    wire N__48815;
    wire N__48810;
    wire N__48807;
    wire N__48804;
    wire N__48795;
    wire N__48786;
    wire N__48783;
    wire N__48776;
    wire N__48767;
    wire N__48762;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48740;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48735;
    wire N__48734;
    wire N__48731;
    wire N__48730;
    wire N__48729;
    wire N__48728;
    wire N__48727;
    wire N__48724;
    wire N__48723;
    wire N__48720;
    wire N__48719;
    wire N__48718;
    wire N__48715;
    wire N__48714;
    wire N__48709;
    wire N__48704;
    wire N__48703;
    wire N__48702;
    wire N__48701;
    wire N__48700;
    wire N__48697;
    wire N__48692;
    wire N__48689;
    wire N__48688;
    wire N__48687;
    wire N__48686;
    wire N__48685;
    wire N__48682;
    wire N__48681;
    wire N__48678;
    wire N__48677;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48669;
    wire N__48668;
    wire N__48665;
    wire N__48662;
    wire N__48659;
    wire N__48656;
    wire N__48653;
    wire N__48650;
    wire N__48645;
    wire N__48642;
    wire N__48639;
    wire N__48636;
    wire N__48633;
    wire N__48626;
    wire N__48621;
    wire N__48620;
    wire N__48619;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48607;
    wire N__48602;
    wire N__48599;
    wire N__48598;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48585;
    wire N__48578;
    wire N__48575;
    wire N__48574;
    wire N__48569;
    wire N__48564;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48533;
    wire N__48528;
    wire N__48523;
    wire N__48518;
    wire N__48515;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48503;
    wire N__48496;
    wire N__48493;
    wire N__48488;
    wire N__48485;
    wire N__48482;
    wire N__48477;
    wire N__48468;
    wire N__48465;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48440;
    wire N__48425;
    wire N__48424;
    wire N__48423;
    wire N__48420;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48408;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48398;
    wire N__48395;
    wire N__48388;
    wire N__48385;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48377;
    wire N__48376;
    wire N__48375;
    wire N__48374;
    wire N__48373;
    wire N__48372;
    wire N__48371;
    wire N__48370;
    wire N__48369;
    wire N__48366;
    wire N__48365;
    wire N__48364;
    wire N__48363;
    wire N__48362;
    wire N__48361;
    wire N__48360;
    wire N__48359;
    wire N__48354;
    wire N__48351;
    wire N__48348;
    wire N__48345;
    wire N__48344;
    wire N__48343;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48339;
    wire N__48338;
    wire N__48337;
    wire N__48336;
    wire N__48335;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48318;
    wire N__48317;
    wire N__48316;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48312;
    wire N__48311;
    wire N__48310;
    wire N__48309;
    wire N__48308;
    wire N__48305;
    wire N__48300;
    wire N__48299;
    wire N__48298;
    wire N__48297;
    wire N__48296;
    wire N__48295;
    wire N__48294;
    wire N__48293;
    wire N__48292;
    wire N__48289;
    wire N__48286;
    wire N__48285;
    wire N__48278;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48266;
    wire N__48259;
    wire N__48256;
    wire N__48253;
    wire N__48248;
    wire N__48243;
    wire N__48236;
    wire N__48233;
    wire N__48232;
    wire N__48229;
    wire N__48228;
    wire N__48223;
    wire N__48218;
    wire N__48217;
    wire N__48216;
    wire N__48215;
    wire N__48212;
    wire N__48203;
    wire N__48196;
    wire N__48195;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48180;
    wire N__48177;
    wire N__48172;
    wire N__48171;
    wire N__48170;
    wire N__48167;
    wire N__48164;
    wire N__48161;
    wire N__48154;
    wire N__48153;
    wire N__48152;
    wire N__48151;
    wire N__48148;
    wire N__48141;
    wire N__48136;
    wire N__48133;
    wire N__48128;
    wire N__48123;
    wire N__48120;
    wire N__48117;
    wire N__48114;
    wire N__48111;
    wire N__48102;
    wire N__48099;
    wire N__48098;
    wire N__48095;
    wire N__48094;
    wire N__48091;
    wire N__48090;
    wire N__48085;
    wire N__48078;
    wire N__48073;
    wire N__48070;
    wire N__48065;
    wire N__48054;
    wire N__48051;
    wire N__48046;
    wire N__48037;
    wire N__48030;
    wire N__48027;
    wire N__48024;
    wire N__48021;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__47999;
    wire N__47998;
    wire N__47997;
    wire N__47994;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47975;
    wire N__47970;
    wire N__47961;
    wire N__47950;
    wire N__47943;
    wire N__47938;
    wire N__47915;
    wire N__47912;
    wire N__47911;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47887;
    wire N__47884;
    wire N__47881;
    wire N__47876;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47866;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47851;
    wire N__47848;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47832;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47818;
    wire N__47815;
    wire N__47812;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47795;
    wire N__47794;
    wire N__47791;
    wire N__47788;
    wire N__47787;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47773;
    wire N__47770;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47752;
    wire N__47749;
    wire N__47746;
    wire N__47745;
    wire N__47740;
    wire N__47737;
    wire N__47732;
    wire N__47731;
    wire N__47730;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47697;
    wire N__47692;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47680;
    wire N__47677;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47669;
    wire N__47666;
    wire N__47663;
    wire N__47660;
    wire N__47657;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47634;
    wire N__47631;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47621;
    wire N__47618;
    wire N__47613;
    wire N__47606;
    wire N__47603;
    wire N__47600;
    wire N__47597;
    wire N__47594;
    wire N__47591;
    wire N__47588;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47576;
    wire N__47575;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47560;
    wire N__47555;
    wire N__47552;
    wire N__47551;
    wire N__47548;
    wire N__47547;
    wire N__47544;
    wire N__47541;
    wire N__47538;
    wire N__47531;
    wire N__47530;
    wire N__47527;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47510;
    wire N__47507;
    wire N__47506;
    wire N__47503;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47486;
    wire N__47485;
    wire N__47482;
    wire N__47479;
    wire N__47476;
    wire N__47471;
    wire N__47468;
    wire N__47465;
    wire N__47462;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47452;
    wire N__47449;
    wire N__47446;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47432;
    wire N__47429;
    wire N__47428;
    wire N__47427;
    wire N__47424;
    wire N__47419;
    wire N__47414;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47406;
    wire N__47401;
    wire N__47398;
    wire N__47397;
    wire N__47396;
    wire N__47395;
    wire N__47392;
    wire N__47389;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47377;
    wire N__47376;
    wire N__47375;
    wire N__47372;
    wire N__47367;
    wire N__47358;
    wire N__47351;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47339;
    wire N__47336;
    wire N__47327;
    wire N__47326;
    wire N__47323;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47296;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47284;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47263;
    wire N__47260;
    wire N__47255;
    wire N__47252;
    wire N__47249;
    wire N__47248;
    wire N__47247;
    wire N__47246;
    wire N__47243;
    wire N__47242;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47234;
    wire N__47231;
    wire N__47228;
    wire N__47225;
    wire N__47222;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47212;
    wire N__47209;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47153;
    wire N__47150;
    wire N__47147;
    wire N__47144;
    wire N__47143;
    wire N__47140;
    wire N__47139;
    wire N__47136;
    wire N__47135;
    wire N__47134;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47124;
    wire N__47121;
    wire N__47118;
    wire N__47115;
    wire N__47110;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47096;
    wire N__47093;
    wire N__47090;
    wire N__47087;
    wire N__47084;
    wire N__47075;
    wire N__47072;
    wire N__47071;
    wire N__47070;
    wire N__47069;
    wire N__47068;
    wire N__47065;
    wire N__47062;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47054;
    wire N__47053;
    wire N__47050;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47029;
    wire N__47022;
    wire N__47015;
    wire N__47012;
    wire N__47009;
    wire N__47000;
    wire N__46997;
    wire N__46996;
    wire N__46995;
    wire N__46994;
    wire N__46993;
    wire N__46990;
    wire N__46989;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46970;
    wire N__46969;
    wire N__46966;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46952;
    wire N__46949;
    wire N__46946;
    wire N__46941;
    wire N__46936;
    wire N__46933;
    wire N__46930;
    wire N__46927;
    wire N__46916;
    wire N__46913;
    wire N__46910;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46880;
    wire N__46877;
    wire N__46874;
    wire N__46871;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46850;
    wire N__46849;
    wire N__46846;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46823;
    wire N__46820;
    wire N__46817;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46799;
    wire N__46796;
    wire N__46795;
    wire N__46792;
    wire N__46789;
    wire N__46786;
    wire N__46783;
    wire N__46780;
    wire N__46777;
    wire N__46772;
    wire N__46769;
    wire N__46768;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46752;
    wire N__46745;
    wire N__46744;
    wire N__46741;
    wire N__46740;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46724;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46694;
    wire N__46691;
    wire N__46690;
    wire N__46689;
    wire N__46686;
    wire N__46681;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46667;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46649;
    wire N__46646;
    wire N__46643;
    wire N__46642;
    wire N__46639;
    wire N__46636;
    wire N__46635;
    wire N__46630;
    wire N__46627;
    wire N__46624;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46609;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46586;
    wire N__46585;
    wire N__46582;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46571;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46555;
    wire N__46550;
    wire N__46547;
    wire N__46544;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46532;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46522;
    wire N__46521;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46499;
    wire N__46496;
    wire N__46493;
    wire N__46492;
    wire N__46491;
    wire N__46488;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46469;
    wire N__46466;
    wire N__46465;
    wire N__46462;
    wire N__46461;
    wire N__46458;
    wire N__46455;
    wire N__46450;
    wire N__46445;
    wire N__46442;
    wire N__46439;
    wire N__46436;
    wire N__46433;
    wire N__46430;
    wire N__46427;
    wire N__46424;
    wire N__46421;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46410;
    wire N__46407;
    wire N__46406;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46379;
    wire N__46376;
    wire N__46371;
    wire N__46368;
    wire N__46367;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46355;
    wire N__46352;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46336;
    wire N__46331;
    wire N__46328;
    wire N__46325;
    wire N__46324;
    wire N__46323;
    wire N__46320;
    wire N__46315;
    wire N__46310;
    wire N__46309;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46299;
    wire N__46292;
    wire N__46289;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46262;
    wire N__46259;
    wire N__46256;
    wire N__46253;
    wire N__46250;
    wire N__46247;
    wire N__46244;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46226;
    wire N__46223;
    wire N__46220;
    wire N__46219;
    wire N__46218;
    wire N__46215;
    wire N__46214;
    wire N__46213;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46205;
    wire N__46202;
    wire N__46199;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46161;
    wire N__46156;
    wire N__46149;
    wire N__46142;
    wire N__46141;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46133;
    wire N__46132;
    wire N__46129;
    wire N__46126;
    wire N__46123;
    wire N__46120;
    wire N__46117;
    wire N__46116;
    wire N__46115;
    wire N__46112;
    wire N__46103;
    wire N__46100;
    wire N__46097;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46085;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46067;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46059;
    wire N__46058;
    wire N__46055;
    wire N__46052;
    wire N__46049;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46032;
    wire N__46029;
    wire N__46028;
    wire N__46025;
    wire N__46022;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45997;
    wire N__45994;
    wire N__45991;
    wire N__45986;
    wire N__45983;
    wire N__45978;
    wire N__45975;
    wire N__45970;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45956;
    wire N__45953;
    wire N__45950;
    wire N__45947;
    wire N__45944;
    wire N__45941;
    wire N__45938;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45916;
    wire N__45913;
    wire N__45912;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45893;
    wire N__45890;
    wire N__45887;
    wire N__45886;
    wire N__45883;
    wire N__45880;
    wire N__45877;
    wire N__45874;
    wire N__45871;
    wire N__45868;
    wire N__45863;
    wire N__45854;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45820;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45800;
    wire N__45799;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45776;
    wire N__45773;
    wire N__45770;
    wire N__45767;
    wire N__45764;
    wire N__45761;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45749;
    wire N__45746;
    wire N__45743;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45719;
    wire N__45716;
    wire N__45713;
    wire N__45710;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45622;
    wire N__45619;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45577;
    wire N__45576;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45566;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45556;
    wire N__45553;
    wire N__45546;
    wire N__45545;
    wire N__45544;
    wire N__45541;
    wire N__45538;
    wire N__45537;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45522;
    wire N__45521;
    wire N__45518;
    wire N__45515;
    wire N__45510;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45477;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45450;
    wire N__45441;
    wire N__45438;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45413;
    wire N__45410;
    wire N__45407;
    wire N__45404;
    wire N__45401;
    wire N__45398;
    wire N__45395;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45376;
    wire N__45373;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45365;
    wire N__45364;
    wire N__45363;
    wire N__45362;
    wire N__45359;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45330;
    wire N__45323;
    wire N__45322;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45306;
    wire N__45303;
    wire N__45290;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45254;
    wire N__45251;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45230;
    wire N__45227;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45215;
    wire N__45212;
    wire N__45209;
    wire N__45206;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45194;
    wire N__45193;
    wire N__45188;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45167;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45137;
    wire N__45134;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45090;
    wire N__45087;
    wire N__45086;
    wire N__45085;
    wire N__45084;
    wire N__45083;
    wire N__45082;
    wire N__45081;
    wire N__45080;
    wire N__45079;
    wire N__45078;
    wire N__45075;
    wire N__45074;
    wire N__45073;
    wire N__45072;
    wire N__45071;
    wire N__45070;
    wire N__45035;
    wire N__45032;
    wire N__45029;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45017;
    wire N__45016;
    wire N__45013;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44989;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44969;
    wire N__44966;
    wire N__44963;
    wire N__44960;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44927;
    wire N__44924;
    wire N__44921;
    wire N__44918;
    wire N__44915;
    wire N__44912;
    wire N__44909;
    wire N__44906;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44898;
    wire N__44897;
    wire N__44894;
    wire N__44891;
    wire N__44886;
    wire N__44879;
    wire N__44876;
    wire N__44873;
    wire N__44870;
    wire N__44869;
    wire N__44866;
    wire N__44863;
    wire N__44862;
    wire N__44861;
    wire N__44854;
    wire N__44851;
    wire N__44846;
    wire N__44845;
    wire N__44844;
    wire N__44841;
    wire N__44836;
    wire N__44833;
    wire N__44828;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44816;
    wire N__44815;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44789;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44765;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44753;
    wire N__44752;
    wire N__44751;
    wire N__44750;
    wire N__44749;
    wire N__44742;
    wire N__44737;
    wire N__44732;
    wire N__44729;
    wire N__44728;
    wire N__44725;
    wire N__44722;
    wire N__44719;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44696;
    wire N__44693;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44681;
    wire N__44678;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44666;
    wire N__44663;
    wire N__44660;
    wire N__44657;
    wire N__44654;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44643;
    wire N__44640;
    wire N__44637;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44608;
    wire N__44607;
    wire N__44604;
    wire N__44599;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44587;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44572;
    wire N__44567;
    wire N__44564;
    wire N__44563;
    wire N__44562;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44540;
    wire N__44537;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44492;
    wire N__44489;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44478;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44467;
    wire N__44464;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44441;
    wire N__44440;
    wire N__44439;
    wire N__44438;
    wire N__44435;
    wire N__44434;
    wire N__44431;
    wire N__44430;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44415;
    wire N__44410;
    wire N__44405;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44393;
    wire N__44390;
    wire N__44387;
    wire N__44382;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44308;
    wire N__44307;
    wire N__44304;
    wire N__44303;
    wire N__44302;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44281;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44233;
    wire N__44228;
    wire N__44223;
    wire N__44220;
    wire N__44215;
    wire N__44208;
    wire N__44201;
    wire N__44198;
    wire N__44197;
    wire N__44194;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44174;
    wire N__44173;
    wire N__44170;
    wire N__44169;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44128;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44120;
    wire N__44113;
    wire N__44110;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44078;
    wire N__44077;
    wire N__44074;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44059;
    wire N__44054;
    wire N__44051;
    wire N__44050;
    wire N__44047;
    wire N__44044;
    wire N__44041;
    wire N__44038;
    wire N__44035;
    wire N__44032;
    wire N__44029;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43979;
    wire N__43978;
    wire N__43975;
    wire N__43972;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43947;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43924;
    wire N__43921;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43909;
    wire N__43904;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43896;
    wire N__43891;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43879;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43820;
    wire N__43817;
    wire N__43816;
    wire N__43815;
    wire N__43814;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43806;
    wire N__43805;
    wire N__43804;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43780;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43762;
    wire N__43761;
    wire N__43760;
    wire N__43759;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43744;
    wire N__43741;
    wire N__43740;
    wire N__43737;
    wire N__43736;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43706;
    wire N__43703;
    wire N__43698;
    wire N__43693;
    wire N__43688;
    wire N__43685;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43668;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43583;
    wire N__43580;
    wire N__43579;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43547;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43535;
    wire N__43532;
    wire N__43529;
    wire N__43528;
    wire N__43525;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43507;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43489;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43469;
    wire N__43466;
    wire N__43463;
    wire N__43460;
    wire N__43459;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43439;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43424;
    wire N__43421;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43381;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43346;
    wire N__43343;
    wire N__43340;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43307;
    wire N__43304;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43283;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43253;
    wire N__43250;
    wire N__43247;
    wire N__43244;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43202;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43178;
    wire N__43175;
    wire N__43172;
    wire N__43169;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43161;
    wire N__43156;
    wire N__43155;
    wire N__43154;
    wire N__43153;
    wire N__43150;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43136;
    wire N__43133;
    wire N__43130;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43111;
    wire N__43108;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43089;
    wire N__43086;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43067;
    wire N__43064;
    wire N__43063;
    wire N__43060;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43022;
    wire N__43019;
    wire N__43016;
    wire N__43013;
    wire N__43010;
    wire N__43009;
    wire N__43006;
    wire N__43005;
    wire N__43004;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42987;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42972;
    wire N__42971;
    wire N__42970;
    wire N__42967;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42906;
    wire N__42903;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42856;
    wire N__42853;
    wire N__42852;
    wire N__42851;
    wire N__42848;
    wire N__42847;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42831;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42803;
    wire N__42800;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42784;
    wire N__42783;
    wire N__42782;
    wire N__42779;
    wire N__42778;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42741;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42724;
    wire N__42723;
    wire N__42722;
    wire N__42721;
    wire N__42718;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42659;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42626;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42610;
    wire N__42609;
    wire N__42608;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42604;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42582;
    wire N__42575;
    wire N__42574;
    wire N__42573;
    wire N__42568;
    wire N__42565;
    wire N__42560;
    wire N__42559;
    wire N__42558;
    wire N__42557;
    wire N__42550;
    wire N__42547;
    wire N__42542;
    wire N__42539;
    wire N__42538;
    wire N__42537;
    wire N__42536;
    wire N__42535;
    wire N__42526;
    wire N__42523;
    wire N__42518;
    wire N__42515;
    wire N__42512;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42500;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42488;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42473;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42461;
    wire N__42458;
    wire N__42457;
    wire N__42454;
    wire N__42451;
    wire N__42448;
    wire N__42443;
    wire N__42440;
    wire N__42439;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42421;
    wire N__42416;
    wire N__42415;
    wire N__42412;
    wire N__42409;
    wire N__42404;
    wire N__42403;
    wire N__42400;
    wire N__42397;
    wire N__42392;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42377;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42365;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42353;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42341;
    wire N__42338;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42220;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42190;
    wire N__42187;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42170;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42130;
    wire N__42127;
    wire N__42124;
    wire N__42121;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42088;
    wire N__42085;
    wire N__42080;
    wire N__42079;
    wire N__42076;
    wire N__42073;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42061;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42041;
    wire N__42040;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42017;
    wire N__42014;
    wire N__42013;
    wire N__42010;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41983;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41966;
    wire N__41963;
    wire N__41962;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41935;
    wire N__41930;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41918;
    wire N__41915;
    wire N__41912;
    wire N__41909;
    wire N__41906;
    wire N__41903;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41857;
    wire N__41848;
    wire N__41845;
    wire N__41840;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41832;
    wire N__41829;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41811;
    wire N__41806;
    wire N__41803;
    wire N__41798;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41786;
    wire N__41785;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41758;
    wire N__41755;
    wire N__41750;
    wire N__41749;
    wire N__41748;
    wire N__41747;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41734;
    wire N__41731;
    wire N__41730;
    wire N__41729;
    wire N__41728;
    wire N__41725;
    wire N__41722;
    wire N__41715;
    wire N__41710;
    wire N__41709;
    wire N__41708;
    wire N__41705;
    wire N__41696;
    wire N__41691;
    wire N__41684;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41669;
    wire N__41666;
    wire N__41663;
    wire N__41660;
    wire N__41657;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41637;
    wire N__41630;
    wire N__41627;
    wire N__41626;
    wire N__41625;
    wire N__41624;
    wire N__41623;
    wire N__41620;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41506;
    wire N__41501;
    wire N__41500;
    wire N__41499;
    wire N__41498;
    wire N__41495;
    wire N__41494;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41461;
    wire N__41456;
    wire N__41451;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41437;
    wire N__41434;
    wire N__41433;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41419;
    wire N__41418;
    wire N__41415;
    wire N__41412;
    wire N__41407;
    wire N__41402;
    wire N__41395;
    wire N__41390;
    wire N__41389;
    wire N__41388;
    wire N__41383;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41375;
    wire N__41372;
    wire N__41371;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41353;
    wire N__41348;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41323;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41308;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41294;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41284;
    wire N__41283;
    wire N__41280;
    wire N__41275;
    wire N__41270;
    wire N__41267;
    wire N__41264;
    wire N__41261;
    wire N__41258;
    wire N__41255;
    wire N__41252;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41234;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41216;
    wire N__41213;
    wire N__41210;
    wire N__41207;
    wire N__41204;
    wire N__41201;
    wire N__41198;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41167;
    wire N__41164;
    wire N__41163;
    wire N__41162;
    wire N__41159;
    wire N__41158;
    wire N__41157;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41108;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41077;
    wire N__41074;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41054;
    wire N__41053;
    wire N__41052;
    wire N__41051;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41042;
    wire N__41037;
    wire N__41036;
    wire N__41035;
    wire N__41032;
    wire N__41027;
    wire N__41024;
    wire N__41023;
    wire N__41022;
    wire N__41021;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40973;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40909;
    wire N__40906;
    wire N__40903;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40893;
    wire N__40890;
    wire N__40887;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40829;
    wire N__40826;
    wire N__40823;
    wire N__40820;
    wire N__40817;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40802;
    wire N__40801;
    wire N__40798;
    wire N__40797;
    wire N__40794;
    wire N__40793;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40758;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40727;
    wire N__40724;
    wire N__40721;
    wire N__40718;
    wire N__40715;
    wire N__40700;
    wire N__40697;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40673;
    wire N__40670;
    wire N__40667;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40654;
    wire N__40651;
    wire N__40650;
    wire N__40647;
    wire N__40646;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40624;
    wire N__40621;
    wire N__40620;
    wire N__40619;
    wire N__40614;
    wire N__40611;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40586;
    wire N__40583;
    wire N__40574;
    wire N__40571;
    wire N__40570;
    wire N__40569;
    wire N__40564;
    wire N__40563;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40551;
    wire N__40548;
    wire N__40543;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40526;
    wire N__40525;
    wire N__40524;
    wire N__40523;
    wire N__40522;
    wire N__40521;
    wire N__40520;
    wire N__40519;
    wire N__40516;
    wire N__40501;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40483;
    wire N__40480;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40457;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40449;
    wire N__40446;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40427;
    wire N__40424;
    wire N__40421;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40385;
    wire N__40382;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40340;
    wire N__40337;
    wire N__40334;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40307;
    wire N__40304;
    wire N__40301;
    wire N__40298;
    wire N__40295;
    wire N__40294;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40246;
    wire N__40245;
    wire N__40244;
    wire N__40241;
    wire N__40238;
    wire N__40235;
    wire N__40234;
    wire N__40233;
    wire N__40230;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40216;
    wire N__40215;
    wire N__40212;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40198;
    wire N__40197;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40175;
    wire N__40172;
    wire N__40171;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40163;
    wire N__40162;
    wire N__40161;
    wire N__40160;
    wire N__40157;
    wire N__40152;
    wire N__40143;
    wire N__40136;
    wire N__40135;
    wire N__40134;
    wire N__40133;
    wire N__40132;
    wire N__40131;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40119;
    wire N__40118;
    wire N__40117;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40111;
    wire N__40110;
    wire N__40109;
    wire N__40108;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40093;
    wire N__40090;
    wire N__40089;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40070;
    wire N__40067;
    wire N__40064;
    wire N__40061;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40053;
    wire N__40050;
    wire N__40049;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40035;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40018;
    wire N__40015;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39962;
    wire N__39957;
    wire N__39946;
    wire N__39939;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39904;
    wire N__39899;
    wire N__39896;
    wire N__39887;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39875;
    wire N__39872;
    wire N__39871;
    wire N__39868;
    wire N__39865;
    wire N__39860;
    wire N__39857;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39845;
    wire N__39842;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39827;
    wire N__39824;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39812;
    wire N__39809;
    wire N__39808;
    wire N__39805;
    wire N__39802;
    wire N__39797;
    wire N__39794;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39764;
    wire N__39763;
    wire N__39760;
    wire N__39757;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39746;
    wire N__39743;
    wire N__39740;
    wire N__39737;
    wire N__39734;
    wire N__39725;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39713;
    wire N__39710;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39698;
    wire N__39695;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39683;
    wire N__39680;
    wire N__39679;
    wire N__39676;
    wire N__39673;
    wire N__39670;
    wire N__39665;
    wire N__39662;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39650;
    wire N__39647;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39632;
    wire N__39629;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39614;
    wire N__39611;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39589;
    wire N__39586;
    wire N__39583;
    wire N__39578;
    wire N__39575;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39560;
    wire N__39557;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39545;
    wire N__39542;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39530;
    wire N__39527;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39515;
    wire N__39512;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39500;
    wire N__39497;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39467;
    wire N__39464;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39431;
    wire N__39428;
    wire N__39427;
    wire N__39424;
    wire N__39421;
    wire N__39418;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39322;
    wire N__39317;
    wire N__39314;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39289;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39275;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39253;
    wire N__39250;
    wire N__39247;
    wire N__39244;
    wire N__39239;
    wire N__39236;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39226;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39206;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39194;
    wire N__39191;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39157;
    wire N__39154;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39143;
    wire N__39142;
    wire N__39141;
    wire N__39140;
    wire N__39139;
    wire N__39138;
    wire N__39137;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39085;
    wire N__39076;
    wire N__39065;
    wire N__39062;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39035;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39016;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__38999;
    wire N__38996;
    wire N__38995;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38972;
    wire N__38969;
    wire N__38968;
    wire N__38967;
    wire N__38966;
    wire N__38965;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38957;
    wire N__38956;
    wire N__38955;
    wire N__38954;
    wire N__38951;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38936;
    wire N__38935;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38897;
    wire N__38894;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38876;
    wire N__38861;
    wire N__38858;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38843;
    wire N__38840;
    wire N__38839;
    wire N__38836;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38810;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38788;
    wire N__38785;
    wire N__38782;
    wire N__38779;
    wire N__38774;
    wire N__38771;
    wire N__38768;
    wire N__38767;
    wire N__38764;
    wire N__38761;
    wire N__38756;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38746;
    wire N__38741;
    wire N__38740;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38725;
    wire N__38722;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38618;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38594;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38579;
    wire N__38578;
    wire N__38575;
    wire N__38574;
    wire N__38573;
    wire N__38572;
    wire N__38571;
    wire N__38568;
    wire N__38567;
    wire N__38564;
    wire N__38563;
    wire N__38562;
    wire N__38561;
    wire N__38560;
    wire N__38559;
    wire N__38558;
    wire N__38557;
    wire N__38556;
    wire N__38555;
    wire N__38552;
    wire N__38549;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38524;
    wire N__38521;
    wire N__38516;
    wire N__38511;
    wire N__38502;
    wire N__38497;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38472;
    wire N__38471;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38456;
    wire N__38455;
    wire N__38454;
    wire N__38453;
    wire N__38452;
    wire N__38451;
    wire N__38450;
    wire N__38449;
    wire N__38448;
    wire N__38445;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38426;
    wire N__38423;
    wire N__38416;
    wire N__38399;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38352;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38336;
    wire N__38333;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38290;
    wire N__38287;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38263;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38237;
    wire N__38234;
    wire N__38231;
    wire N__38228;
    wire N__38225;
    wire N__38222;
    wire N__38219;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38186;
    wire N__38183;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38165;
    wire N__38162;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38148;
    wire N__38145;
    wire N__38142;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38126;
    wire N__38123;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38102;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38077;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38056;
    wire N__38051;
    wire N__38048;
    wire N__38045;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38014;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37971;
    wire N__37970;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37931;
    wire N__37930;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37912;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37865;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37799;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37786;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37742;
    wire N__37739;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37724;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37649;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37618;
    wire N__37615;
    wire N__37612;
    wire N__37609;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37516;
    wire N__37513;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37483;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37265;
    wire N__37264;
    wire N__37261;
    wire N__37258;
    wire N__37253;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37232;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37220;
    wire N__37217;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37202;
    wire N__37199;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37187;
    wire N__37186;
    wire N__37183;
    wire N__37180;
    wire N__37175;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37160;
    wire N__37157;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37124;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37112;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37102;
    wire N__37097;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37064;
    wire N__37061;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37049;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37034;
    wire N__37031;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36931;
    wire N__36926;
    wire N__36925;
    wire N__36922;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36824;
    wire N__36821;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36795;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36724;
    wire N__36721;
    wire N__36720;
    wire N__36719;
    wire N__36718;
    wire N__36717;
    wire N__36716;
    wire N__36715;
    wire N__36710;
    wire N__36709;
    wire N__36708;
    wire N__36707;
    wire N__36702;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36686;
    wire N__36685;
    wire N__36680;
    wire N__36677;
    wire N__36676;
    wire N__36675;
    wire N__36674;
    wire N__36669;
    wire N__36666;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36648;
    wire N__36635;
    wire N__36634;
    wire N__36631;
    wire N__36628;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36617;
    wire N__36614;
    wire N__36609;
    wire N__36606;
    wire N__36599;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36587;
    wire N__36586;
    wire N__36583;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36572;
    wire N__36569;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36548;
    wire N__36547;
    wire N__36544;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36482;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36433;
    wire N__36432;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36421;
    wire N__36420;
    wire N__36419;
    wire N__36418;
    wire N__36417;
    wire N__36416;
    wire N__36415;
    wire N__36414;
    wire N__36411;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36391;
    wire N__36382;
    wire N__36379;
    wire N__36370;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36345;
    wire N__36344;
    wire N__36339;
    wire N__36338;
    wire N__36337;
    wire N__36336;
    wire N__36335;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36316;
    wire N__36313;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36295;
    wire N__36292;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36275;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36254;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36221;
    wire N__36218;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36190;
    wire N__36185;
    wire N__36182;
    wire N__36181;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36166;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36121;
    wire N__36120;
    wire N__36119;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36111;
    wire N__36106;
    wire N__36103;
    wire N__36096;
    wire N__36093;
    wire N__36086;
    wire N__36085;
    wire N__36084;
    wire N__36083;
    wire N__36082;
    wire N__36081;
    wire N__36072;
    wire N__36067;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36039;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36013;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35869;
    wire N__35868;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35852;
    wire N__35851;
    wire N__35848;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35836;
    wire N__35831;
    wire N__35828;
    wire N__35817;
    wire N__35804;
    wire N__35803;
    wire N__35800;
    wire N__35799;
    wire N__35796;
    wire N__35793;
    wire N__35792;
    wire N__35791;
    wire N__35790;
    wire N__35789;
    wire N__35788;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35781;
    wire N__35776;
    wire N__35769;
    wire N__35766;
    wire N__35761;
    wire N__35754;
    wire N__35741;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35699;
    wire N__35698;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35674;
    wire N__35673;
    wire N__35670;
    wire N__35665;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35653;
    wire N__35650;
    wire N__35647;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35593;
    wire N__35590;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35573;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35567;
    wire N__35566;
    wire N__35563;
    wire N__35562;
    wire N__35559;
    wire N__35558;
    wire N__35555;
    wire N__35554;
    wire N__35551;
    wire N__35550;
    wire N__35547;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35510;
    wire N__35507;
    wire N__35506;
    wire N__35501;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35489;
    wire N__35484;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35468;
    wire N__35463;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35421;
    wire N__35420;
    wire N__35419;
    wire N__35418;
    wire N__35417;
    wire N__35416;
    wire N__35413;
    wire N__35412;
    wire N__35411;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35405;
    wire N__35404;
    wire N__35403;
    wire N__35402;
    wire N__35401;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35393;
    wire N__35392;
    wire N__35391;
    wire N__35390;
    wire N__35387;
    wire N__35382;
    wire N__35377;
    wire N__35376;
    wire N__35373;
    wire N__35372;
    wire N__35371;
    wire N__35370;
    wire N__35369;
    wire N__35368;
    wire N__35367;
    wire N__35366;
    wire N__35365;
    wire N__35364;
    wire N__35363;
    wire N__35362;
    wire N__35361;
    wire N__35358;
    wire N__35353;
    wire N__35348;
    wire N__35347;
    wire N__35346;
    wire N__35345;
    wire N__35344;
    wire N__35343;
    wire N__35342;
    wire N__35341;
    wire N__35332;
    wire N__35321;
    wire N__35320;
    wire N__35319;
    wire N__35316;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35298;
    wire N__35291;
    wire N__35288;
    wire N__35285;
    wire N__35270;
    wire N__35259;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35243;
    wire N__35234;
    wire N__35229;
    wire N__35224;
    wire N__35219;
    wire N__35218;
    wire N__35217;
    wire N__35216;
    wire N__35215;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35197;
    wire N__35192;
    wire N__35185;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35171;
    wire N__35170;
    wire N__35169;
    wire N__35168;
    wire N__35167;
    wire N__35166;
    wire N__35165;
    wire N__35158;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35140;
    wire N__35139;
    wire N__35134;
    wire N__35131;
    wire N__35130;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35096;
    wire N__35091;
    wire N__35088;
    wire N__35083;
    wire N__35076;
    wire N__35069;
    wire N__35048;
    wire N__35045;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35031;
    wire N__35030;
    wire N__35029;
    wire N__35026;
    wire N__35025;
    wire N__35024;
    wire N__35021;
    wire N__35020;
    wire N__35019;
    wire N__35018;
    wire N__35017;
    wire N__35014;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35000;
    wire N__34997;
    wire N__34988;
    wire N__34983;
    wire N__34980;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34960;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34942;
    wire N__34941;
    wire N__34940;
    wire N__34939;
    wire N__34938;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34926;
    wire N__34925;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34913;
    wire N__34910;
    wire N__34905;
    wire N__34896;
    wire N__34893;
    wire N__34888;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34834;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34796;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34762;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34750;
    wire N__34745;
    wire N__34742;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34720;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34702;
    wire N__34701;
    wire N__34698;
    wire N__34693;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34661;
    wire N__34660;
    wire N__34659;
    wire N__34658;
    wire N__34657;
    wire N__34656;
    wire N__34655;
    wire N__34654;
    wire N__34653;
    wire N__34652;
    wire N__34651;
    wire N__34650;
    wire N__34649;
    wire N__34648;
    wire N__34641;
    wire N__34638;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34622;
    wire N__34621;
    wire N__34618;
    wire N__34609;
    wire N__34606;
    wire N__34599;
    wire N__34596;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34588;
    wire N__34585;
    wire N__34584;
    wire N__34583;
    wire N__34580;
    wire N__34577;
    wire N__34574;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34558;
    wire N__34553;
    wire N__34548;
    wire N__34543;
    wire N__34538;
    wire N__34535;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34487;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34468;
    wire N__34465;
    wire N__34460;
    wire N__34457;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34440;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34424;
    wire N__34419;
    wire N__34416;
    wire N__34411;
    wire N__34410;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34388;
    wire N__34383;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34377;
    wire N__34370;
    wire N__34367;
    wire N__34362;
    wire N__34357;
    wire N__34350;
    wire N__34343;
    wire N__34340;
    wire N__34339;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34317;
    wire N__34314;
    wire N__34305;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34286;
    wire N__34283;
    wire N__34276;
    wire N__34271;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34251;
    wire N__34244;
    wire N__34241;
    wire N__34240;
    wire N__34235;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34217;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34193;
    wire N__34190;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34166;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34145;
    wire N__34142;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34052;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33986;
    wire N__33983;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33965;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33881;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33873;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33850;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33824;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33809;
    wire N__33808;
    wire N__33807;
    wire N__33806;
    wire N__33799;
    wire N__33796;
    wire N__33791;
    wire N__33790;
    wire N__33789;
    wire N__33784;
    wire N__33781;
    wire N__33776;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33768;
    wire N__33767;
    wire N__33766;
    wire N__33757;
    wire N__33754;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33673;
    wire N__33670;
    wire N__33669;
    wire N__33668;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33654;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33631;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33589;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33560;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33532;
    wire N__33529;
    wire N__33524;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33520;
    wire N__33519;
    wire N__33518;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33494;
    wire N__33493;
    wire N__33492;
    wire N__33491;
    wire N__33488;
    wire N__33481;
    wire N__33478;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33474;
    wire N__33473;
    wire N__33472;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33451;
    wire N__33448;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33421;
    wire N__33412;
    wire N__33409;
    wire N__33400;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33373;
    wire N__33372;
    wire N__33371;
    wire N__33368;
    wire N__33367;
    wire N__33366;
    wire N__33365;
    wire N__33364;
    wire N__33363;
    wire N__33362;
    wire N__33359;
    wire N__33358;
    wire N__33355;
    wire N__33354;
    wire N__33351;
    wire N__33350;
    wire N__33349;
    wire N__33348;
    wire N__33347;
    wire N__33346;
    wire N__33345;
    wire N__33344;
    wire N__33341;
    wire N__33340;
    wire N__33339;
    wire N__33338;
    wire N__33337;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33311;
    wire N__33302;
    wire N__33301;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33286;
    wire N__33285;
    wire N__33284;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33267;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33249;
    wire N__33246;
    wire N__33241;
    wire N__33240;
    wire N__33239;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33234;
    wire N__33217;
    wire N__33214;
    wire N__33207;
    wire N__33202;
    wire N__33191;
    wire N__33180;
    wire N__33175;
    wire N__33172;
    wire N__33167;
    wire N__33164;
    wire N__33157;
    wire N__33146;
    wire N__33141;
    wire N__33128;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33124;
    wire N__33123;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33119;
    wire N__33118;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33114;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33110;
    wire N__33109;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33101;
    wire N__33100;
    wire N__33099;
    wire N__33098;
    wire N__33097;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33086;
    wire N__33085;
    wire N__33084;
    wire N__33083;
    wire N__33082;
    wire N__33081;
    wire N__33076;
    wire N__33063;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33043;
    wire N__33042;
    wire N__33035;
    wire N__33028;
    wire N__33023;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33012;
    wire N__33011;
    wire N__33008;
    wire N__32997;
    wire N__32994;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32984;
    wire N__32983;
    wire N__32974;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32956;
    wire N__32951;
    wire N__32942;
    wire N__32929;
    wire N__32924;
    wire N__32909;
    wire N__32906;
    wire N__32905;
    wire N__32904;
    wire N__32903;
    wire N__32902;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32887;
    wire N__32884;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32870;
    wire N__32869;
    wire N__32868;
    wire N__32867;
    wire N__32866;
    wire N__32861;
    wire N__32860;
    wire N__32859;
    wire N__32858;
    wire N__32857;
    wire N__32852;
    wire N__32847;
    wire N__32846;
    wire N__32845;
    wire N__32842;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32799;
    wire N__32794;
    wire N__32785;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32734;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32693;
    wire N__32690;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32678;
    wire N__32677;
    wire N__32674;
    wire N__32671;
    wire N__32666;
    wire N__32665;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32651;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32639;
    wire N__32636;
    wire N__32633;
    wire N__32630;
    wire N__32627;
    wire N__32624;
    wire N__32621;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32609;
    wire N__32608;
    wire N__32605;
    wire N__32602;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32584;
    wire N__32579;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32567;
    wire N__32564;
    wire N__32561;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32549;
    wire N__32546;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32533;
    wire N__32530;
    wire N__32527;
    wire N__32524;
    wire N__32519;
    wire N__32516;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32468;
    wire N__32465;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32450;
    wire N__32447;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32380;
    wire N__32375;
    wire N__32372;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32338;
    wire N__32337;
    wire N__32334;
    wire N__32329;
    wire N__32324;
    wire N__32321;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32255;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32231;
    wire N__32228;
    wire N__32227;
    wire N__32226;
    wire N__32221;
    wire N__32218;
    wire N__32217;
    wire N__32214;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32181;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32149;
    wire N__32146;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32129;
    wire N__32126;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32105;
    wire N__32102;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32091;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32065;
    wire N__32054;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32046;
    wire N__32045;
    wire N__32044;
    wire N__32041;
    wire N__32038;
    wire N__32033;
    wire N__32032;
    wire N__32029;
    wire N__32028;
    wire N__32027;
    wire N__32020;
    wire N__32013;
    wire N__32010;
    wire N__32003;
    wire N__32002;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31990;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31966;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31936;
    wire N__31933;
    wire N__31928;
    wire N__31925;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31913;
    wire N__31910;
    wire N__31907;
    wire N__31904;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31889;
    wire N__31886;
    wire N__31883;
    wire N__31882;
    wire N__31881;
    wire N__31880;
    wire N__31877;
    wire N__31874;
    wire N__31869;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31768;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31745;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31706;
    wire N__31703;
    wire N__31702;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31684;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31619;
    wire N__31616;
    wire N__31613;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31457;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31394;
    wire N__31391;
    wire N__31390;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31373;
    wire N__31370;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31301;
    wire N__31300;
    wire N__31299;
    wire N__31296;
    wire N__31291;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31276;
    wire N__31275;
    wire N__31272;
    wire N__31267;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31249;
    wire N__31246;
    wire N__31245;
    wire N__31244;
    wire N__31241;
    wire N__31234;
    wire N__31229;
    wire N__31228;
    wire N__31227;
    wire N__31226;
    wire N__31223;
    wire N__31216;
    wire N__31211;
    wire N__31208;
    wire N__31207;
    wire N__31206;
    wire N__31203;
    wire N__31198;
    wire N__31193;
    wire N__31190;
    wire N__31189;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31174;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31118;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31067;
    wire N__31066;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31051;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31034;
    wire N__31031;
    wire N__31030;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31013;
    wire N__31010;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30995;
    wire N__30994;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30979;
    wire N__30974;
    wire N__30971;
    wire N__30968;
    wire N__30967;
    wire N__30966;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30947;
    wire N__30946;
    wire N__30943;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30923;
    wire N__30920;
    wire N__30917;
    wire N__30914;
    wire N__30911;
    wire N__30910;
    wire N__30909;
    wire N__30904;
    wire N__30901;
    wire N__30896;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30881;
    wire N__30878;
    wire N__30877;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30859;
    wire N__30854;
    wire N__30851;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30833;
    wire N__30830;
    wire N__30827;
    wire N__30824;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30813;
    wire N__30808;
    wire N__30805;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30584;
    wire N__30581;
    wire N__30580;
    wire N__30577;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30536;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30511;
    wire N__30510;
    wire N__30507;
    wire N__30502;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30460;
    wire N__30459;
    wire N__30456;
    wire N__30451;
    wire N__30446;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30434;
    wire N__30431;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30398;
    wire N__30397;
    wire N__30396;
    wire N__30393;
    wire N__30388;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30280;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30175;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30061;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29961;
    wire N__29958;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29899;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29786;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29524;
    wire N__29519;
    wire N__29516;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29468;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29434;
    wire N__29429;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29399;
    wire N__29398;
    wire N__29395;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29369;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29345;
    wire N__29342;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29311;
    wire N__29310;
    wire N__29307;
    wire N__29302;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29261;
    wire N__29260;
    wire N__29257;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29245;
    wire N__29240;
    wire N__29239;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29216;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29204;
    wire N__29201;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29177;
    wire N__29174;
    wire N__29173;
    wire N__29172;
    wire N__29171;
    wire N__29170;
    wire N__29169;
    wire N__29168;
    wire N__29167;
    wire N__29166;
    wire N__29165;
    wire N__29164;
    wire N__29163;
    wire N__29162;
    wire N__29161;
    wire N__29160;
    wire N__29159;
    wire N__29154;
    wire N__29151;
    wire N__29150;
    wire N__29147;
    wire N__29132;
    wire N__29131;
    wire N__29128;
    wire N__29127;
    wire N__29126;
    wire N__29125;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29111;
    wire N__29110;
    wire N__29107;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29093;
    wire N__29090;
    wire N__29073;
    wire N__29068;
    wire N__29065;
    wire N__29058;
    wire N__29045;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29033;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29006;
    wire N__29005;
    wire N__29002;
    wire N__29001;
    wire N__29000;
    wire N__28997;
    wire N__28996;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28979;
    wire N__28974;
    wire N__28969;
    wire N__28964;
    wire N__28961;
    wire N__28958;
    wire N__28955;
    wire N__28952;
    wire N__28947;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28906;
    wire N__28905;
    wire N__28902;
    wire N__28897;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28874;
    wire N__28871;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28859;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28847;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28835;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28824;
    wire N__28821;
    wire N__28818;
    wire N__28815;
    wire N__28810;
    wire N__28807;
    wire N__28802;
    wire N__28799;
    wire N__28796;
    wire N__28795;
    wire N__28794;
    wire N__28791;
    wire N__28786;
    wire N__28781;
    wire N__28780;
    wire N__28777;
    wire N__28776;
    wire N__28773;
    wire N__28766;
    wire N__28763;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28697;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28670;
    wire N__28669;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28610;
    wire N__28607;
    wire N__28606;
    wire N__28605;
    wire N__28602;
    wire N__28597;
    wire N__28592;
    wire N__28589;
    wire N__28586;
    wire N__28585;
    wire N__28582;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28537;
    wire N__28532;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28514;
    wire N__28511;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28465;
    wire N__28464;
    wire N__28461;
    wire N__28456;
    wire N__28451;
    wire N__28448;
    wire N__28445;
    wire N__28442;
    wire N__28441;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28414;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28376;
    wire N__28373;
    wire N__28372;
    wire N__28369;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28357;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28339;
    wire N__28336;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28288;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28148;
    wire N__28145;
    wire N__28144;
    wire N__28143;
    wire N__28140;
    wire N__28135;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28117;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28102;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28060;
    wire N__28057;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28034;
    wire N__28031;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27985;
    wire N__27984;
    wire N__27981;
    wire N__27976;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27912;
    wire N__27907;
    wire N__27904;
    wire N__27899;
    wire N__27898;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27883;
    wire N__27880;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27863;
    wire N__27862;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27845;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27716;
    wire N__27713;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27674;
    wire N__27673;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27626;
    wire N__27623;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27572;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27538;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27506;
    wire N__27505;
    wire N__27502;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27484;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27473;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27455;
    wire N__27452;
    wire N__27451;
    wire N__27448;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27403;
    wire N__27400;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27272;
    wire N__27271;
    wire N__27270;
    wire N__27265;
    wire N__27262;
    wire N__27257;
    wire N__27256;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27173;
    wire N__27172;
    wire N__27171;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27117;
    wire N__27114;
    wire N__27107;
    wire N__27106;
    wire N__27105;
    wire N__27104;
    wire N__27101;
    wire N__27100;
    wire N__27099;
    wire N__27096;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27055;
    wire N__27052;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26971;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26948;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26846;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26825;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26807;
    wire N__26804;
    wire N__26803;
    wire N__26802;
    wire N__26799;
    wire N__26794;
    wire N__26791;
    wire N__26786;
    wire N__26783;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26771;
    wire N__26768;
    wire N__26767;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26752;
    wire N__26749;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26726;
    wire N__26723;
    wire N__26722;
    wire N__26721;
    wire N__26718;
    wire N__26713;
    wire N__26710;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26684;
    wire N__26681;
    wire N__26680;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26642;
    wire N__26639;
    wire N__26638;
    wire N__26637;
    wire N__26634;
    wire N__26629;
    wire N__26626;
    wire N__26621;
    wire N__26618;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26569;
    wire N__26568;
    wire N__26565;
    wire N__26560;
    wire N__26557;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26524;
    wire N__26521;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26491;
    wire N__26488;
    wire N__26487;
    wire N__26484;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26455;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26392;
    wire N__26391;
    wire N__26388;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26372;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26364;
    wire N__26361;
    wire N__26356;
    wire N__26353;
    wire N__26348;
    wire N__26345;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26328;
    wire N__26323;
    wire N__26320;
    wire N__26315;
    wire N__26312;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26299;
    wire N__26294;
    wire N__26291;
    wire N__26290;
    wire N__26289;
    wire N__26288;
    wire N__26285;
    wire N__26284;
    wire N__26281;
    wire N__26280;
    wire N__26279;
    wire N__26278;
    wire N__26277;
    wire N__26276;
    wire N__26275;
    wire N__26274;
    wire N__26273;
    wire N__26262;
    wire N__26259;
    wire N__26256;
    wire N__26255;
    wire N__26254;
    wire N__26251;
    wire N__26250;
    wire N__26247;
    wire N__26246;
    wire N__26243;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26237;
    wire N__26236;
    wire N__26233;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26215;
    wire N__26202;
    wire N__26189;
    wire N__26180;
    wire N__26179;
    wire N__26176;
    wire N__26175;
    wire N__26172;
    wire N__26167;
    wire N__26164;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26152;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26122;
    wire N__26121;
    wire N__26118;
    wire N__26113;
    wire N__26110;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26095;
    wire N__26092;
    wire N__26091;
    wire N__26088;
    wire N__26083;
    wire N__26080;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26065;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26035;
    wire N__26032;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26002;
    wire N__26001;
    wire N__25998;
    wire N__25993;
    wire N__25990;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25945;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25927;
    wire N__25922;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25901;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25889;
    wire N__25886;
    wire N__25885;
    wire N__25882;
    wire N__25879;
    wire N__25878;
    wire N__25875;
    wire N__25870;
    wire N__25865;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25846;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25798;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25781;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25744;
    wire N__25741;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25609;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25592;
    wire N__25591;
    wire N__25588;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25550;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25439;
    wire N__25436;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25340;
    wire N__25333;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25280;
    wire N__25277;
    wire N__25276;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25261;
    wire N__25256;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25229;
    wire N__25228;
    wire N__25225;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25205;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25197;
    wire N__25196;
    wire N__25191;
    wire N__25188;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25163;
    wire N__25160;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25121;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25103;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25085;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25048;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25040;
    wire N__25039;
    wire N__25038;
    wire N__25035;
    wire N__25034;
    wire N__25033;
    wire N__25032;
    wire N__25031;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25017;
    wire N__25016;
    wire N__25015;
    wire N__25014;
    wire N__25013;
    wire N__25012;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24989;
    wire N__24984;
    wire N__24981;
    wire N__24976;
    wire N__24969;
    wire N__24960;
    wire N__24953;
    wire N__24944;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24893;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24871;
    wire N__24866;
    wire N__24865;
    wire N__24864;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24850;
    wire N__24849;
    wire N__24848;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24844;
    wire N__24843;
    wire N__24842;
    wire N__24841;
    wire N__24840;
    wire N__24839;
    wire N__24826;
    wire N__24823;
    wire N__24814;
    wire N__24809;
    wire N__24808;
    wire N__24807;
    wire N__24806;
    wire N__24805;
    wire N__24804;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24793;
    wire N__24786;
    wire N__24781;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24769;
    wire N__24766;
    wire N__24765;
    wire N__24756;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24731;
    wire N__24724;
    wire N__24721;
    wire N__24716;
    wire N__24711;
    wire N__24708;
    wire N__24683;
    wire N__24682;
    wire N__24681;
    wire N__24680;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24676;
    wire N__24675;
    wire N__24674;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24666;
    wire N__24665;
    wire N__24664;
    wire N__24661;
    wire N__24660;
    wire N__24659;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24648;
    wire N__24645;
    wire N__24644;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24636;
    wire N__24635;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24621;
    wire N__24616;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24592;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24584;
    wire N__24579;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24561;
    wire N__24554;
    wire N__24551;
    wire N__24546;
    wire N__24543;
    wire N__24538;
    wire N__24529;
    wire N__24518;
    wire N__24515;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24473;
    wire N__24472;
    wire N__24471;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24467;
    wire N__24466;
    wire N__24463;
    wire N__24456;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24448;
    wire N__24447;
    wire N__24446;
    wire N__24445;
    wire N__24444;
    wire N__24443;
    wire N__24442;
    wire N__24441;
    wire N__24440;
    wire N__24439;
    wire N__24438;
    wire N__24437;
    wire N__24436;
    wire N__24435;
    wire N__24434;
    wire N__24433;
    wire N__24432;
    wire N__24431;
    wire N__24428;
    wire N__24427;
    wire N__24426;
    wire N__24425;
    wire N__24424;
    wire N__24423;
    wire N__24422;
    wire N__24421;
    wire N__24420;
    wire N__24419;
    wire N__24418;
    wire N__24417;
    wire N__24414;
    wire N__24413;
    wire N__24412;
    wire N__24411;
    wire N__24410;
    wire N__24409;
    wire N__24406;
    wire N__24401;
    wire N__24394;
    wire N__24383;
    wire N__24372;
    wire N__24371;
    wire N__24370;
    wire N__24369;
    wire N__24362;
    wire N__24351;
    wire N__24334;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24316;
    wire N__24311;
    wire N__24302;
    wire N__24299;
    wire N__24292;
    wire N__24287;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24241;
    wire N__24236;
    wire N__24235;
    wire N__24234;
    wire N__24233;
    wire N__24230;
    wire N__24229;
    wire N__24228;
    wire N__24227;
    wire N__24224;
    wire N__24223;
    wire N__24222;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24218;
    wire N__24213;
    wire N__24208;
    wire N__24203;
    wire N__24202;
    wire N__24201;
    wire N__24194;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24156;
    wire N__24143;
    wire N__24142;
    wire N__24141;
    wire N__24140;
    wire N__24139;
    wire N__24128;
    wire N__24127;
    wire N__24126;
    wire N__24125;
    wire N__24122;
    wire N__24115;
    wire N__24110;
    wire N__24109;
    wire N__24108;
    wire N__24107;
    wire N__24106;
    wire N__24105;
    wire N__24104;
    wire N__24103;
    wire N__24102;
    wire N__24091;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24065;
    wire N__24064;
    wire N__24063;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24051;
    wire N__24048;
    wire N__24047;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24026;
    wire N__24023;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23977;
    wire N__23976;
    wire N__23973;
    wire N__23968;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23939;
    wire N__23936;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23926;
    wire N__23925;
    wire N__23922;
    wire N__23917;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23858;
    wire N__23855;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23840;
    wire N__23837;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23801;
    wire N__23798;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23767;
    wire N__23766;
    wire N__23763;
    wire N__23758;
    wire N__23755;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23731;
    wire N__23728;
    wire N__23727;
    wire N__23720;
    wire N__23717;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23709;
    wire N__23706;
    wire N__23701;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23687;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23675;
    wire N__23672;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23654;
    wire N__23651;
    wire N__23650;
    wire N__23647;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23623;
    wire N__23622;
    wire N__23619;
    wire N__23614;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23512;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23497;
    wire N__23496;
    wire N__23495;
    wire N__23494;
    wire N__23491;
    wire N__23490;
    wire N__23489;
    wire N__23488;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23465;
    wire N__23460;
    wire N__23451;
    wire N__23444;
    wire N__23441;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23421;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23377;
    wire N__23372;
    wire N__23367;
    wire N__23360;
    wire N__23359;
    wire N__23358;
    wire N__23357;
    wire N__23354;
    wire N__23353;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23342;
    wire N__23341;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23334;
    wire N__23333;
    wire N__23332;
    wire N__23331;
    wire N__23328;
    wire N__23327;
    wire N__23326;
    wire N__23325;
    wire N__23324;
    wire N__23323;
    wire N__23320;
    wire N__23319;
    wire N__23318;
    wire N__23317;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23305;
    wire N__23302;
    wire N__23287;
    wire N__23278;
    wire N__23275;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23240;
    wire N__23229;
    wire N__23228;
    wire N__23217;
    wire N__23214;
    wire N__23207;
    wire N__23204;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23170;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23145;
    wire N__23144;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23126;
    wire N__23125;
    wire N__23122;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23100;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23011;
    wire N__23008;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22954;
    wire N__22951;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22931;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22906;
    wire N__22905;
    wire N__22902;
    wire N__22897;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22849;
    wire N__22848;
    wire N__22845;
    wire N__22840;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22819;
    wire N__22818;
    wire N__22815;
    wire N__22810;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22783;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22744;
    wire N__22743;
    wire N__22740;
    wire N__22735;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22684;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22633;
    wire N__22632;
    wire N__22629;
    wire N__22624;
    wire N__22619;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22582;
    wire N__22581;
    wire N__22580;
    wire N__22577;
    wire N__22576;
    wire N__22575;
    wire N__22574;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22543;
    wire N__22540;
    wire N__22533;
    wire N__22532;
    wire N__22529;
    wire N__22524;
    wire N__22521;
    wire N__22516;
    wire N__22513;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22493;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22469;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22440;
    wire N__22437;
    wire N__22430;
    wire N__22427;
    wire N__22426;
    wire N__22425;
    wire N__22422;
    wire N__22417;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22390;
    wire N__22389;
    wire N__22388;
    wire N__22387;
    wire N__22384;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22264;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22249;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22168;
    wire N__22167;
    wire N__22166;
    wire N__22165;
    wire N__22164;
    wire N__22163;
    wire N__22162;
    wire N__22161;
    wire N__22160;
    wire N__22159;
    wire N__22158;
    wire N__22157;
    wire N__22156;
    wire N__22155;
    wire N__22154;
    wire N__22147;
    wire N__22140;
    wire N__22133;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22098;
    wire N__22095;
    wire N__22088;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22076;
    wire N__22073;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22043;
    wire N__22040;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21973;
    wire N__21970;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21928;
    wire N__21923;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21886;
    wire N__21885;
    wire N__21882;
    wire N__21877;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21862;
    wire N__21861;
    wire N__21858;
    wire N__21853;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21815;
    wire N__21814;
    wire N__21811;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21736;
    wire N__21735;
    wire N__21730;
    wire N__21727;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21704;
    wire N__21701;
    wire N__21700;
    wire N__21699;
    wire N__21696;
    wire N__21691;
    wire N__21686;
    wire N__21685;
    wire N__21682;
    wire N__21681;
    wire N__21678;
    wire N__21671;
    wire N__21668;
    wire N__21667;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21655;
    wire N__21652;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21621;
    wire N__21618;
    wire N__21613;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21586;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21568;
    wire N__21563;
    wire N__21562;
    wire N__21561;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21546;
    wire N__21545;
    wire N__21542;
    wire N__21529;
    wire N__21526;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21513;
    wire N__21510;
    wire N__21505;
    wire N__21498;
    wire N__21493;
    wire N__21490;
    wire N__21479;
    wire N__21478;
    wire N__21477;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21463;
    wire N__21462;
    wire N__21459;
    wire N__21454;
    wire N__21449;
    wire N__21448;
    wire N__21445;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21433;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21334;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21287;
    wire N__21284;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21272;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21260;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21238;
    wire N__21235;
    wire N__21232;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21192;
    wire N__21189;
    wire N__21182;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21170;
    wire N__21167;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21115;
    wire N__21112;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21100;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21071;
    wire N__21070;
    wire N__21069;
    wire N__21068;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21053;
    wire N__21050;
    wire N__21041;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21029;
    wire N__21028;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21020;
    wire N__21017;
    wire N__21016;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20973;
    wire N__20972;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20960;
    wire N__20957;
    wire N__20948;
    wire N__20947;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20893;
    wire N__20888;
    wire N__20885;
    wire N__20884;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20855;
    wire N__20852;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20840;
    wire N__20837;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20759;
    wire N__20756;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20710;
    wire N__20707;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20687;
    wire N__20684;
    wire N__20683;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20671;
    wire N__20670;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20658;
    wire N__20657;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20594;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20582;
    wire N__20579;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20564;
    wire N__20561;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20549;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20523;
    wire N__20520;
    wire N__20515;
    wire N__20510;
    wire N__20507;
    wire N__20506;
    wire N__20505;
    wire N__20502;
    wire N__20497;
    wire N__20492;
    wire N__20491;
    wire N__20490;
    wire N__20487;
    wire N__20486;
    wire N__20483;
    wire N__20482;
    wire N__20471;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20447;
    wire N__20444;
    wire N__20443;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20419;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20381;
    wire N__20378;
    wire N__20377;
    wire N__20372;
    wire N__20369;
    wire N__20368;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20314;
    wire N__20311;
    wire N__20310;
    wire N__20309;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20294;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20262;
    wire N__20259;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20188;
    wire N__20183;
    wire N__20180;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20170;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20143;
    wire N__20142;
    wire N__20139;
    wire N__20134;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20124;
    wire N__20119;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20029;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19994;
    wire N__19993;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19975;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19910;
    wire N__19909;
    wire N__19908;
    wire N__19901;
    wire N__19900;
    wire N__19899;
    wire N__19896;
    wire N__19891;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19853;
    wire N__19852;
    wire N__19849;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19784;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19769;
    wire N__19766;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19751;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19736;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19721;
    wire N__19720;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19706;
    wire N__19703;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19688;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19627;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19610;
    wire N__19609;
    wire N__19608;
    wire N__19605;
    wire N__19600;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19576;
    wire N__19573;
    wire N__19568;
    wire N__19567;
    wire N__19566;
    wire N__19563;
    wire N__19562;
    wire N__19559;
    wire N__19552;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19421;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19409;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19366;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19343;
    wire N__19342;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19330;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19274;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19259;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19247;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19235;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19220;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire ICE_GPMO_2;
    wire VCCG0;
    wire INViac_raw_buf_vac_raw_buf_merged11WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged3WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged10WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged8WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged4WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged9WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged5WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged0WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged6WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged1WCLKN_net;
    wire ICE_SYSCLK;
    wire INViac_raw_buf_vac_raw_buf_merged7WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged2WCLKN_net;
    wire bfn_2_7_0_;
    wire \ADC_VAC.n19408 ;
    wire \ADC_VAC.n19409 ;
    wire \ADC_VAC.n19410 ;
    wire \ADC_VAC.n19411 ;
    wire \ADC_VAC.n19412 ;
    wire \ADC_VAC.n19413 ;
    wire \ADC_VAC.n19414 ;
    wire \ADC_VAC.bit_cnt_0 ;
    wire \ADC_VAC.bit_cnt_6 ;
    wire \ADC_VAC.bit_cnt_4 ;
    wire \ADC_VAC.bit_cnt_3 ;
    wire \ADC_VAC.bit_cnt_5 ;
    wire \ADC_VAC.bit_cnt_2 ;
    wire \ADC_VAC.bit_cnt_7 ;
    wire \ADC_VAC.bit_cnt_1 ;
    wire \ADC_VAC.n21054_cascade_ ;
    wire \ADC_VAC.n16 ;
    wire VAC_MISO;
    wire cmd_rdadctmp_0;
    wire cmd_rdadctmp_1;
    wire cmd_rdadctmp_2;
    wire cmd_rdadctmp_3;
    wire \ADC_VAC.n14822 ;
    wire \ADC_VAC.n20715_cascade_ ;
    wire \ADC_VAC.n21053 ;
    wire \ADC_VAC.n20716 ;
    wire \ADC_VAC.n17_cascade_ ;
    wire \ADC_VAC.n12 ;
    wire \ADC_VAC.n12489 ;
    wire VAC_SCLK;
    wire n14_adj_1606_cascade_;
    wire VAC_CS;
    wire n20615;
    wire VAC_DRDY;
    wire n20615_cascade_;
    wire bit_cnt_2;
    wire bit_cnt_1;
    wire \CLK_DDS.n16766 ;
    wire bfn_5_5_0_;
    wire \ADC_VDC.n19457 ;
    wire \ADC_VDC.n19458 ;
    wire \ADC_VDC.n19459 ;
    wire \ADC_VDC.n19460 ;
    wire \ADC_VDC.n19461 ;
    wire \ADC_VDC.n19462 ;
    wire \ADC_VDC.n19463 ;
    wire \ADC_VDC.n19464 ;
    wire bfn_5_6_0_;
    wire \ADC_VDC.n19465 ;
    wire \ADC_VDC.n19466 ;
    wire \ADC_VDC.n19467 ;
    wire \ADC_VDC.avg_cnt_4 ;
    wire \ADC_VDC.avg_cnt_7 ;
    wire \ADC_VDC.avg_cnt_3 ;
    wire \ADC_VDC.avg_cnt_5 ;
    wire \ADC_VDC.avg_cnt_9 ;
    wire \ADC_VDC.avg_cnt_0 ;
    wire \ADC_VDC.avg_cnt_8 ;
    wire \ADC_VDC.avg_cnt_10 ;
    wire \ADC_VDC.n20 ;
    wire \ADC_VDC.n19_adj_1412_cascade_ ;
    wire \ADC_VDC.n18479_cascade_ ;
    wire DDS_CS1;
    wire RTD_SDO;
    wire \CLK_DDS.tmp_buf_0 ;
    wire bit_cnt_3;
    wire bit_cnt_0_adj_1456;
    wire \ADC_IAC.n17_cascade_ ;
    wire DDS_SCK1;
    wire cmd_rdadctmp_6_adj_1444;
    wire \ADC_IAC.n12 ;
    wire n20612_cascade_;
    wire \ADC_IAC.n20713 ;
    wire \ADC_IAC.n20783_cascade_ ;
    wire \ADC_IAC.n20795_cascade_ ;
    wire \ADC_IAC.n21068_cascade_ ;
    wire \ADC_IAC.n20714 ;
    wire IAC_MISO;
    wire cmd_rdadctmp_0_adj_1450;
    wire IAC_SCLK;
    wire cmd_rdadctmp_28;
    wire bfn_6_6_0_;
    wire \ADC_VDC.n19531 ;
    wire \ADC_VDC.n19532 ;
    wire \ADC_VDC.n19533 ;
    wire \ADC_VDC.n19534 ;
    wire \ADC_VDC.n19535 ;
    wire \ADC_VDC.n19536 ;
    wire \ADC_VDC.n19537 ;
    wire \ADC_VDC.bit_cnt_5 ;
    wire \ADC_VDC.n20534_cascade_ ;
    wire \ADC_VDC.n10 ;
    wire \ADC_VDC.bit_cnt_7 ;
    wire \ADC_VDC.bit_cnt_6 ;
    wire \ADC_VDC.n21082 ;
    wire \ADC_VDC.n21079 ;
    wire \ADC_VDC.n21977_cascade_ ;
    wire \ADC_VDC.n18482 ;
    wire \ADC_VDC.bit_cnt_2 ;
    wire \ADC_VDC.n6 ;
    wire \ADC_VDC.n10552_cascade_ ;
    wire \ADC_VDC.n21974 ;
    wire \ADC_VDC.bit_cnt_3 ;
    wire \ADC_VDC.n20562 ;
    wire \ADC_VDC.n21224_cascade_ ;
    wire \ADC_VDC.n20748 ;
    wire \ADC_VDC.n31_cascade_ ;
    wire \ADC_VDC.n20555 ;
    wire read_buf_12;
    wire adress_3;
    wire adress_2;
    wire adress_4;
    wire adress_5;
    wire RTD_SDI;
    wire \RTD.n21309_cascade_ ;
    wire \RTD.n12 ;
    wire \RTD.n19_cascade_ ;
    wire read_buf_9;
    wire adress_1;
    wire read_buf_1;
    wire read_buf_13;
    wire read_buf_8;
    wire n20754;
    wire cmd_rdadctmp_5_adj_1445;
    wire cmd_rdadctmp_4_adj_1446;
    wire cmd_rdadctmp_3_adj_1447;
    wire IAC_DRDY;
    wire n20612;
    wire n14_adj_1604_cascade_;
    wire IAC_CS;
    wire \ADC_IAC.bit_cnt_0 ;
    wire bfn_6_15_0_;
    wire \ADC_IAC.bit_cnt_1 ;
    wire \ADC_IAC.n19415 ;
    wire \ADC_IAC.bit_cnt_2 ;
    wire \ADC_IAC.n19416 ;
    wire \ADC_IAC.bit_cnt_3 ;
    wire \ADC_IAC.n19417 ;
    wire \ADC_IAC.bit_cnt_4 ;
    wire \ADC_IAC.n19418 ;
    wire \ADC_IAC.bit_cnt_5 ;
    wire \ADC_IAC.n19419 ;
    wire \ADC_IAC.bit_cnt_6 ;
    wire \ADC_IAC.n19420 ;
    wire \ADC_IAC.n19421 ;
    wire \ADC_IAC.bit_cnt_7 ;
    wire \ADC_IAC.n12586 ;
    wire \ADC_IAC.n14860 ;
    wire cmd_rdadctmp_1_adj_1449;
    wire cmd_rdadctmp_2_adj_1448;
    wire DDS_MCLK1;
    wire cmd_rdadctmp_28_adj_1422;
    wire \ADC_VDC.n19_adj_1413_cascade_ ;
    wire \ADC_VDC.n17 ;
    wire \ADC_VDC.n4 ;
    wire \ADC_VDC.n10132_cascade_ ;
    wire \ADC_VDC.n7_adj_1411 ;
    wire \ADC_VDC.n20750 ;
    wire \ADC_VDC.n12 ;
    wire \ADC_VDC.n20750_cascade_ ;
    wire \ADC_VDC.n11692_cascade_ ;
    wire VDC_SCLK;
    wire \ADC_VDC.bit_cnt_1 ;
    wire \ADC_VDC.n20534 ;
    wire \ADC_VDC.bit_cnt_4 ;
    wire \ADC_VDC.n6_adj_1410 ;
    wire \ADC_VDC.n11281_cascade_ ;
    wire \ADC_VDC.bit_cnt_0 ;
    wire \ADC_VDC.n15 ;
    wire \ADC_VDC.n15_cascade_ ;
    wire \ADC_VDC.n20746_cascade_ ;
    wire \ADC_VDC.n72 ;
    wire \ADC_VDC.n12823 ;
    wire \ADC_VDC.n13038_cascade_ ;
    wire \ADC_VDC.n20659 ;
    wire \ADC_VDC.n17432_cascade_ ;
    wire \ADC_VDC.n18466 ;
    wire read_buf_11;
    wire read_buf_15;
    wire n11730_cascade_;
    wire adress_6;
    wire \RTD.cfg_buf_6 ;
    wire \RTD.cfg_buf_0 ;
    wire \RTD.n9_cascade_ ;
    wire \RTD.adress_7_N_1340_7_cascade_ ;
    wire \RTD.adress_7 ;
    wire adress_0;
    wire n13181;
    wire \RTD.cfg_buf_5 ;
    wire \RTD.cfg_buf_3 ;
    wire \RTD.n11 ;
    wire \RTD.n7333_cascade_ ;
    wire \RTD.n13_cascade_ ;
    wire \RTD.n11734 ;
    wire \RTD.n7333 ;
    wire \RTD.cfg_tmp_1 ;
    wire \RTD.cfg_tmp_2 ;
    wire \RTD.cfg_tmp_3 ;
    wire \RTD.cfg_tmp_4 ;
    wire \RTD.cfg_tmp_5 ;
    wire \RTD.cfg_tmp_6 ;
    wire \RTD.cfg_tmp_7 ;
    wire \RTD.cfg_tmp_0 ;
    wire \RTD.n13228 ;
    wire \RTD.n15015 ;
    wire read_buf_7;
    wire read_buf_2;
    wire read_buf_3;
    wire n1_adj_1601;
    wire read_buf_4;
    wire n1_adj_1601_cascade_;
    wire read_buf_5;
    wire cmd_rdadctmp_29_adj_1421;
    wire cmd_rdadctmp_30_adj_1420;
    wire DDS_MOSI1;
    wire cmd_rdadctmp_23_adj_1427;
    wire cmd_rdadctmp_24_adj_1426;
    wire cmd_rdadctmp_26_adj_1424;
    wire \CLK_DDS.tmp_buf_1 ;
    wire \CLK_DDS.tmp_buf_2 ;
    wire \CLK_DDS.tmp_buf_3 ;
    wire \CLK_DDS.tmp_buf_4 ;
    wire \CLK_DDS.tmp_buf_5 ;
    wire \CLK_DDS.tmp_buf_6 ;
    wire \CLK_DDS.tmp_buf_7 ;
    wire \CLK_DDS.n9_adj_1395 ;
    wire buf_adcdata_vac_4;
    wire n19_adj_1636_cascade_;
    wire buf_adcdata_iac_4;
    wire buf_data_iac_4;
    wire n22_adj_1637_cascade_;
    wire cmd_rdadctmp_4;
    wire cmd_rdadctmp_5;
    wire cmd_rdadctmp_15;
    wire n19_adj_1631;
    wire buf_adcdata_vac_5;
    wire buf_adcdata_vac_20;
    wire cmd_rdadctmp_29;
    wire cmd_rdadctmp_30;
    wire cmd_rdadctmp_31;
    wire buf_adcdata_vdc_5;
    wire buf_adcdata_vdc_4;
    wire buf_adcdata_vdc_20;
    wire \ADC_VDC.n47 ;
    wire RTD_SCLK;
    wire \RTD.n8 ;
    wire n13309;
    wire RTD_DRDY;
    wire \RTD.adress_7_N_1340_7 ;
    wire \RTD.n16669 ;
    wire \RTD.n16669_cascade_ ;
    wire RTD_CS;
    wire \RTD.n11703 ;
    wire \RTD.cfg_buf_1 ;
    wire \RTD.n12_adj_1397 ;
    wire buf_adcdata_vdc_23;
    wire buf_adcdata_vac_23;
    wire n19_adj_1526_cascade_;
    wire n22076_cascade_;
    wire buf_readRTD_15;
    wire n20;
    wire \RTD.n22370 ;
    wire \RTD.n21323_cascade_ ;
    wire \RTD.n26 ;
    wire \RTD.n21325_cascade_ ;
    wire \RTD.n4 ;
    wire \RTD.n1 ;
    wire \RTD.n1_cascade_ ;
    wire \RTD.n20587 ;
    wire n8_adj_1608;
    wire n21227;
    wire dds_state_0_adj_1454;
    wire \CLK_DDS.n9 ;
    wire \RTD.mode ;
    wire \RTD.n21276_cascade_ ;
    wire \RTD.n21275 ;
    wire \RTD.adc_state_3_N_1368_1 ;
    wire \RTD.adc_state_3_N_1368_1_cascade_ ;
    wire \RTD.n7 ;
    wire \RTD.n20762 ;
    wire \RTD.n11742 ;
    wire n16_adj_1512_cascade_;
    wire cmd_rdadctmp_25_adj_1425;
    wire cmd_rdadctmp_31_adj_1419;
    wire VAC_OSR1;
    wire buf_adcdata_iac_21;
    wire buf_adcdata_iac_23;
    wire VAC_FLT1;
    wire n17_adj_1525;
    wire buf_adcdata_iac_16;
    wire IAC_OSR0;
    wire n22100;
    wire SELIRNG0;
    wire \CLK_DDS.tmp_buf_10 ;
    wire \CLK_DDS.tmp_buf_11 ;
    wire \CLK_DDS.tmp_buf_12 ;
    wire \CLK_DDS.tmp_buf_13 ;
    wire \CLK_DDS.tmp_buf_14 ;
    wire tmp_buf_15_adj_1455;
    wire dds_state_2_adj_1452;
    wire dds_state_1_adj_1453;
    wire \CLK_DDS.tmp_buf_8 ;
    wire \CLK_DDS.tmp_buf_9 ;
    wire \CLK_DDS.n12800 ;
    wire trig_dds1;
    wire ICE_GPMO_1;
    wire IAC_CLK;
    wire cmd_rdadctmp_14;
    wire buf_adcdata_vdc_7;
    wire buf_adcdata_vac_7;
    wire buf_adcdata_iac_7;
    wire n19_adj_1625_cascade_;
    wire buf_data_iac_7;
    wire n22_adj_1626_cascade_;
    wire buf_adcdata_vac_6;
    wire buf_adcdata_vdc_6;
    wire buf_adcdata_iac_6;
    wire n19_adj_1628_cascade_;
    wire buf_data_iac_6;
    wire n22_adj_1629_cascade_;
    wire cmd_rdadctmp_14_adj_1436;
    wire cmd_rdadctmp_15_adj_1435;
    wire n12875_cascade_;
    wire buf_adcdata_vdc_19;
    wire \ADC_VDC.avg_cnt_11 ;
    wire \ADC_VDC.avg_cnt_2 ;
    wire \ADC_VDC.avg_cnt_1 ;
    wire \ADC_VDC.avg_cnt_6 ;
    wire \ADC_VDC.n21 ;
    wire \ADC_VDC.n18479 ;
    wire \ADC_VDC.n21145_cascade_ ;
    wire \ADC_VDC.n13050 ;
    wire read_buf_10;
    wire buf_adcdata_vdc_18;
    wire n20833_cascade_;
    wire read_buf_14;
    wire buf_readRTD_11;
    wire n22214;
    wire \RTD.n10 ;
    wire \RTD.cfg_buf_2 ;
    wire read_buf_0;
    wire \RTD.adc_state_0 ;
    wire adc_state_3_adj_1481;
    wire \RTD.n14717 ;
    wire n16_adj_1524;
    wire \RTD.cfg_buf_4 ;
    wire adc_state_2_adj_1482;
    wire read_buf_6;
    wire n11730;
    wire \RTD.n13192 ;
    wire \RTD.n20631 ;
    wire buf_cfgRTD_7;
    wire \RTD.cfg_buf_7 ;
    wire buf_cfgRTD_3;
    wire cmd_rdadctmp_7_adj_1443;
    wire buf_readRTD_13;
    wire buf_readRTD_10;
    wire buf_cfgRTD_2;
    wire n20834;
    wire adc_state_1_adj_1483;
    wire \RTD.n20656 ;
    wire n12397_cascade_;
    wire buf_adcdata_vac_21;
    wire buf_adcdata_vdc_21;
    wire n22184;
    wire buf_readRTD_12;
    wire n22202;
    wire buf_readRTD_8;
    wire buf_cfgRTD_0;
    wire cmd_rdadctmp_27_adj_1423;
    wire buf_dds1_15;
    wire buf_cfgRTD_4;
    wire n20849;
    wire n22103;
    wire buf_adcdata_iac_17;
    wire buf_data_iac_21;
    wire n20876_cascade_;
    wire n22106;
    wire n20875;
    wire n22022;
    wire buf_dds1_4;
    wire n8_adj_1555_cascade_;
    wire data_index_9_N_216_8;
    wire n8_adj_1555;
    wire n22040;
    wire buf_dds1_9;
    wire buf_dds1_8;
    wire n12383_cascade_;
    wire buf_dds1_10;
    wire n20673;
    wire n11412_cascade_;
    wire AC_ADC_SYNC;
    wire cmd_rdadctmp_12;
    wire cmd_rdadctmp_13;
    wire cmd_rdadctmp_6;
    wire cmd_rdadctmp_7;
    wire cmd_rdadctmp_13_adj_1437;
    wire buf_adcdata_iac_5;
    wire buf_data_iac_5;
    wire n22_adj_1632;
    wire \ADC_VDC.n21718 ;
    wire n12875;
    wire cmd_rdadctmp_0_adj_1479;
    wire \ADC_VDC.cmd_rdadcbuf_0 ;
    wire bfn_10_5_0_;
    wire cmd_rdadctmp_1_adj_1478;
    wire \ADC_VDC.cmd_rdadcbuf_1 ;
    wire \ADC_VDC.n19422 ;
    wire cmd_rdadctmp_2_adj_1477;
    wire \ADC_VDC.cmd_rdadcbuf_2 ;
    wire \ADC_VDC.n19423 ;
    wire cmd_rdadctmp_3_adj_1476;
    wire \ADC_VDC.cmd_rdadcbuf_3 ;
    wire \ADC_VDC.n19424 ;
    wire cmd_rdadctmp_4_adj_1475;
    wire \ADC_VDC.cmd_rdadcbuf_4 ;
    wire \ADC_VDC.n19425 ;
    wire cmd_rdadctmp_5_adj_1474;
    wire \ADC_VDC.cmd_rdadcbuf_5 ;
    wire \ADC_VDC.n19426 ;
    wire cmd_rdadctmp_6_adj_1473;
    wire \ADC_VDC.cmd_rdadcbuf_6 ;
    wire \ADC_VDC.n19427 ;
    wire cmd_rdadctmp_7_adj_1472;
    wire \ADC_VDC.cmd_rdadcbuf_7 ;
    wire \ADC_VDC.n19428 ;
    wire \ADC_VDC.n19429 ;
    wire cmd_rdadctmp_8_adj_1471;
    wire \ADC_VDC.cmd_rdadcbuf_8 ;
    wire bfn_10_6_0_;
    wire cmd_rdadctmp_9_adj_1470;
    wire \ADC_VDC.cmd_rdadcbuf_9 ;
    wire \ADC_VDC.n19430 ;
    wire cmd_rdadctmp_10_adj_1469;
    wire \ADC_VDC.cmd_rdadcbuf_10 ;
    wire \ADC_VDC.n19431 ;
    wire cmd_rdadctmp_11_adj_1468;
    wire \ADC_VDC.n19432 ;
    wire cmd_rdadctmp_12_adj_1467;
    wire cmd_rdadcbuf_12;
    wire \ADC_VDC.n19433 ;
    wire cmd_rdadctmp_13_adj_1466;
    wire cmd_rdadcbuf_13;
    wire \ADC_VDC.n19434 ;
    wire cmd_rdadctmp_14_adj_1465;
    wire cmd_rdadcbuf_14;
    wire \ADC_VDC.n19435 ;
    wire cmd_rdadctmp_15_adj_1464;
    wire cmd_rdadcbuf_15;
    wire \ADC_VDC.n19436 ;
    wire \ADC_VDC.n19437 ;
    wire cmd_rdadctmp_16_adj_1463;
    wire cmd_rdadcbuf_16;
    wire bfn_10_7_0_;
    wire cmd_rdadctmp_17_adj_1462;
    wire cmd_rdadcbuf_17;
    wire \ADC_VDC.n19438 ;
    wire cmd_rdadctmp_18_adj_1461;
    wire cmd_rdadcbuf_18;
    wire \ADC_VDC.n19439 ;
    wire cmd_rdadctmp_19_adj_1460;
    wire cmd_rdadcbuf_19;
    wire \ADC_VDC.n19440 ;
    wire cmd_rdadctmp_20_adj_1459;
    wire \ADC_VDC.n19441 ;
    wire cmd_rdadctmp_21_adj_1458;
    wire cmd_rdadcbuf_21;
    wire \ADC_VDC.n19442 ;
    wire cmd_rdadcbuf_22;
    wire \ADC_VDC.n19443 ;
    wire cmd_rdadcbuf_23;
    wire \ADC_VDC.n19444 ;
    wire \ADC_VDC.n19445 ;
    wire bfn_10_8_0_;
    wire \ADC_VDC.n19446 ;
    wire \ADC_VDC.n19447 ;
    wire \ADC_VDC.n19448 ;
    wire cmd_rdadcbuf_28;
    wire \ADC_VDC.n19449 ;
    wire cmd_rdadcbuf_29;
    wire \ADC_VDC.n19450 ;
    wire cmd_rdadcbuf_30;
    wire \ADC_VDC.n19451 ;
    wire cmd_rdadcbuf_31;
    wire \ADC_VDC.n19452 ;
    wire \ADC_VDC.n19453 ;
    wire cmd_rdadcbuf_32;
    wire bfn_10_9_0_;
    wire \ADC_VDC.n19454 ;
    wire \ADC_VDC.n13038 ;
    wire \ADC_VDC.n14931 ;
    wire cmd_rdadcbuf_34;
    wire \ADC_VDC.n19455 ;
    wire \ADC_VDC.cmd_rdadcbuf_35_N_1139_34 ;
    wire n20824;
    wire n22118;
    wire cmd_rdadctmp_8;
    wire buf_cfgRTD_5;
    wire buf_adcdata_iac_18;
    wire IAC_FLT0;
    wire n20825;
    wire data_index_9_N_216_0;
    wire comm_cmd_5;
    wire comm_cmd_6;
    wire IAC_OSR1;
    wire comm_cmd_4;
    wire buf_dds1_3;
    wire buf_cfgRTD_1;
    wire buf_readRTD_9;
    wire n9_adj_1416;
    wire buf_dds1_0;
    wire n20663_cascade_;
    wire bfn_10_14_0_;
    wire n19384;
    wire n19385;
    wire n19386;
    wire n19387;
    wire n19388;
    wire n19389;
    wire n19390;
    wire n19391;
    wire data_index_8;
    wire n7_adj_1554;
    wire bfn_10_15_0_;
    wire n19392;
    wire buf_dds1_2;
    wire data_index_7;
    wire n8_adj_1557;
    wire n8_adj_1557_cascade_;
    wire n7_adj_1556;
    wire data_index_9_N_216_7;
    wire n8_adj_1553_cascade_;
    wire data_index_9;
    wire ICE_GPMI_0;
    wire n11401;
    wire n20772_cascade_;
    wire n11835_cascade_;
    wire buf_dds0_10;
    wire \SIG_DDS.tmp_buf_10 ;
    wire buf_dds0_13;
    wire \SIG_DDS.tmp_buf_13 ;
    wire \SIG_DDS.tmp_buf_11 ;
    wire \SIG_DDS.tmp_buf_12 ;
    wire \SIG_DDS.tmp_buf_14 ;
    wire buf_dds0_15;
    wire buf_dds0_9;
    wire \SIG_DDS.tmp_buf_9 ;
    wire \SIG_DDS.tmp_buf_6 ;
    wire \SIG_DDS.tmp_buf_5 ;
    wire buf_dds0_2;
    wire buf_dds0_4;
    wire \SIG_DDS.tmp_buf_4 ;
    wire \SIG_DDS.tmp_buf_7 ;
    wire buf_dds0_8;
    wire \SIG_DDS.tmp_buf_8 ;
    wire buf_dds0_1;
    wire \SIG_DDS.tmp_buf_1 ;
    wire \SIG_DDS.tmp_buf_2 ;
    wire buf_dds0_3;
    wire \SIG_DDS.tmp_buf_3 ;
    wire n8_adj_1553;
    wire n7_adj_1552;
    wire data_index_9_N_216_9;
    wire buf_adcdata_vdc_2;
    wire buf_adcdata_vac_2;
    wire buf_adcdata_iac_2;
    wire n19_adj_1646_cascade_;
    wire buf_data_iac_2;
    wire n22_adj_1647_cascade_;
    wire cmd_rdadctmp_10;
    wire buf_adcdata_vdc_3;
    wire n19_adj_1642_cascade_;
    wire buf_data_iac_3;
    wire n22_adj_1643_cascade_;
    wire buf_adcdata_iac_3;
    wire cmd_rdadctmp_11;
    wire buf_adcdata_vac_3;
    wire cmd_rdadctmp_11_adj_1439;
    wire cmd_rdadctmp_12_adj_1438;
    wire buf_data_vac_7;
    wire buf_data_vac_6;
    wire buf_data_vac_5;
    wire cmd_rdadctmp_10_adj_1440;
    wire n30_adj_1480_cascade_;
    wire buf_adcdata_vdc_1;
    wire n19_adj_1491_cascade_;
    wire buf_adcdata_iac_1;
    wire buf_readRTD_14;
    wire cmd_rdadcbuf_26;
    wire cmd_rdadcbuf_25;
    wire cmd_rdadcbuf_24;
    wire cmd_rdadcbuf_27;
    wire cmd_rdadcbuf_11;
    wire cmd_rdadcbuf_33;
    wire n13109;
    wire cmd_rdadcbuf_20;
    wire buf_adcdata_vac_18;
    wire n12411;
    wire buf_cfgRTD_6;
    wire cmd_rdadctmp_27;
    wire buf_adcdata_vac_19;
    wire cmd_rdadctmp_8_adj_1442;
    wire cmd_rdadctmp_9_adj_1441;
    wire buf_adcdata_vdc_15;
    wire buf_adcdata_vac_15;
    wire n22016;
    wire buf_adcdata_vdc_16;
    wire cmd_rdadctmp_23;
    wire cmd_rdadctmp_24;
    wire n20590_cascade_;
    wire buf_adcdata_vac_16;
    wire data_count_0;
    wire bfn_11_11_0_;
    wire data_count_1;
    wire n19345;
    wire data_count_2;
    wire n19346;
    wire data_count_3;
    wire n19347;
    wire data_count_4;
    wire n19348;
    wire data_count_5;
    wire n19349;
    wire data_count_6;
    wire n19350;
    wire data_count_7;
    wire n19351;
    wire n19352;
    wire INVdata_count_i0_i0C_net;
    wire data_count_8;
    wire bfn_11_12_0_;
    wire n19353;
    wire data_count_9;
    wire INVdata_count_i0_i8C_net;
    wire cmd_rdadctmp_16;
    wire buf_adcdata_vdc_8;
    wire buf_adcdata_vac_8;
    wire buf_adcdata_vdc_10;
    wire buf_adcdata_vac_10;
    wire cmd_rdadctmp_17;
    wire cmd_rdadctmp_18;
    wire AMPV_POW;
    wire n23_adj_1536;
    wire cmd_rdadctmp_21_adj_1429;
    wire n7_adj_1531;
    wire cmd_rdadctmp_22_adj_1428;
    wire buf_adcdata_vdc_9;
    wire buf_adcdata_vac_9;
    wire n17411_cascade_;
    wire data_index_9_N_216_5;
    wire n17409;
    wire n17411;
    wire data_index_5;
    wire n8828_cascade_;
    wire data_index_0;
    wire n8_adj_1532;
    wire buf_dds1_13;
    wire buf_dds0_6;
    wire buf_dds1_6;
    wire n11757;
    wire wdtick_cnt_0;
    wire wdtick_cnt_1;
    wire wdtick_cnt_2;
    wire buf_dds0_0;
    wire \SIG_DDS.tmp_buf_0 ;
    wire \SIG_DDS.n12738 ;
    wire EIS_SYNCCLK;
    wire OUT_SYNCCLK;
    wire bfn_12_3_0_;
    wire \ADC_VDC.genclk.n19468 ;
    wire \ADC_VDC.genclk.t0off_2 ;
    wire \ADC_VDC.genclk.n19469 ;
    wire \ADC_VDC.genclk.n19470 ;
    wire \ADC_VDC.genclk.n19471 ;
    wire \ADC_VDC.genclk.n19472 ;
    wire \ADC_VDC.genclk.n19473 ;
    wire \ADC_VDC.genclk.t0off_7 ;
    wire \ADC_VDC.genclk.n19474 ;
    wire \ADC_VDC.genclk.n19475 ;
    wire \INVADC_VDC.genclk.t0off_i0C_net ;
    wire bfn_12_4_0_;
    wire \ADC_VDC.genclk.n19476 ;
    wire \ADC_VDC.genclk.t0off_10 ;
    wire \ADC_VDC.genclk.n19477 ;
    wire \ADC_VDC.genclk.n19478 ;
    wire \ADC_VDC.genclk.t0off_12 ;
    wire \ADC_VDC.genclk.n19479 ;
    wire \ADC_VDC.genclk.n19480 ;
    wire \ADC_VDC.genclk.n19481 ;
    wire \ADC_VDC.genclk.n19482 ;
    wire \INVADC_VDC.genclk.t0off_i8C_net ;
    wire \ADC_VDC.genclk.n11751 ;
    wire n12_adj_1615_cascade_;
    wire n12236_cascade_;
    wire buf_data_vac_0;
    wire buf_data_vac_1;
    wire buf_data_vac_2;
    wire buf_data_vac_3;
    wire buf_data_vac_4;
    wire n12236;
    wire n14801;
    wire n2_adj_1587_cascade_;
    wire comm_buf_5_4;
    wire n21324;
    wire n4_adj_1588_cascade_;
    wire n22136;
    wire n1_adj_1586;
    wire n19006;
    wire n19006_cascade_;
    wire n30_adj_1627;
    wire n30_adj_1630;
    wire n30_adj_1634;
    wire n30_adj_1638;
    wire comm_buf_2_4;
    wire n30_adj_1644;
    wire n30_adj_1648;
    wire cmd_rdadctmp_22_adj_1457;
    wire \ADC_VDC.n10552 ;
    wire \ADC_VDC.cmd_rdadctmp_23 ;
    wire \ADC_VDC.n12915 ;
    wire \ADC_VDC.n20392 ;
    wire \RTD.n17720 ;
    wire buf_adcdata_vac_22;
    wire buf_adcdata_vdc_22;
    wire n22160;
    wire comm_buf_6_4;
    wire n20646;
    wire n14522;
    wire n11918;
    wire cmd_rdadctmp_22;
    wire bfn_12_11_0_;
    wire n19393;
    wire n19394;
    wire n19395;
    wire n19396;
    wire n19397;
    wire n19398;
    wire n19399;
    wire n19400;
    wire bfn_12_12_0_;
    wire n19401;
    wire n19402;
    wire n19403;
    wire n19404;
    wire data_idxvec_13;
    wire n19405;
    wire n19406;
    wire n19407;
    wire n22169_cascade_;
    wire n22079;
    wire n20568_cascade_;
    wire data_idxvec_15;
    wire eis_end;
    wire n26_adj_1528_cascade_;
    wire n22166;
    wire n20742;
    wire acadc_trig;
    wire INVeis_end_309C_net;
    wire n16594_cascade_;
    wire n22196;
    wire n16602_cascade_;
    wire INVeis_state_i0C_net;
    wire n16602;
    wire acadc_skipCount_14;
    wire acadc_skipCount_10;
    wire acadc_skipcnt_0;
    wire bfn_12_16_0_;
    wire INVacadc_skipcnt_i0_i0C_net;
    wire n19369;
    wire n19369_THRU_CRY_0_THRU_CO;
    wire n19369_THRU_CRY_1_THRU_CO;
    wire n19369_THRU_CRY_2_THRU_CO;
    wire n19369_THRU_CRY_3_THRU_CO;
    wire n19369_THRU_CRY_4_THRU_CO;
    wire GNDG0;
    wire n19369_THRU_CRY_5_THRU_CO;
    wire n19369_THRU_CRY_6_THRU_CO;
    wire bfn_12_17_0_;
    wire n19370;
    wire n19371;
    wire n19372;
    wire n19373;
    wire acadc_skipcnt_6;
    wire n19374;
    wire n19375;
    wire n19376;
    wire n19377;
    wire INVacadc_skipcnt_i0_i1C_net;
    wire bfn_12_18_0_;
    wire acadc_skipcnt_10;
    wire n19378;
    wire acadc_skipcnt_11;
    wire n19379;
    wire acadc_skipcnt_12;
    wire n19380;
    wire n19381;
    wire acadc_skipcnt_14;
    wire n19382;
    wire n19383;
    wire INVacadc_skipcnt_i0_i9C_net;
    wire TEST_LED;
    wire \ADC_VDC.genclk.t0off_13 ;
    wire \ADC_VDC.genclk.t0off_3 ;
    wire \ADC_VDC.genclk.t0off_5 ;
    wire \ADC_VDC.genclk.t0off_8 ;
    wire \ADC_VDC.genclk.n27 ;
    wire \ADC_VDC.genclk.n26_cascade_ ;
    wire \ADC_VDC.genclk.n21206_cascade_ ;
    wire \INVADC_VDC.genclk.div_state_i0C_net ;
    wire \ADC_VDC.genclk.t0off_6 ;
    wire \ADC_VDC.genclk.t0off_0 ;
    wire \ADC_VDC.genclk.t0off_4 ;
    wire \ADC_VDC.genclk.t0off_1 ;
    wire \ADC_VDC.genclk.n21208 ;
    wire \ADC_VDC.genclk.t0off_14 ;
    wire \ADC_VDC.genclk.t0off_9 ;
    wire \ADC_VDC.genclk.t0off_15 ;
    wire \ADC_VDC.genclk.t0off_11 ;
    wire \ADC_VDC.genclk.n28 ;
    wire \ADC_VDC.genclk.n21206 ;
    wire \INVADC_VDC.genclk.div_state_i1C_net ;
    wire \ADC_VDC.genclk.n6 ;
    wire \ADC_VDC.genclk.div_state_0 ;
    wire \ADC_VDC.n11766 ;
    wire VDC_SDO;
    wire \ADC_VDC.adc_state_0 ;
    wire \ADC_VDC.n62 ;
    wire adc_state_2;
    wire adc_state_3;
    wire \ADC_VDC.n62_cascade_ ;
    wire \ADC_VDC.adc_state_1 ;
    wire \ADC_VDC.n11 ;
    wire bfn_13_5_0_;
    wire \ADC_VDC.genclk.n19483 ;
    wire \ADC_VDC.genclk.n19484 ;
    wire \ADC_VDC.genclk.n19485 ;
    wire \ADC_VDC.genclk.n19486 ;
    wire \ADC_VDC.genclk.n19487 ;
    wire \ADC_VDC.genclk.n19488 ;
    wire \ADC_VDC.genclk.n19489 ;
    wire \ADC_VDC.genclk.n19490 ;
    wire \INVADC_VDC.genclk.t0on_i0C_net ;
    wire bfn_13_6_0_;
    wire \ADC_VDC.genclk.n19491 ;
    wire \ADC_VDC.genclk.n19492 ;
    wire \ADC_VDC.genclk.n19493 ;
    wire \ADC_VDC.genclk.n19494 ;
    wire \ADC_VDC.genclk.n19495 ;
    wire \ADC_VDC.genclk.n19496 ;
    wire \ADC_VDC.genclk.n19497 ;
    wire \INVADC_VDC.genclk.t0on_i8C_net ;
    wire \ADC_VDC.genclk.div_state_1__N_1275 ;
    wire \ADC_VDC.genclk.n15067 ;
    wire \RTD.bit_cnt_3 ;
    wire \RTD.bit_cnt_1 ;
    wire \RTD.bit_cnt_2 ;
    wire \RTD.bit_cnt_0 ;
    wire \RTD.n11756 ;
    wire \RTD.n15081 ;
    wire n12152_cascade_;
    wire n12_adj_1639;
    wire n12194_cascade_;
    wire buf_adcdata_iac_0;
    wire n22_cascade_;
    wire buf_data_iac_0;
    wire n30_adj_1484_cascade_;
    wire n22_adj_1489;
    wire buf_data_iac_1;
    wire n30_adj_1504_cascade_;
    wire buf_adcdata_vdc_0;
    wire buf_adcdata_vac_0;
    wire n19_adj_1485;
    wire n12110;
    wire n12110_cascade_;
    wire n14780;
    wire data_idxvec_10;
    wire n20905_cascade_;
    wire n20839;
    wire n22148_cascade_;
    wire n22121;
    wire n22151_cascade_;
    wire n20889_cascade_;
    wire buf_data_iac_18;
    wire n20906;
    wire n20670;
    wire n20672;
    wire cmd_rdadctmp_9;
    wire buf_adcdata_vac_1;
    wire n20840;
    wire cmd_rdadctmp_21;
    wire cmd_rdadctmp_20;
    wire n20590;
    wire cmd_rdadctmp_19;
    wire cmd_rdadctmp_25;
    wire n12534;
    wire cmd_rdadctmp_26;
    wire n24_adj_1622_cascade_;
    wire buf_adcdata_vdc_12;
    wire buf_adcdata_vac_12;
    wire n35_cascade_;
    wire iac_raw_buf_N_735;
    wire n17_adj_1645;
    wire adc_state_0;
    wire adc_state_1;
    wire DTRIG_N_919;
    wire n8;
    wire n11354;
    wire n10534_cascade_;
    wire n16598;
    wire n20957;
    wire DTRIG_N_919_adj_1451;
    wire adc_state_1_adj_1417;
    wire ICE_GPMO_0;
    wire auxmode;
    wire acadc_rst_cascade_;
    wire tacadc_rst;
    wire buf_readRTD_7;
    wire n19_adj_1502;
    wire n11_cascade_;
    wire n21099_cascade_;
    wire n13;
    wire INVeis_state_i2C_net;
    wire n11760;
    wire n17430;
    wire acadc_dtrig_v;
    wire acadc_dtrig_i;
    wire n4_adj_1569;
    wire data_index_3;
    wire n8_adj_1563;
    wire n8_adj_1563_cascade_;
    wire n7_adj_1562;
    wire data_index_9_N_216_3;
    wire acadc_skipcnt_5;
    wire acadc_skipcnt_3;
    wire acadc_skipcnt_8;
    wire n20_adj_1617_cascade_;
    wire n17_adj_1612;
    wire n26_adj_1640_cascade_;
    wire n31;
    wire data_index_2;
    wire acadc_skipcnt_15;
    wire acadc_skipcnt_9;
    wire n21;
    wire n24_adj_1537_cascade_;
    wire n23_adj_1624;
    wire n30;
    wire n20789;
    wire eis_state_0;
    wire acadc_rst;
    wire buf_dds1_5;
    wire data_idxvec_14;
    wire eis_end_N_725;
    wire n11670;
    wire n14687;
    wire n10733;
    wire buf_dds0_5;
    wire n27_adj_1551_cascade_;
    wire n25;
    wire n19608_cascade_;
    wire n10_adj_1594;
    wire n26_adj_1543;
    wire n28_adj_1621;
    wire n14_adj_1592;
    wire buf_dds1_14;
    wire buf_dds0_14;
    wire n22115_cascade_;
    wire n22163;
    wire VAC_FLT0;
    wire buf_adcdata_iac_22;
    wire n22112;
    wire n21037;
    wire n23_adj_1534;
    wire n22070_cascade_;
    wire n20856;
    wire n22073_cascade_;
    wire n30_adj_1535_cascade_;
    wire \ADC_VDC.genclk.t0on_6 ;
    wire \ADC_VDC.genclk.t0on_1 ;
    wire \ADC_VDC.genclk.t0on_4 ;
    wire \ADC_VDC.genclk.t0on_0 ;
    wire \ADC_VDC.genclk.n21211_cascade_ ;
    wire \ADC_VDC.genclk.n21205 ;
    wire \ADC_VDC.genclk.t0on_13 ;
    wire \ADC_VDC.genclk.t0on_3 ;
    wire \ADC_VDC.genclk.t0on_5 ;
    wire \ADC_VDC.genclk.t0on_8 ;
    wire \ADC_VDC.genclk.n26_adj_1408 ;
    wire \ADC_VDC.genclk.t0on_14 ;
    wire \ADC_VDC.genclk.t0on_9 ;
    wire \ADC_VDC.genclk.t0on_15 ;
    wire \ADC_VDC.genclk.t0on_11 ;
    wire \ADC_VDC.genclk.n28_adj_1407 ;
    wire \ADC_VDC.genclk.t0on_12 ;
    wire \ADC_VDC.genclk.t0on_2 ;
    wire \ADC_VDC.genclk.t0on_7 ;
    wire \ADC_VDC.genclk.t0on_10 ;
    wire \ADC_VDC.genclk.n27_adj_1409 ;
    wire buf_data_vac_16;
    wire buf_data_vac_20;
    wire comm_buf_3_4;
    wire buf_data_vac_23;
    wire buf_data_vac_22;
    wire buf_data_vac_21;
    wire buf_data_vac_19;
    wire buf_data_vac_18;
    wire buf_data_vac_17;
    wire n12152;
    wire n14787;
    wire n1_cascade_;
    wire comm_buf_2_0;
    wire comm_buf_3_0;
    wire n2;
    wire comm_buf_5_0;
    wire n20970;
    wire n4_adj_1507_cascade_;
    wire n21980;
    wire n21116_cascade_;
    wire n10713;
    wire n12_adj_1602;
    wire buf_data_vac_8;
    wire comm_buf_4_0;
    wire buf_data_vac_15;
    wire buf_data_vac_14;
    wire buf_data_vac_13;
    wire buf_data_vac_12;
    wire comm_buf_4_4;
    wire buf_data_vac_11;
    wire buf_data_vac_10;
    wire buf_data_vac_9;
    wire n12194;
    wire n14794;
    wire n1_adj_1589_cascade_;
    wire comm_buf_6_3;
    wire n21296_cascade_;
    wire n22154;
    wire comm_buf_4_3;
    wire comm_buf_5_3;
    wire n4_adj_1591;
    wire comm_buf_3_3;
    wire comm_buf_2_3;
    wire n2_adj_1590;
    wire n21102_cascade_;
    wire n21_adj_1618;
    wire n16_adj_1599;
    wire data_idxvec_6;
    wire buf_data_iac_14;
    wire n26_adj_1505_cascade_;
    wire n20930_cascade_;
    wire n21962_cascade_;
    wire n21965_cascade_;
    wire buf_adcdata_vdc_14;
    wire buf_adcdata_vac_14;
    wire buf_readRTD_6;
    wire n19_cascade_;
    wire n20954;
    wire acadc_skipCount_6;
    wire n20929;
    wire comm_buf_1_3;
    wire acadc_skipCount_3;
    wire n20884_cascade_;
    wire n20878;
    wire n22124_cascade_;
    wire n22127;
    wire data_idxvec_3;
    wire buf_data_iac_11;
    wire n26_adj_1514_cascade_;
    wire n20885;
    wire buf_readRTD_3;
    wire n20879;
    wire buf_adcdata_vac_11;
    wire buf_adcdata_vdc_11;
    wire n19_adj_1513;
    wire n22178_cascade_;
    wire n22181_cascade_;
    wire n30_adj_1511_cascade_;
    wire data_idxvec_4;
    wire n26_adj_1510;
    wire n19_adj_1509;
    wire buf_readRTD_4;
    wire buf_adcdata_iac_12;
    wire n22010_cascade_;
    wire n16_adj_1508;
    wire n22013;
    wire n12441_cascade_;
    wire n8_adj_1567_cascade_;
    wire data_index_1;
    wire n11835;
    wire n16763;
    wire buf_dds1_1;
    wire buf_adcdata_iac_14;
    wire n16;
    wire n20953;
    wire n10614;
    wire n12312;
    wire VDC_RNG0;
    wire acadc_skipCount_12;
    wire n12383;
    wire acadc_skipcnt_13;
    wire acadc_skipCount_13;
    wire n14;
    wire acadc_skipcnt_1;
    wire acadc_skipcnt_4;
    wire n18_adj_1611;
    wire data_index_4;
    wire n7_adj_1560;
    wire n8_adj_1561;
    wire data_index_9_N_216_4;
    wire n8_adj_1565;
    wire n7_adj_1564;
    wire data_index_9_N_216_2;
    wire n14_adj_1573;
    wire n14_adj_1572;
    wire acadc_skipcnt_7;
    wire acadc_skipcnt_2;
    wire n22_adj_1620;
    wire n9_adj_1415;
    wire n14_adj_1570;
    wire n21048;
    wire n10_adj_1613;
    wire bfn_14_17_0_;
    wire n19498;
    wire n19499;
    wire n19500;
    wire n19501;
    wire n19502;
    wire n10;
    wire n19503;
    wire n19504;
    wire INVdds0_mclkcnt_i7_3783__i0C_net;
    wire secclk_cnt_0;
    wire bfn_14_18_0_;
    wire secclk_cnt_1;
    wire n19509;
    wire secclk_cnt_2;
    wire n19510;
    wire secclk_cnt_3;
    wire n19511;
    wire secclk_cnt_4;
    wire n19512;
    wire secclk_cnt_5;
    wire n19513;
    wire secclk_cnt_6;
    wire n19514;
    wire secclk_cnt_7;
    wire n19515;
    wire n19516;
    wire secclk_cnt_8;
    wire bfn_14_19_0_;
    wire secclk_cnt_9;
    wire n19517;
    wire secclk_cnt_10;
    wire n19518;
    wire secclk_cnt_11;
    wire n19519;
    wire secclk_cnt_12;
    wire n19520;
    wire secclk_cnt_13;
    wire n19521;
    wire secclk_cnt_14;
    wire n19522;
    wire secclk_cnt_15;
    wire n19523;
    wire n19524;
    wire secclk_cnt_16;
    wire bfn_14_20_0_;
    wire secclk_cnt_17;
    wire n19525;
    wire secclk_cnt_18;
    wire n19526;
    wire secclk_cnt_19;
    wire n19527;
    wire secclk_cnt_20;
    wire n19528;
    wire secclk_cnt_21;
    wire n19529;
    wire n19530;
    wire secclk_cnt_22;
    wire n14731;
    wire comm_rx_buf_6;
    wire \ADC_VDC.genclk.div_state_1 ;
    wire VDC_CLK;
    wire \INVADC_VDC.genclk.t_clk_24C_net ;
    wire n21506_cascade_;
    wire n21067;
    wire n23_adj_1538;
    wire n22028;
    wire buf_adcdata_iac_20;
    wire buf_dds0_12;
    wire n22088_cascade_;
    wire buf_dds1_12;
    wire n22091_cascade_;
    wire n22205;
    wire n22031;
    wire n20844_cascade_;
    wire comm_rx_buf_4;
    wire n30_adj_1539_cascade_;
    wire comm_cmd_7;
    wire n20621_cascade_;
    wire n25_adj_1619_cascade_;
    wire \comm_spi.n16869 ;
    wire \INVcomm_spi.data_valid_85C_net ;
    wire n7_adj_1609;
    wire buf_dds1_11;
    wire buf_dds0_11;
    wire buf_adcdata_iac_19;
    wire n22082;
    wire data_idxvec_11;
    wire buf_data_iac_19;
    wire n26_adj_1541_cascade_;
    wire n20837_cascade_;
    wire n22085;
    wire n22094_cascade_;
    wire n20828;
    wire comm_rx_buf_3;
    wire n22097_cascade_;
    wire flagcntwd;
    wire n11406;
    wire n12242_cascade_;
    wire n20599_cascade_;
    wire n5;
    wire IAC_FLT1;
    wire eis_state_1;
    wire buf_data_iac_8;
    wire data_idxvec_12;
    wire n20983;
    wire n12397;
    wire VAC_OSR0;
    wire n21046;
    wire acadc_skipCount_0;
    wire n19_adj_1487;
    wire buf_readRTD_0;
    wire data_idxvec_0;
    wire n20973;
    wire n26_cascade_;
    wire n21998;
    wire n16_adj_1488;
    wire n22004;
    wire n22007_cascade_;
    wire n22001;
    wire n30_adj_1486_cascade_;
    wire comm_buf_1_0;
    wire acadc_skipCount_8;
    wire eis_start;
    wire n21992;
    wire data_idxvec_8;
    wire buf_data_iac_16;
    wire n20917_cascade_;
    wire n21995;
    wire n20919_cascade_;
    wire n22043;
    wire n22019;
    wire n22220_cascade_;
    wire n22223_cascade_;
    wire comm_buf_0_0;
    wire iac_raw_buf_N_737;
    wire bfn_15_13_0_;
    wire n19354;
    wire n19355;
    wire n19356;
    wire n19357;
    wire n19358;
    wire n19359;
    wire n19360;
    wire n19361;
    wire INVdata_cntvec_i0_i0C_net;
    wire bfn_15_14_0_;
    wire n19362;
    wire n19363;
    wire n19364;
    wire n19365;
    wire n19366;
    wire n19367;
    wire n19368;
    wire INVdata_cntvec_i0_i8C_net;
    wire n13473;
    wire n14663;
    wire data_cntvec_14;
    wire data_cntvec_11;
    wire req_data_cnt_14;
    wire n8828;
    wire n8_adj_1559_cascade_;
    wire data_index_9_N_216_6;
    wire n8_adj_1567;
    wire n7_adj_1566;
    wire data_index_9_N_216_1;
    wire data_cntvec_12;
    wire data_cntvec_10;
    wire req_data_cnt_12;
    wire req_data_cnt_10;
    wire n8_adj_1559;
    wire n7_adj_1558;
    wire data_index_6;
    wire \comm_spi.data_tx_7__N_771 ;
    wire bfn_15_16_0_;
    wire n19505;
    wire n19506;
    wire n19507;
    wire n19508;
    wire clk_cnt_0;
    wire clk_cnt_4;
    wire clk_cnt_1;
    wire clk_cnt_3;
    wire n6_cascade_;
    wire clk_cnt_2;
    wire acadc_skipCount_11;
    wire dds0_mclkcnt_3;
    wire dds0_mclkcnt_5;
    wire dds0_mclkcnt_1;
    wire dds0_mclkcnt_4;
    wire dds0_mclkcnt_2;
    wire dds0_mclkcnt_0;
    wire n12_cascade_;
    wire dds0_mclkcnt_7;
    wire n20543;
    wire n20543_cascade_;
    wire dds0_mclkcnt_6;
    wire INVdds0_mclk_304C_net;
    wire buf_data_iac_22;
    wire n21038;
    wire \comm_spi.bit_cnt_3 ;
    wire \comm_spi.bit_cnt_2 ;
    wire \comm_spi.bit_cnt_1 ;
    wire \comm_spi.bit_cnt_0 ;
    wire \INVcomm_spi.bit_cnt_3778__i3C_net ;
    wire n30_adj_1529;
    wire n22109;
    wire n14766;
    wire n21199_cascade_;
    wire n20681_cascade_;
    wire n20599;
    wire n12108_cascade_;
    wire n4_adj_1616;
    wire n11977;
    wire comm_buf_3_6;
    wire comm_buf_2_6;
    wire comm_buf_6_6;
    wire n21329_cascade_;
    wire n21986_cascade_;
    wire n2_adj_1584;
    wire comm_buf_0_6;
    wire n1_adj_1583;
    wire n20621;
    wire n7_cascade_;
    wire comm_buf_2_2;
    wire comm_buf_3_2;
    wire comm_buf_0_2;
    wire n22046_cascade_;
    wire comm_buf_5_2;
    wire comm_buf_4_2;
    wire comm_buf_6_2;
    wire n4_adj_1593_cascade_;
    wire n22049;
    wire n20801_cascade_;
    wire n20596;
    wire n21094;
    wire n21092_cascade_;
    wire n20_adj_1610;
    wire n20883;
    wire n20695_cascade_;
    wire n20881;
    wire n14545_cascade_;
    wire data_idxvec_1;
    wire n26_adj_1522_cascade_;
    wire acadc_skipCount_1;
    wire n22190_cascade_;
    wire n22193_cascade_;
    wire n30_adj_1523_cascade_;
    wire n19_adj_1520;
    wire buf_readRTD_1;
    wire n22064_cascade_;
    wire n16_adj_1519;
    wire n22067;
    wire buf_readRTD_5;
    wire buf_adcdata_iac_13;
    wire n22142_cascade_;
    wire n16_adj_1496;
    wire acadc_skipCount_5;
    wire n22145;
    wire n22133_cascade_;
    wire n30_adj_1499_cascade_;
    wire data_idxvec_5;
    wire n26_adj_1498_cascade_;
    wire n22130;
    wire data_cntvec_8;
    wire data_cntvec_13;
    wire n19_adj_1597_cascade_;
    wire n29_adj_1635_cascade_;
    wire n16_adj_1623;
    wire req_data_cnt_8;
    wire n10534;
    wire n20798;
    wire n22061;
    wire n14730;
    wire clk_RTD;
    wire n23;
    wire n21_adj_1521;
    wire n22_adj_1568_cascade_;
    wire n30_adj_1641;
    wire data_idxvec_9;
    wire buf_data_iac_17;
    wire n20812_cascade_;
    wire comm_buf_0_3;
    wire SELIRNG1;
    wire comm_buf_0_4;
    wire n14_adj_1571;
    wire n14_adj_1549;
    wire n20814;
    wire n22025;
    wire n22232_cascade_;
    wire n22235;
    wire buf_adcdata_vdc_17;
    wire buf_adcdata_vac_17;
    wire n22226;
    wire n22229;
    wire DDS_RNG_0;
    wire acadc_skipCount_9;
    wire n22037;
    wire buf_dds1_7;
    wire buf_dds0_7;
    wire req_data_cnt_11;
    wire n23_adj_1540;
    wire n20836;
    wire n14_adj_1545;
    wire n11931;
    wire n21073_cascade_;
    wire n21072_cascade_;
    wire clk_16MHz;
    wire dds0_mclk;
    wire buf_control_6;
    wire DDS_MCLK;
    wire buf_adcdata_iac_15;
    wire n16_adj_1503;
    wire n20797;
    wire eis_stop;
    wire n22034;
    wire \SIG_DDS.bit_cnt_1 ;
    wire \SIG_DDS.bit_cnt_2 ;
    wire \SIG_DDS.bit_cnt_3 ;
    wire trig_dds0;
    wire n14900;
    wire bit_cnt_0;
    wire tmp_buf_15;
    wire DDS_MOSI;
    wire DDS_CS;
    wire \SIG_DDS.n9_adj_1394 ;
    wire buf_data_iac_20;
    wire n20984;
    wire n17738;
    wire n14146;
    wire comm_state_3_N_436_2;
    wire n15_cascade_;
    wire n12_adj_1649;
    wire comm_buf_4_1;
    wire comm_buf_5_1;
    wire n4_adj_1595_cascade_;
    wire comm_buf_2_1;
    wire comm_buf_3_1;
    wire comm_buf_0_1;
    wire n22052_cascade_;
    wire comm_buf_1_1;
    wire n20807;
    wire n22055_cascade_;
    wire comm_buf_5_5;
    wire comm_buf_3_5;
    wire n17404_cascade_;
    wire n20951_cascade_;
    wire comm_rx_buf_1;
    wire comm_buf_6_1;
    wire n4_adj_1598_cascade_;
    wire n20573;
    wire comm_state_3_N_420_3;
    wire n1272_cascade_;
    wire comm_buf_4_5;
    wire n22175;
    wire n20551;
    wire n11420;
    wire n20551_cascade_;
    wire n20717;
    wire n20575;
    wire n20962;
    wire n14545;
    wire n22238;
    wire n2_adj_1575_cascade_;
    wire n22241_cascade_;
    wire n8_adj_1576;
    wire n1272;
    wire n20697;
    wire n4_adj_1614;
    wire n20668;
    wire n11866;
    wire n14753;
    wire n8_adj_1530;
    wire comm_buf_3_7;
    wire comm_buf_2_7;
    wire n2_adj_1581_cascade_;
    wire n11503;
    wire n14815;
    wire comm_buf_0_7;
    wire n1_adj_1580;
    wire comm_buf_5_7;
    wire comm_buf_4_7;
    wire n20966;
    wire n4_adj_1582_cascade_;
    wire n21968;
    wire comm_buf_1_5;
    wire buf_data_iac_9;
    wire n21270;
    wire n9;
    wire n20663;
    wire n12467_cascade_;
    wire n14_adj_1533;
    wire data_cntvec_6;
    wire data_cntvec_0;
    wire req_data_cnt_0;
    wire n17;
    wire n16_adj_1515;
    wire comm_buf_0_5;
    wire req_data_cnt_6;
    wire req_data_cnt_2;
    wire n22208_cascade_;
    wire acadc_skipCount_2;
    wire n21959;
    wire n22211_cascade_;
    wire comm_rx_buf_2;
    wire n30_adj_1518_cascade_;
    wire comm_buf_1_2;
    wire n12047;
    wire n14773;
    wire n19_adj_1516;
    wire buf_readRTD_2;
    wire n21956;
    wire data_idxvec_2;
    wire data_cntvec_2;
    wire n26_adj_1517;
    wire n14_adj_1550;
    wire n14_adj_1544;
    wire data_cntvec_1;
    wire data_cntvec_4;
    wire req_data_cnt_4;
    wire req_data_cnt_1;
    wire n18;
    wire buf_adcdata_vdc_13;
    wire buf_adcdata_vac_13;
    wire n19_adj_1497;
    wire n14_adj_1579;
    wire acadc_skipCount_15;
    wire n23_adj_1527;
    wire data_cntvec_5;
    wire data_cntvec_3;
    wire req_data_cnt_3;
    wire n20_adj_1596;
    wire comm_buf_1_7;
    wire n14_adj_1546;
    wire n14_adj_1546_cascade_;
    wire n14_adj_1577;
    wire req_data_cnt_13;
    wire data_cntvec_9;
    wire req_data_cnt_15;
    wire data_cntvec_15;
    wire n24;
    wire n14_adj_1574;
    wire req_data_cnt_9;
    wire n12467;
    wire n14_adj_1578;
    wire req_data_cnt_5;
    wire n9321;
    wire n12441;
    wire acadc_skipCount_4;
    wire data_idxvec_7;
    wire data_cntvec_7;
    wire buf_data_iac_15;
    wire n26_adj_1500_cascade_;
    wire n20810_cascade_;
    wire n22058;
    wire acadc_skipCount_7;
    wire req_data_cnt_7;
    wire n20809;
    wire comm_cmd_2;
    wire comm_cmd_3;
    wire comm_cmd_1;
    wire comm_length_1;
    wire comm_length_2;
    wire comm_length_0;
    wire n4;
    wire n14671;
    wire \SIG_DDS.n21331 ;
    wire \SIG_DDS.n10 ;
    wire \SIG_DDS.n9 ;
    wire dds_state_0;
    wire dds_state_2;
    wire dds_state_1;
    wire DDS_SCK;
    wire wdtick_flag;
    wire buf_control_0;
    wire CONT_SD;
    wire n20608;
    wire n23_adj_1501;
    wire n21_adj_1600_cascade_;
    wire n17485;
    wire n18_adj_1633;
    wire \comm_spi.imosi_cascade_ ;
    wire \comm_spi.n22667 ;
    wire \comm_spi.n14630 ;
    wire \comm_spi.n22667_cascade_ ;
    wire comm_rx_buf_0;
    wire comm_rx_buf_0_cascade_;
    wire comm_buf_6_0;
    wire comm_index_2;
    wire comm_buf_2_5;
    wire comm_index_1;
    wire n22172;
    wire comm_rx_buf_5;
    wire comm_buf_6_5;
    wire n2369_cascade_;
    wire n21130_cascade_;
    wire n14_adj_1506;
    wire n3;
    wire n20681;
    wire n3_cascade_;
    wire n2369;
    wire n19655;
    wire ICE_SPI_CE0;
    wire comm_data_vld;
    wire n21129;
    wire n20740;
    wire n11363_cascade_;
    wire n12242;
    wire n12235;
    wire n11869;
    wire n11876;
    wire comm_rx_buf_7;
    wire n12244;
    wire comm_buf_6_7;
    wire THERMOSTAT;
    wire buf_control_7;
    wire n11935;
    wire n19904;
    wire comm_buf_1_4;
    wire n14_adj_1548;
    wire cmd_rdadctmp_20_adj_1430;
    wire comm_buf_1_6;
    wire comm_state_2;
    wire n14_adj_1547;
    wire buf_adcdata_iac_8;
    wire cmd_rdadctmp_16_adj_1434;
    wire n12663;
    wire cmd_rdadctmp_18_adj_1432;
    wire buf_adcdata_iac_10;
    wire cmd_rdadctmp_19_adj_1431;
    wire buf_adcdata_iac_11;
    wire n20584;
    wire adc_state_0_adj_1418;
    wire cmd_rdadctmp_17_adj_1433;
    wire buf_adcdata_iac_9;
    wire buf_data_iac_12;
    wire n21230;
    wire buf_data_iac_13;
    wire n21297;
    wire \comm_spi.DOUT_7__N_747 ;
    wire comm_state_3;
    wire n11377;
    wire \comm_spi.data_tx_7__N_770 ;
    wire comm_buf_5_6;
    wire comm_buf_4_6;
    wire comm_index_0;
    wire n4_adj_1585;
    wire comm_state_1;
    wire comm_state_0;
    wire n9270;
    wire \comm_spi.n22670 ;
    wire \comm_spi.n14631 ;
    wire \comm_spi.n14616 ;
    wire \comm_spi.n14617 ;
    wire \INVcomm_spi.imiso_83_12208_12209_setC_net ;
    wire comm_tx_buf_2;
    wire \comm_spi.imosi ;
    wire \comm_spi.DOUT_7__N_748 ;
    wire \comm_spi.imosi_N_753 ;
    wire \comm_spi.data_tx_7__N_790 ;
    wire \comm_spi.n22685 ;
    wire \comm_spi.data_tx_7__N_772 ;
    wire \comm_spi.n14634 ;
    wire comm_tx_buf_1;
    wire \comm_spi.data_tx_7__N_773 ;
    wire \comm_spi.n22682 ;
    wire \comm_spi.n14638 ;
    wire \comm_spi.n14639 ;
    wire \comm_spi.data_tx_7__N_787 ;
    wire comm_tx_buf_3;
    wire comm_tx_buf_4;
    wire comm_tx_buf_5;
    wire \comm_spi.n22679 ;
    wire \comm_spi.n14642 ;
    wire \comm_spi.n14643 ;
    wire \comm_spi.data_tx_7__N_784 ;
    wire \comm_spi.data_tx_7__N_781 ;
    wire buf_data_iac_23;
    wire n21204;
    wire ICE_SPI_MISO;
    wire \comm_spi.n14621 ;
    wire \INVcomm_spi.MISO_48_12202_12203_resetC_net ;
    wire \comm_spi.n14626 ;
    wire \comm_spi.n14620 ;
    wire \INVcomm_spi.MISO_48_12202_12203_setC_net ;
    wire comm_tx_buf_6;
    wire \comm_spi.n14619 ;
    wire \comm_spi.n14627 ;
    wire \INVcomm_spi.imiso_83_12208_12209_resetC_net ;
    wire \comm_spi.n14624 ;
    wire \comm_spi.n22661 ;
    wire \comm_spi.n14623 ;
    wire \comm_spi.data_tx_7__N_767 ;
    wire comm_tx_buf_7;
    wire \comm_spi.data_tx_7__N_775 ;
    wire \comm_spi.n14635 ;
    wire \comm_spi.data_tx_7__N_793 ;
    wire \comm_spi.n22664 ;
    wire \comm_spi.n14612 ;
    wire \comm_spi.iclk_N_763 ;
    wire \comm_spi.n22688 ;
    wire comm_cmd_0;
    wire buf_data_iac_10;
    wire n21320;
    wire \comm_spi.n14655 ;
    wire \comm_spi.data_tx_7__N_778 ;
    wire \comm_spi.n22673 ;
    wire \comm_spi.n14651 ;
    wire \comm_spi.n14654 ;
    wire \comm_spi.data_tx_7__N_768 ;
    wire \comm_spi.n22676 ;
    wire \comm_spi.n14646 ;
    wire \comm_spi.n14647 ;
    wire \comm_spi.n14650 ;
    wire \comm_spi.data_tx_7__N_769 ;
    wire ICE_SPI_MOSI;
    wire \comm_spi.imosi_N_754 ;
    wire \comm_spi.n14608 ;
    wire \comm_spi.data_tx_7__N_774 ;
    wire ICE_SPI_SCLK;
    wire \comm_spi.n14613 ;
    wire clk_32MHz;
    wire \comm_spi.iclk_N_764 ;
    wire CONSTANT_ONE_NET;
    wire \comm_spi.n14609 ;
    wire \comm_spi.iclk ;
    wire comm_clear;
    wire comm_tx_buf_0;
    wire \comm_spi.data_tx_7__N_796 ;
    wire _gnd_net_;

    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_main.zim_pll_inst .TEST_MODE=1'b0;
    defparam \pll_main.zim_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll_main.zim_pll_inst .FILTER_RANGE=3'b011;
    defparam \pll_main.zim_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_main.zim_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_main.zim_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll_main.zim_pll_inst .DIVR=4'b0000;
    defparam \pll_main.zim_pll_inst .DIVQ=3'b101;
    defparam \pll_main.zim_pll_inst .DIVF=7'b0011111;
    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll_main.zim_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(),
            .REFERENCECLK(N__19205),
            .RESETB(N__57232),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(clk_16MHz),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(clk_32MHz),
            .SCLK(GNDG0));
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged2_physical (
            .RDATA({dangling_wire_0,dangling_wire_1,buf_data_iac_19,dangling_wire_2,dangling_wire_3,dangling_wire_4,buf_data_vac_19,dangling_wire_5,dangling_wire_6,dangling_wire_7,buf_data_iac_18,dangling_wire_8,dangling_wire_9,dangling_wire_10,buf_data_vac_18,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__28217,N__25697,N__27800,N__42278,N__31142,N__38690,N__35978,N__39389,N__42152,N__27350}),
            .WADDR({dangling_wire_13,N__30668,N__30776,N__29600,N__29708,N__29810,N__29924,N__30029,N__30143,N__30251,N__30359}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__40913,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__29429,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__27455,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__29033,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__57931),
            .RE(N__57187),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .WE(N__35539));
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged7_physical (
            .RDATA({dangling_wire_42,dangling_wire_43,buf_data_iac_9,dangling_wire_44,dangling_wire_45,dangling_wire_46,buf_data_vac_9,dangling_wire_47,dangling_wire_48,dangling_wire_49,buf_data_iac_8,dangling_wire_50,dangling_wire_51,dangling_wire_52,buf_data_vac_8,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__28171,N__25660,N__27760,N__42238,N__31108,N__38653,N__35938,N__39352,N__42115,N__27313}),
            .WADDR({dangling_wire_55,N__30631,N__30733,N__29563,N__29668,N__29776,N__29890,N__29998,N__30112,N__30214,N__30322}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__52613,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__30833,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__52153,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__30524,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__57982),
            .RE(N__57379),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .WE(N__35568));
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged1_physical (
            .RDATA({dangling_wire_84,dangling_wire_85,buf_data_iac_21,dangling_wire_86,dangling_wire_87,dangling_wire_88,buf_data_vac_21,dangling_wire_89,dangling_wire_90,dangling_wire_91,buf_data_iac_20,dangling_wire_92,dangling_wire_93,dangling_wire_94,buf_data_vac_20,dangling_wire_95}),
            .RADDR({dangling_wire_96,N__28235,N__25715,N__27818,N__42296,N__31160,N__38708,N__35996,N__39407,N__42170,N__27368}),
            .WADDR({dangling_wire_97,N__30686,N__30794,N__29618,N__29726,N__29828,N__29942,N__30047,N__30161,N__30269,N__30377}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({dangling_wire_114,dangling_wire_115,N__22892,dangling_wire_116,dangling_wire_117,dangling_wire_118,N__25487,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__40382,dangling_wire_122,dangling_wire_123,dangling_wire_124,N__21953,dangling_wire_125}),
            .RCLKE(),
            .RCLK(N__57858),
            .RE(N__57147),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .WE(N__35567));
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged6_physical (
            .RDATA({dangling_wire_126,dangling_wire_127,buf_data_iac_11,dangling_wire_128,dangling_wire_129,dangling_wire_130,buf_data_vac_11,dangling_wire_131,dangling_wire_132,dangling_wire_133,buf_data_iac_10,dangling_wire_134,dangling_wire_135,dangling_wire_136,buf_data_vac_10,dangling_wire_137}),
            .RADDR({dangling_wire_138,N__28183,N__25672,N__27772,N__42250,N__31118,N__38665,N__35950,N__39364,N__42127,N__27325}),
            .WADDR({dangling_wire_139,N__30643,N__30745,N__29575,N__29680,N__29786,N__29900,N__30005,N__30119,N__30226,N__30334}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({dangling_wire_156,dangling_wire_157,N__53237,dangling_wire_158,dangling_wire_159,dangling_wire_160,N__38294,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__51875,dangling_wire_164,dangling_wire_165,dangling_wire_166,N__30473,dangling_wire_167}),
            .RCLKE(),
            .RCLK(N__57980),
            .RE(N__57320),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .WE(N__35566));
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged0_physical (
            .RDATA({dangling_wire_168,dangling_wire_169,buf_data_iac_23,dangling_wire_170,dangling_wire_171,dangling_wire_172,buf_data_vac_23,dangling_wire_173,dangling_wire_174,dangling_wire_175,buf_data_iac_22,dangling_wire_176,dangling_wire_177,dangling_wire_178,buf_data_vac_22,dangling_wire_179}),
            .RADDR({dangling_wire_180,N__28241,N__25721,N__27824,N__42302,N__31166,N__38714,N__36002,N__39413,N__42176,N__27374}),
            .WADDR({dangling_wire_181,N__30692,N__30800,N__29624,N__29732,N__29834,N__29948,N__30053,N__30167,N__30275,N__30383}),
            .MASK({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .WDATA({dangling_wire_198,dangling_wire_199,N__22859,dangling_wire_200,dangling_wire_201,dangling_wire_202,N__22277,dangling_wire_203,dangling_wire_204,dangling_wire_205,N__36820,dangling_wire_206,dangling_wire_207,dangling_wire_208,N__31967,dangling_wire_209}),
            .RCLKE(),
            .RCLK(N__57837),
            .RE(N__57167),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .WE(N__35570));
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged5_physical (
            .RDATA({dangling_wire_210,dangling_wire_211,buf_data_iac_13,dangling_wire_212,dangling_wire_213,dangling_wire_214,buf_data_vac_13,dangling_wire_215,dangling_wire_216,dangling_wire_217,buf_data_iac_12,dangling_wire_218,dangling_wire_219,dangling_wire_220,buf_data_vac_12,dangling_wire_221}),
            .RADDR({dangling_wire_222,N__28195,N__25679,N__27782,N__42260,N__31124,N__38672,N__35960,N__39371,N__42134,N__27332}),
            .WADDR({dangling_wire_223,N__30650,N__30757,N__29582,N__29690,N__29792,N__29906,N__30011,N__30125,N__30233,N__30341}),
            .MASK({dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .WDATA({dangling_wire_240,dangling_wire_241,N__43579,dangling_wire_242,dangling_wire_243,dangling_wire_244,N__46649,dangling_wire_245,dangling_wire_246,dangling_wire_247,N__38165,dangling_wire_248,dangling_wire_249,dangling_wire_250,N__35603,dangling_wire_251}),
            .RCLKE(),
            .RCLK(N__57977),
            .RE(N__57319),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .WE(N__35554));
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged9_physical (
            .RDATA({dangling_wire_252,dangling_wire_253,buf_data_iac_5,dangling_wire_254,dangling_wire_255,dangling_wire_256,buf_data_vac_5,dangling_wire_257,dangling_wire_258,dangling_wire_259,buf_data_iac_4,dangling_wire_260,dangling_wire_261,dangling_wire_262,buf_data_vac_4,dangling_wire_263}),
            .RADDR({dangling_wire_264,N__28192,N__25663,N__27769,N__42247,N__31105,N__38656,N__35947,N__39355,N__42118,N__27316}),
            .WADDR({dangling_wire_265,N__30634,N__30748,N__29566,N__29677,N__29773,N__29887,N__29989,N__30103,N__30217,N__30325}),
            .MASK({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .WDATA({dangling_wire_282,dangling_wire_283,N__25865,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__21977,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__21869,dangling_wire_290,dangling_wire_291,dangling_wire_292,N__21893,dangling_wire_293}),
            .RCLKE(),
            .RCLK(N__57848),
            .RE(N__57380),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .WE(N__35558));
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged4_physical (
            .RDATA({dangling_wire_294,dangling_wire_295,buf_data_iac_15,dangling_wire_296,dangling_wire_297,dangling_wire_298,buf_data_vac_15,dangling_wire_299,dangling_wire_300,dangling_wire_301,buf_data_iac_14,dangling_wire_302,dangling_wire_303,dangling_wire_304,buf_data_vac_14,dangling_wire_305}),
            .RADDR({dangling_wire_306,N__28205,N__25685,N__27788,N__42266,N__31130,N__38678,N__35966,N__39377,N__42140,N__27338}),
            .WADDR({dangling_wire_307,N__30656,N__30764,N__29588,N__29696,N__29798,N__29912,N__30017,N__30131,N__30239,N__30347}),
            .MASK({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323}),
            .WDATA({dangling_wire_324,dangling_wire_325,N__44959,dangling_wire_326,dangling_wire_327,dangling_wire_328,N__29324,dangling_wire_329,dangling_wire_330,dangling_wire_331,N__38366,dangling_wire_332,dangling_wire_333,dangling_wire_334,N__38084,dangling_wire_335}),
            .RCLKE(),
            .RCLK(N__57968),
            .RE(N__57238),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .WE(N__35546));
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged8_physical (
            .RDATA({dangling_wire_336,dangling_wire_337,buf_data_iac_7,dangling_wire_338,dangling_wire_339,dangling_wire_340,buf_data_vac_7,dangling_wire_341,dangling_wire_342,dangling_wire_343,buf_data_iac_6,dangling_wire_344,dangling_wire_345,dangling_wire_346,buf_data_vac_6,dangling_wire_347}),
            .RADDR({dangling_wire_348,N__28204,N__25675,N__27781,N__42259,N__31117,N__38668,N__35959,N__39367,N__42130,N__27328}),
            .WADDR({dangling_wire_349,N__30646,N__30760,N__29578,N__29689,N__29785,N__29899,N__30001,N__30115,N__30229,N__30337}),
            .MASK({dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .WDATA({dangling_wire_366,dangling_wire_367,N__23630,dangling_wire_368,dangling_wire_369,dangling_wire_370,N__23654,dangling_wire_371,dangling_wire_372,dangling_wire_373,N__23771,dangling_wire_374,dangling_wire_375,dangling_wire_376,N__23591,dangling_wire_377}),
            .RCLKE(),
            .RCLK(N__57827),
            .RE(N__57318),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .WE(N__35569));
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged10_physical (
            .RDATA({dangling_wire_378,dangling_wire_379,buf_data_iac_3,dangling_wire_380,dangling_wire_381,dangling_wire_382,buf_data_vac_3,dangling_wire_383,dangling_wire_384,dangling_wire_385,buf_data_iac_2,dangling_wire_386,dangling_wire_387,dangling_wire_388,buf_data_vac_2,dangling_wire_389}),
            .RADDR({dangling_wire_390,N__28229,N__25709,N__27812,N__42290,N__31154,N__38702,N__35990,N__39401,N__42164,N__27362}),
            .WADDR({dangling_wire_391,N__30680,N__30788,N__29612,N__29720,N__29822,N__29936,N__30041,N__30155,N__30263,N__30371}),
            .MASK({dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407}),
            .WDATA({dangling_wire_408,dangling_wire_409,N__28472,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__28802,dangling_wire_413,dangling_wire_414,dangling_wire_415,N__28592,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__28619,dangling_wire_419}),
            .RCLKE(),
            .RCLK(N__57877),
            .RE(N__57148),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .WE(N__35562));
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged3_physical (
            .RDATA({dangling_wire_420,dangling_wire_421,buf_data_iac_17,dangling_wire_422,dangling_wire_423,dangling_wire_424,buf_data_vac_17,dangling_wire_425,dangling_wire_426,dangling_wire_427,buf_data_iac_16,dangling_wire_428,dangling_wire_429,dangling_wire_430,buf_data_vac_16,dangling_wire_431}),
            .RADDR({dangling_wire_432,N__28211,N__25691,N__27794,N__42272,N__31136,N__38684,N__35972,N__39383,N__42146,N__27344}),
            .WADDR({dangling_wire_433,N__30662,N__30770,N__29594,N__29702,N__29804,N__29918,N__30023,N__30137,N__30245,N__30353}),
            .MASK({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .WDATA({dangling_wire_450,dangling_wire_451,N__25556,dangling_wire_452,dangling_wire_453,dangling_wire_454,N__43967,dangling_wire_455,dangling_wire_456,dangling_wire_457,N__22793,dangling_wire_458,dangling_wire_459,dangling_wire_460,N__30410,dangling_wire_461}),
            .RCLKE(),
            .RCLK(N__57954),
            .RE(N__57236),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .WE(N__35506));
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged11_physical (
            .RDATA({dangling_wire_462,dangling_wire_463,buf_data_iac_1,dangling_wire_464,dangling_wire_465,dangling_wire_466,buf_data_vac_1,dangling_wire_467,dangling_wire_468,dangling_wire_469,buf_data_iac_0,dangling_wire_470,dangling_wire_471,dangling_wire_472,buf_data_vac_0,dangling_wire_473}),
            .RADDR({dangling_wire_474,N__28223,N__25703,N__27806,N__42284,N__31148,N__38696,N__35984,N__39395,N__42158,N__27356}),
            .WADDR({dangling_wire_475,N__30674,N__30782,N__29606,N__29714,N__29816,N__29930,N__30035,N__30149,N__30257,N__30365}),
            .MASK({dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .WDATA({dangling_wire_492,dangling_wire_493,N__28913,dangling_wire_494,dangling_wire_495,dangling_wire_496,N__34745,dangling_wire_497,dangling_wire_498,dangling_wire_499,N__34070,dangling_wire_500,dangling_wire_501,dangling_wire_502,N__33964,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__57905),
            .RE(N__57185),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .WE(N__35550));
    IO_PAD ipInertedIOPad_VAC_DRDY_iopad (
            .OE(N__59184),
            .DIN(N__59183),
            .DOUT(N__59182),
            .PACKAGEPIN(VAC_DRDY));
    defparam ipInertedIOPad_VAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_DRDY_preio (
            .PADOEN(N__59184),
            .PADOUT(N__59183),
            .PADIN(N__59182),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT1_iopad (
            .OE(N__59175),
            .DIN(N__59174),
            .DOUT(N__59173),
            .PACKAGEPIN(IAC_FLT1));
    defparam ipInertedIOPad_IAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT1_preio (
            .PADOEN(N__59175),
            .PADOUT(N__59174),
            .PADIN(N__59173),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__41093),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK_iopad (
            .OE(N__59166),
            .DIN(N__59165),
            .DOUT(N__59164),
            .PACKAGEPIN(DDS_SCK));
    defparam ipInertedIOPad_DDS_SCK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK_preio (
            .PADOEN(N__59166),
            .PADOUT(N__59165),
            .PADIN(N__59164),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__50039),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_166_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_166_iopad (
            .OE(N__59157),
            .DIN(N__59156),
            .DOUT(N__59155),
            .PACKAGEPIN(ICE_IOR_166));
    defparam ipInertedIOPad_ICE_IOR_166_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_166_preio (
            .PADOEN(N__59157),
            .PADOUT(N__59156),
            .PADIN(N__59155),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_119_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_119_iopad (
            .OE(N__59148),
            .DIN(N__59147),
            .DOUT(N__59146),
            .PACKAGEPIN(ICE_IOR_119));
    defparam ipInertedIOPad_ICE_IOR_119_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_119_preio (
            .PADOEN(N__59148),
            .PADOUT(N__59147),
            .PADIN(N__59146),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI_iopad (
            .OE(N__59139),
            .DIN(N__59138),
            .DOUT(N__59137),
            .PACKAGEPIN(DDS_MOSI));
    defparam ipInertedIOPad_DDS_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI_preio (
            .PADOEN(N__59139),
            .PADOUT(N__59138),
            .PADIN(N__59137),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44705),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MISO_iopad (
            .OE(N__59130),
            .DIN(N__59129),
            .DOUT(N__59128),
            .PACKAGEPIN(VAC_MISO));
    defparam ipInertedIOPad_VAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_MISO_preio (
            .PADOEN(N__59130),
            .PADOUT(N__59129),
            .PADIN(N__59128),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI1_iopad (
            .OE(N__59121),
            .DIN(N__59120),
            .DOUT(N__59119),
            .PACKAGEPIN(DDS_MOSI1));
    defparam ipInertedIOPad_DDS_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI1_preio (
            .PADOEN(N__59121),
            .PADOUT(N__59120),
            .PADIN(N__59119),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21722),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_146_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_146_iopad (
            .OE(N__59112),
            .DIN(N__59111),
            .DOUT(N__59110),
            .PACKAGEPIN(ICE_IOR_146));
    defparam ipInertedIOPad_ICE_IOR_146_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_146_preio (
            .PADOEN(N__59112),
            .PADOUT(N__59111),
            .PADIN(N__59110),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_CLK_iopad (
            .OE(N__59103),
            .DIN(N__59102),
            .DOUT(N__59101),
            .PACKAGEPIN(VDC_CLK));
    defparam ipInertedIOPad_VDC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_CLK_preio (
            .PADOEN(N__59103),
            .PADOUT(N__59102),
            .PADIN(N__59101),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__40089),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_222_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_222_iopad (
            .OE(N__59094),
            .DIN(N__59093),
            .DOUT(N__59092),
            .PACKAGEPIN(ICE_IOT_222));
    defparam ipInertedIOPad_ICE_IOT_222_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_222_preio (
            .PADOEN(N__59094),
            .PADOUT(N__59093),
            .PADIN(N__59092),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CS_iopad (
            .OE(N__59085),
            .DIN(N__59084),
            .DOUT(N__59083),
            .PACKAGEPIN(IAC_CS));
    defparam ipInertedIOPad_IAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CS_preio (
            .PADOEN(N__59085),
            .PADOUT(N__59084),
            .PADIN(N__59083),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20621),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_18B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_18B_iopad (
            .OE(N__59076),
            .DIN(N__59075),
            .DOUT(N__59074),
            .PACKAGEPIN(ICE_IOL_18B));
    defparam ipInertedIOPad_ICE_IOL_18B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_18B_preio (
            .PADOEN(N__59076),
            .PADOUT(N__59075),
            .PADIN(N__59074),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13A_iopad (
            .OE(N__59067),
            .DIN(N__59066),
            .DOUT(N__59065),
            .PACKAGEPIN(ICE_IOL_13A));
    defparam ipInertedIOPad_ICE_IOL_13A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13A_preio (
            .PADOEN(N__59067),
            .PADOUT(N__59066),
            .PADIN(N__59065),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_81_iopad (
            .OE(N__59058),
            .DIN(N__59057),
            .DOUT(N__59056),
            .PACKAGEPIN(ICE_IOB_81));
    defparam ipInertedIOPad_ICE_IOB_81_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_81_preio (
            .PADOEN(N__59058),
            .PADOUT(N__59057),
            .PADIN(N__59056),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR1_iopad (
            .OE(N__59049),
            .DIN(N__59048),
            .DOUT(N__59047),
            .PACKAGEPIN(VAC_OSR1));
    defparam ipInertedIOPad_VAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR1_preio (
            .PADOEN(N__59049),
            .PADOUT(N__59048),
            .PADIN(N__59047),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22913),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MOSI_iopad (
            .OE(N__59040),
            .DIN(N__59039),
            .DOUT(N__59038),
            .PACKAGEPIN(IAC_MOSI));
    defparam ipInertedIOPad_IAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_MOSI_preio (
            .PADOEN(N__59040),
            .PADOUT(N__59039),
            .PADIN(N__59038),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS1_iopad (
            .OE(N__59031),
            .DIN(N__59030),
            .DOUT(N__59029),
            .PACKAGEPIN(DDS_CS1));
    defparam ipInertedIOPad_DDS_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS1_preio (
            .PADOEN(N__59031),
            .PADOUT(N__59030),
            .PADIN(N__59029),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19841),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4B_iopad (
            .OE(N__59022),
            .DIN(N__59021),
            .DOUT(N__59020),
            .PACKAGEPIN(ICE_IOL_4B));
    defparam ipInertedIOPad_ICE_IOL_4B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4B_preio (
            .PADOEN(N__59022),
            .PADOUT(N__59021),
            .PADIN(N__59020),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_94_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_94_iopad (
            .OE(N__59013),
            .DIN(N__59012),
            .DOUT(N__59011),
            .PACKAGEPIN(ICE_IOB_94));
    defparam ipInertedIOPad_ICE_IOB_94_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_94_preio (
            .PADOEN(N__59013),
            .PADOUT(N__59012),
            .PADIN(N__59011),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CS_iopad (
            .OE(N__59004),
            .DIN(N__59003),
            .DOUT(N__59002),
            .PACKAGEPIN(VAC_CS));
    defparam ipInertedIOPad_VAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CS_preio (
            .PADOEN(N__59004),
            .PADOUT(N__59003),
            .PADIN(N__59002),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19448),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CLK_iopad (
            .OE(N__58995),
            .DIN(N__58994),
            .DOUT(N__58993),
            .PACKAGEPIN(VAC_CLK));
    defparam ipInertedIOPad_VAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CLK_preio (
            .PADOEN(N__58995),
            .PADOUT(N__58994),
            .PADIN(N__58993),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23068),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_CE0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_CE0_iopad (
            .OE(N__58986),
            .DIN(N__58985),
            .DOUT(N__58984),
            .PACKAGEPIN(ICE_SPI_CE0));
    defparam ipInertedIOPad_ICE_SPI_CE0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_CE0_preio (
            .PADOEN(N__58986),
            .PADOUT(N__58985),
            .PADIN(N__58984),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_CE0),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_167_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_167_iopad (
            .OE(N__58977),
            .DIN(N__58976),
            .DOUT(N__58975),
            .PACKAGEPIN(ICE_IOR_167));
    defparam ipInertedIOPad_ICE_IOR_167_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_167_preio (
            .PADOEN(N__58977),
            .PADOUT(N__58976),
            .PADIN(N__58975),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_118_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_118_iopad (
            .OE(N__58968),
            .DIN(N__58967),
            .DOUT(N__58966),
            .PACKAGEPIN(ICE_IOR_118));
    defparam ipInertedIOPad_ICE_IOR_118_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_118_preio (
            .PADOEN(N__58968),
            .PADOUT(N__58967),
            .PADIN(N__58966),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_SDO_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_SDO_iopad (
            .OE(N__58959),
            .DIN(N__58958),
            .DOUT(N__58957),
            .PACKAGEPIN(RTD_SDO));
    defparam ipInertedIOPad_RTD_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_SDO_preio (
            .PADOEN(N__58959),
            .PADOUT(N__58958),
            .PADIN(N__58957),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_SDO),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR0_iopad (
            .OE(N__58950),
            .DIN(N__58949),
            .DOUT(N__58948),
            .PACKAGEPIN(IAC_OSR0));
    defparam ipInertedIOPad_IAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR0_preio (
            .PADOEN(N__58950),
            .PADOUT(N__58949),
            .PADIN(N__58948),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22760),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SCLK_iopad (
            .OE(N__58941),
            .DIN(N__58940),
            .DOUT(N__58939),
            .PACKAGEPIN(VDC_SCLK));
    defparam ipInertedIOPad_VDC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_SCLK_preio (
            .PADOEN(N__58941),
            .PADOUT(N__58940),
            .PADIN(N__58939),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21092),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT1_iopad (
            .OE(N__58932),
            .DIN(N__58931),
            .DOUT(N__58930),
            .PACKAGEPIN(VAC_FLT1));
    defparam ipInertedIOPad_VAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT1_preio (
            .PADOEN(N__58932),
            .PADOUT(N__58931),
            .PADIN(N__58930),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22835),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_MOSI_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_MOSI_iopad (
            .OE(N__58923),
            .DIN(N__58922),
            .DOUT(N__58921),
            .PACKAGEPIN(ICE_SPI_MOSI));
    defparam ipInertedIOPad_ICE_SPI_MOSI_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_MOSI_preio (
            .PADOEN(N__58923),
            .PADOUT(N__58922),
            .PADIN(N__58921),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_MOSI),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_165_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_165_iopad (
            .OE(N__58914),
            .DIN(N__58913),
            .DOUT(N__58912),
            .PACKAGEPIN(ICE_IOR_165));
    defparam ipInertedIOPad_ICE_IOR_165_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_165_preio (
            .PADOEN(N__58914),
            .PADOUT(N__58913),
            .PADIN(N__58912),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_147_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_147_iopad (
            .OE(N__58905),
            .DIN(N__58904),
            .DOUT(N__58903),
            .PACKAGEPIN(ICE_IOR_147));
    defparam ipInertedIOPad_ICE_IOR_147_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_147_preio (
            .PADOEN(N__58905),
            .PADOUT(N__58904),
            .PADIN(N__58903),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_14A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_14A_iopad (
            .OE(N__58896),
            .DIN(N__58895),
            .DOUT(N__58894),
            .PACKAGEPIN(ICE_IOL_14A));
    defparam ipInertedIOPad_ICE_IOL_14A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_14A_preio (
            .PADOEN(N__58896),
            .PADOUT(N__58895),
            .PADIN(N__58894),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13B_iopad (
            .OE(N__58887),
            .DIN(N__58886),
            .DOUT(N__58885),
            .PACKAGEPIN(ICE_IOL_13B));
    defparam ipInertedIOPad_ICE_IOL_13B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13B_preio (
            .PADOEN(N__58887),
            .PADOUT(N__58886),
            .PADIN(N__58885),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_91_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_91_iopad (
            .OE(N__58878),
            .DIN(N__58877),
            .DOUT(N__58876),
            .PACKAGEPIN(ICE_IOB_91));
    defparam ipInertedIOPad_ICE_IOB_91_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_91_preio (
            .PADOEN(N__58878),
            .PADOUT(N__58877),
            .PADIN(N__58876),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_0_iopad (
            .OE(N__58869),
            .DIN(N__58868),
            .DOUT(N__58867),
            .PACKAGEPIN(ICE_GPMO_0));
    defparam ipInertedIOPad_ICE_GPMO_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_0_preio (
            .PADOEN(N__58869),
            .PADOUT(N__58868),
            .PADIN(N__58867),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_0),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_RNG_0_iopad (
            .OE(N__58860),
            .DIN(N__58859),
            .DOUT(N__58858),
            .PACKAGEPIN(DDS_RNG_0));
    defparam ipInertedIOPad_DDS_RNG_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_RNG_0_preio (
            .PADOEN(N__58860),
            .PADOUT(N__58859),
            .PADIN(N__58858),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44660),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_RNG0_iopad (
            .OE(N__58851),
            .DIN(N__58850),
            .DOUT(N__58849),
            .PACKAGEPIN(VDC_RNG0));
    defparam ipInertedIOPad_VDC_RNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_RNG0_preio (
            .PADOEN(N__58851),
            .PADOUT(N__58850),
            .PADIN(N__58849),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39035),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_SCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_SCLK_iopad (
            .OE(N__58842),
            .DIN(N__58841),
            .DOUT(N__58840),
            .PACKAGEPIN(ICE_SPI_SCLK));
    defparam ipInertedIOPad_ICE_SPI_SCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_SCLK_preio (
            .PADOEN(N__58842),
            .PADOUT(N__58841),
            .PADIN(N__58840),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_SCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_152_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_152_iopad (
            .OE(N__58833),
            .DIN(N__58832),
            .DOUT(N__58831),
            .PACKAGEPIN(ICE_IOR_152));
    defparam ipInertedIOPad_ICE_IOR_152_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_152_preio (
            .PADOEN(N__58833),
            .PADOUT(N__58832),
            .PADIN(N__58831),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12A_iopad (
            .OE(N__58824),
            .DIN(N__58823),
            .DOUT(N__58822),
            .PACKAGEPIN(ICE_IOL_12A));
    defparam ipInertedIOPad_ICE_IOL_12A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12A_preio (
            .PADOEN(N__58824),
            .PADOUT(N__58823),
            .PADIN(N__58822),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_DRDY_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_DRDY_iopad (
            .OE(N__58815),
            .DIN(N__58814),
            .DOUT(N__58813),
            .PACKAGEPIN(RTD_DRDY));
    defparam ipInertedIOPad_RTD_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_DRDY_preio (
            .PADOEN(N__58815),
            .PADOUT(N__58814),
            .PADIN(N__58813),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SPI_MISO_iopad (
            .OE(N__58806),
            .DIN(N__58805),
            .DOUT(N__58804),
            .PACKAGEPIN(ICE_SPI_MISO));
    defparam ipInertedIOPad_ICE_SPI_MISO_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_SPI_MISO_preio (
            .PADOEN(N__58806),
            .PADOUT(N__58805),
            .PADIN(N__58804),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__55565),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_177_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_177_iopad (
            .OE(N__58797),
            .DIN(N__58796),
            .DOUT(N__58795),
            .PACKAGEPIN(ICE_IOT_177));
    defparam ipInertedIOPad_ICE_IOT_177_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_177_preio (
            .PADOEN(N__58797),
            .PADOUT(N__58796),
            .PADIN(N__58795),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_141_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_141_iopad (
            .OE(N__58788),
            .DIN(N__58787),
            .DOUT(N__58786),
            .PACKAGEPIN(ICE_IOR_141));
    defparam ipInertedIOPad_ICE_IOR_141_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_141_preio (
            .PADOEN(N__58788),
            .PADOUT(N__58787),
            .PADIN(N__58786),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_102_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_102_iopad (
            .OE(N__58779),
            .DIN(N__58778),
            .DOUT(N__58777),
            .PACKAGEPIN(ICE_IOB_102));
    defparam ipInertedIOPad_ICE_IOB_102_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_102_preio (
            .PADOEN(N__58779),
            .PADOUT(N__58778),
            .PADIN(N__58777),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_2_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_2_iopad (
            .OE(N__58770),
            .DIN(N__58769),
            .DOUT(N__58768),
            .PACKAGEPIN(ICE_GPMO_2));
    defparam ipInertedIOPad_ICE_GPMO_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_2_preio (
            .PADOEN(N__58770),
            .PADOUT(N__58769),
            .PADIN(N__58768),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_2),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_GPMI_0_iopad (
            .OE(N__58761),
            .DIN(N__58760),
            .DOUT(N__58759),
            .PACKAGEPIN(ICE_GPMI_0));
    defparam ipInertedIOPad_ICE_GPMI_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_GPMI_0_preio (
            .PADOEN(N__58761),
            .PADOUT(N__58760),
            .PADIN(N__58759),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27971),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MISO_iopad (
            .OE(N__58752),
            .DIN(N__58751),
            .DOUT(N__58750),
            .PACKAGEPIN(IAC_MISO));
    defparam ipInertedIOPad_IAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_MISO_preio (
            .PADOEN(N__58752),
            .PADOUT(N__58751),
            .PADIN(N__58750),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR0_iopad (
            .OE(N__58743),
            .DIN(N__58742),
            .DOUT(N__58741),
            .PACKAGEPIN(VAC_OSR0));
    defparam ipInertedIOPad_VAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR0_preio (
            .PADOEN(N__58743),
            .PADOUT(N__58742),
            .PADIN(N__58741),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__41339),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MOSI_iopad (
            .OE(N__58734),
            .DIN(N__58733),
            .DOUT(N__58732),
            .PACKAGEPIN(VAC_MOSI));
    defparam ipInertedIOPad_VAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_MOSI_preio (
            .PADOEN(N__58734),
            .PADOUT(N__58733),
            .PADIN(N__58732),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TEST_LED_iopad (
            .OE(N__58725),
            .DIN(N__58724),
            .DOUT(N__58723),
            .PACKAGEPIN(TEST_LED));
    defparam ipInertedIOPad_TEST_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_TEST_LED_preio (
            .PADOEN(N__58725),
            .PADOUT(N__58724),
            .PADIN(N__58723),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32741),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_148_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_148_iopad (
            .OE(N__58716),
            .DIN(N__58715),
            .DOUT(N__58714),
            .PACKAGEPIN(ICE_IOR_148));
    defparam ipInertedIOPad_ICE_IOR_148_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_148_preio (
            .PADOEN(N__58716),
            .PADOUT(N__58715),
            .PADIN(N__58714),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_STAT_COMM_iopad (
            .OE(N__58707),
            .DIN(N__58706),
            .DOUT(N__58705),
            .PACKAGEPIN(STAT_COMM));
    defparam ipInertedIOPad_STAT_COMM_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_STAT_COMM_preio (
            .PADOEN(N__58707),
            .PADOUT(N__58706),
            .PADIN(N__58705),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19190),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SYSCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SYSCLK_iopad (
            .OE(N__58698),
            .DIN(N__58697),
            .DOUT(N__58696),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ipInertedIOPad_ICE_SYSCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SYSCLK_preio (
            .PADOEN(N__58698),
            .PADOUT(N__58697),
            .PADIN(N__58696),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SYSCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_161_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_161_iopad (
            .OE(N__58689),
            .DIN(N__58688),
            .DOUT(N__58687),
            .PACKAGEPIN(ICE_IOR_161));
    defparam ipInertedIOPad_ICE_IOR_161_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_161_preio (
            .PADOEN(N__58689),
            .PADOUT(N__58688),
            .PADIN(N__58687),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_95_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_95_iopad (
            .OE(N__58680),
            .DIN(N__58679),
            .DOUT(N__58678),
            .PACKAGEPIN(ICE_IOB_95));
    defparam ipInertedIOPad_ICE_IOB_95_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_95_preio (
            .PADOEN(N__58680),
            .PADOUT(N__58679),
            .PADIN(N__58678),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_82_iopad (
            .OE(N__58671),
            .DIN(N__58670),
            .DOUT(N__58669),
            .PACKAGEPIN(ICE_IOB_82));
    defparam ipInertedIOPad_ICE_IOB_82_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_82_preio (
            .PADOEN(N__58671),
            .PADOUT(N__58670),
            .PADIN(N__58669),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_104_iopad (
            .OE(N__58662),
            .DIN(N__58661),
            .DOUT(N__58660),
            .PACKAGEPIN(ICE_IOB_104));
    defparam ipInertedIOPad_ICE_IOB_104_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_104_preio (
            .PADOEN(N__58662),
            .PADOUT(N__58661),
            .PADIN(N__58660),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CLK_iopad (
            .OE(N__58653),
            .DIN(N__58652),
            .DOUT(N__58651),
            .PACKAGEPIN(IAC_CLK));
    defparam ipInertedIOPad_IAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CLK_preio (
            .PADOEN(N__58653),
            .PADOUT(N__58652),
            .PADIN(N__58651),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23075),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS_iopad (
            .OE(N__58644),
            .DIN(N__58643),
            .DOUT(N__58642),
            .PACKAGEPIN(DDS_CS));
    defparam ipInertedIOPad_DDS_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS_preio (
            .PADOEN(N__58644),
            .PADOUT(N__58643),
            .PADIN(N__58642),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__45278),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG0_iopad (
            .OE(N__58635),
            .DIN(N__58634),
            .DOUT(N__58633),
            .PACKAGEPIN(SELIRNG0));
    defparam ipInertedIOPad_SELIRNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG0_preio (
            .PADOEN(N__58635),
            .PADOUT(N__58634),
            .PADIN(N__58633),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23024),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SDI_iopad (
            .OE(N__58626),
            .DIN(N__58625),
            .DOUT(N__58624),
            .PACKAGEPIN(RTD_SDI));
    defparam ipInertedIOPad_RTD_SDI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SDI_preio (
            .PADOEN(N__58626),
            .PADOUT(N__58625),
            .PADIN(N__58624),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20348),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_221_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_221_iopad (
            .OE(N__58617),
            .DIN(N__58616),
            .DOUT(N__58615),
            .PACKAGEPIN(ICE_IOT_221));
    defparam ipInertedIOPad_ICE_IOT_221_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_221_preio (
            .PADOEN(N__58617),
            .PADOUT(N__58616),
            .PADIN(N__58615),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_197_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_197_iopad (
            .OE(N__58608),
            .DIN(N__58607),
            .DOUT(N__58606),
            .PACKAGEPIN(ICE_IOT_197));
    defparam ipInertedIOPad_ICE_IOT_197_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_197_preio (
            .PADOEN(N__58608),
            .PADOUT(N__58607),
            .PADIN(N__58606),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK_iopad (
            .OE(N__58599),
            .DIN(N__58598),
            .DOUT(N__58597),
            .PACKAGEPIN(DDS_MCLK));
    defparam ipInertedIOPad_DDS_MCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK_preio (
            .PADOEN(N__58599),
            .PADOUT(N__58598),
            .PADIN(N__58597),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44984),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SCLK_iopad (
            .OE(N__58590),
            .DIN(N__58589),
            .DOUT(N__58588),
            .PACKAGEPIN(RTD_SCLK));
    defparam ipInertedIOPad_RTD_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SCLK_preio (
            .PADOEN(N__58590),
            .PADOUT(N__58589),
            .PADIN(N__58588),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22205),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_CS_iopad (
            .OE(N__58581),
            .DIN(N__58580),
            .DOUT(N__58579),
            .PACKAGEPIN(RTD_CS));
    defparam ipInertedIOPad_RTD_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_CS_preio (
            .PADOEN(N__58581),
            .PADOUT(N__58580),
            .PADIN(N__58579),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22355),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_137_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_137_iopad (
            .OE(N__58572),
            .DIN(N__58571),
            .DOUT(N__58570),
            .PACKAGEPIN(ICE_IOR_137));
    defparam ipInertedIOPad_ICE_IOR_137_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_137_preio (
            .PADOEN(N__58572),
            .PADOUT(N__58571),
            .PADIN(N__58570),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR1_iopad (
            .OE(N__58563),
            .DIN(N__58562),
            .DOUT(N__58561),
            .PACKAGEPIN(IAC_OSR1));
    defparam ipInertedIOPad_IAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR1_preio (
            .PADOEN(N__58563),
            .PADOUT(N__58562),
            .PADIN(N__58561),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27713),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT0_iopad (
            .OE(N__58554),
            .DIN(N__58553),
            .DOUT(N__58552),
            .PACKAGEPIN(VAC_FLT0));
    defparam ipInertedIOPad_VAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT0_preio (
            .PADOEN(N__58554),
            .PADOUT(N__58553),
            .PADIN(N__58552),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36869),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_144_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_144_iopad (
            .OE(N__58545),
            .DIN(N__58544),
            .DOUT(N__58543),
            .PACKAGEPIN(ICE_IOR_144));
    defparam ipInertedIOPad_ICE_IOR_144_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_144_preio (
            .PADOEN(N__58545),
            .PADOUT(N__58544),
            .PADIN(N__58543),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_128_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_128_iopad (
            .OE(N__58536),
            .DIN(N__58535),
            .DOUT(N__58534),
            .PACKAGEPIN(ICE_IOR_128));
    defparam ipInertedIOPad_ICE_IOR_128_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_128_preio (
            .PADOEN(N__58536),
            .PADOUT(N__58535),
            .PADIN(N__58534),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_1_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_1_iopad (
            .OE(N__58527),
            .DIN(N__58526),
            .DOUT(N__58525),
            .PACKAGEPIN(ICE_GPMO_1));
    defparam ipInertedIOPad_ICE_GPMO_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_1_preio (
            .PADOEN(N__58527),
            .PADOUT(N__58526),
            .PADIN(N__58525),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_1),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_SCLK_iopad (
            .OE(N__58518),
            .DIN(N__58517),
            .DOUT(N__58516),
            .PACKAGEPIN(IAC_SCLK));
    defparam ipInertedIOPad_IAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_SCLK_preio (
            .PADOEN(N__58518),
            .PADOUT(N__58517),
            .PADIN(N__58516),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20021),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_EIS_SYNCCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_EIS_SYNCCLK_iopad (
            .OE(N__58509),
            .DIN(N__58508),
            .DOUT(N__58507),
            .PACKAGEPIN(EIS_SYNCCLK));
    defparam ipInertedIOPad_EIS_SYNCCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_EIS_SYNCCLK_preio (
            .PADOEN(N__58509),
            .PADOUT(N__58508),
            .PADIN(N__58507),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(EIS_SYNCCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_139_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_139_iopad (
            .OE(N__58500),
            .DIN(N__58499),
            .DOUT(N__58498),
            .PACKAGEPIN(ICE_IOR_139));
    defparam ipInertedIOPad_ICE_IOR_139_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_139_preio (
            .PADOEN(N__58500),
            .PADOUT(N__58499),
            .PADIN(N__58498),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4A_iopad (
            .OE(N__58491),
            .DIN(N__58490),
            .DOUT(N__58489),
            .PACKAGEPIN(ICE_IOL_4A));
    defparam ipInertedIOPad_ICE_IOL_4A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4A_preio (
            .PADOEN(N__58491),
            .PADOUT(N__58490),
            .PADIN(N__58489),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_SCLK_iopad (
            .OE(N__58482),
            .DIN(N__58481),
            .DOUT(N__58480),
            .PACKAGEPIN(VAC_SCLK));
    defparam ipInertedIOPad_VAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_SCLK_preio (
            .PADOEN(N__58482),
            .PADOUT(N__58481),
            .PADIN(N__58480),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19478),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_THERMOSTAT_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_THERMOSTAT_iopad (
            .OE(N__58473),
            .DIN(N__58472),
            .DOUT(N__58471),
            .PACKAGEPIN(THERMOSTAT));
    defparam ipInertedIOPad_THERMOSTAT_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_THERMOSTAT_preio (
            .PADOEN(N__58473),
            .PADOUT(N__58472),
            .PADIN(N__58471),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(THERMOSTAT),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_164_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_164_iopad (
            .OE(N__58464),
            .DIN(N__58463),
            .DOUT(N__58462),
            .PACKAGEPIN(ICE_IOR_164));
    defparam ipInertedIOPad_ICE_IOR_164_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_164_preio (
            .PADOEN(N__58464),
            .PADOUT(N__58463),
            .PADIN(N__58462),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_103_iopad (
            .OE(N__58455),
            .DIN(N__58454),
            .DOUT(N__58453),
            .PACKAGEPIN(ICE_IOB_103));
    defparam ipInertedIOPad_ICE_IOB_103_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_103_preio (
            .PADOEN(N__58455),
            .PADOUT(N__58454),
            .PADIN(N__58453),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_OUT_SYNCCLK_iopad (
            .OE(N__58446),
            .DIN(N__58445),
            .DOUT(N__58444),
            .PACKAGEPIN(OUT_SYNCCLK));
    defparam ipInertedIOPad_OUT_SYNCCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_OUT_SYNCCLK_preio (
            .PADOEN(N__58446),
            .PADOUT(N__58445),
            .PADIN(N__58444),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31346),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AMPV_POW_iopad (
            .OE(N__58437),
            .DIN(N__58436),
            .DOUT(N__58435),
            .PACKAGEPIN(AMPV_POW));
    defparam ipInertedIOPad_AMPV_POW_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AMPV_POW_preio (
            .PADOEN(N__58437),
            .PADOUT(N__58436),
            .PADIN(N__58435),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30956),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SDO_iopad (
            .OE(N__58428),
            .DIN(N__58427),
            .DOUT(N__58426),
            .PACKAGEPIN(VDC_SDO));
    defparam ipInertedIOPad_VDC_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDC_SDO_preio (
            .PADOEN(N__58428),
            .PADOUT(N__58427),
            .PADIN(N__58426),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VDC_SDO),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_174_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_174_iopad (
            .OE(N__58419),
            .DIN(N__58418),
            .DOUT(N__58417),
            .PACKAGEPIN(ICE_IOT_174));
    defparam ipInertedIOPad_ICE_IOT_174_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_174_preio (
            .PADOEN(N__58419),
            .PADOUT(N__58418),
            .PADIN(N__58417),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_140_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_140_iopad (
            .OE(N__58410),
            .DIN(N__58409),
            .DOUT(N__58408),
            .PACKAGEPIN(ICE_IOR_140));
    defparam ipInertedIOPad_ICE_IOR_140_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_140_preio (
            .PADOEN(N__58410),
            .PADOUT(N__58409),
            .PADIN(N__58408),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_96_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_96_iopad (
            .OE(N__58401),
            .DIN(N__58400),
            .DOUT(N__58399),
            .PACKAGEPIN(ICE_IOB_96));
    defparam ipInertedIOPad_ICE_IOB_96_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_96_preio (
            .PADOEN(N__58401),
            .PADOUT(N__58400),
            .PADIN(N__58399),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CONT_SD_iopad (
            .OE(N__58392),
            .DIN(N__58391),
            .DOUT(N__58390),
            .PACKAGEPIN(CONT_SD));
    defparam ipInertedIOPad_CONT_SD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_CONT_SD_preio (
            .PADOEN(N__58392),
            .PADOUT(N__58391),
            .PADIN(N__58390),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__49952),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AC_ADC_SYNC_iopad (
            .OE(N__58383),
            .DIN(N__58382),
            .DOUT(N__58381),
            .PACKAGEPIN(AC_ADC_SYNC));
    defparam ipInertedIOPad_AC_ADC_SYNC_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AC_ADC_SYNC_preio (
            .PADOEN(N__58383),
            .PADOUT(N__58382),
            .PADIN(N__58381),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25766),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG1_iopad (
            .OE(N__58374),
            .DIN(N__58373),
            .DOUT(N__58372),
            .PACKAGEPIN(SELIRNG1));
    defparam ipInertedIOPad_SELIRNG1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG1_preio (
            .PADOEN(N__58374),
            .PADOUT(N__58373),
            .PADIN(N__58372),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44201),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12B_iopad (
            .OE(N__58365),
            .DIN(N__58364),
            .DOUT(N__58363),
            .PACKAGEPIN(ICE_IOL_12B));
    defparam ipInertedIOPad_ICE_IOL_12B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12B_preio (
            .PADOEN(N__58365),
            .PADOUT(N__58364),
            .PADIN(N__58363),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_160_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_160_iopad (
            .OE(N__58356),
            .DIN(N__58355),
            .DOUT(N__58354),
            .PACKAGEPIN(ICE_IOR_160));
    defparam ipInertedIOPad_ICE_IOR_160_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_160_preio (
            .PADOEN(N__58356),
            .PADOUT(N__58355),
            .PADIN(N__58354),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_136_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_136_iopad (
            .OE(N__58347),
            .DIN(N__58346),
            .DOUT(N__58345),
            .PACKAGEPIN(ICE_IOR_136));
    defparam ipInertedIOPad_ICE_IOR_136_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_136_preio (
            .PADOEN(N__58347),
            .PADOUT(N__58346),
            .PADIN(N__58345),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK1_iopad (
            .OE(N__58338),
            .DIN(N__58337),
            .DOUT(N__58336),
            .PACKAGEPIN(DDS_MCLK1));
    defparam ipInertedIOPad_DDS_MCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK1_preio (
            .PADOEN(N__58338),
            .PADOUT(N__58337),
            .PADIN(N__58336),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20738),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_198_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_198_iopad (
            .OE(N__58329),
            .DIN(N__58328),
            .DOUT(N__58327),
            .PACKAGEPIN(ICE_IOT_198));
    defparam ipInertedIOPad_ICE_IOT_198_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_198_preio (
            .PADOEN(N__58329),
            .PADOUT(N__58328),
            .PADIN(N__58327),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_173_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_173_iopad (
            .OE(N__58320),
            .DIN(N__58319),
            .DOUT(N__58318),
            .PACKAGEPIN(ICE_IOT_173));
    defparam ipInertedIOPad_ICE_IOT_173_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_173_preio (
            .PADOEN(N__58320),
            .PADOUT(N__58319),
            .PADIN(N__58318),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_DRDY_iopad (
            .OE(N__58311),
            .DIN(N__58310),
            .DOUT(N__58309),
            .PACKAGEPIN(IAC_DRDY));
    defparam ipInertedIOPad_IAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_DRDY_preio (
            .PADOEN(N__58311),
            .PADOUT(N__58310),
            .PADIN(N__58309),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_DRDY),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_178_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_178_iopad (
            .OE(N__58302),
            .DIN(N__58301),
            .DOUT(N__58300),
            .PACKAGEPIN(ICE_IOT_178));
    defparam ipInertedIOPad_ICE_IOT_178_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_178_preio (
            .PADOEN(N__58302),
            .PADOUT(N__58301),
            .PADIN(N__58300),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_138_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_138_iopad (
            .OE(N__58293),
            .DIN(N__58292),
            .DOUT(N__58291),
            .PACKAGEPIN(ICE_IOR_138));
    defparam ipInertedIOPad_ICE_IOR_138_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_138_preio (
            .PADOEN(N__58293),
            .PADOUT(N__58292),
            .PADIN(N__58291),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_120_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_120_iopad (
            .OE(N__58284),
            .DIN(N__58283),
            .DOUT(N__58282),
            .PACKAGEPIN(ICE_IOR_120));
    defparam ipInertedIOPad_ICE_IOR_120_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_120_preio (
            .PADOEN(N__58284),
            .PADOUT(N__58283),
            .PADIN(N__58282),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT0_iopad (
            .OE(N__58275),
            .DIN(N__58274),
            .DOUT(N__58273),
            .PACKAGEPIN(IAC_FLT0));
    defparam ipInertedIOPad_IAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT0_preio (
            .PADOEN(N__58275),
            .PADOUT(N__58274),
            .PADIN(N__58273),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27416),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK1_iopad (
            .OE(N__58266),
            .DIN(N__58265),
            .DOUT(N__58264),
            .PACKAGEPIN(DDS_SCK1));
    defparam ipInertedIOPad_DDS_SCK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK1_preio (
            .PADOEN(N__58266),
            .PADOUT(N__58265),
            .PADIN(N__58264),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19883),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    SRMux I__14593 (
            .O(N__58247),
            .I(N__58244));
    LocalMux I__14592 (
            .O(N__58244),
            .I(\comm_spi.data_tx_7__N_768 ));
    InMux I__14591 (
            .O(N__58241),
            .I(N__58238));
    LocalMux I__14590 (
            .O(N__58238),
            .I(N__58234));
    InMux I__14589 (
            .O(N__58237),
            .I(N__58231));
    Span4Mux_v I__14588 (
            .O(N__58234),
            .I(N__58228));
    LocalMux I__14587 (
            .O(N__58231),
            .I(N__58225));
    Span4Mux_v I__14586 (
            .O(N__58228),
            .I(N__58221));
    Span4Mux_v I__14585 (
            .O(N__58225),
            .I(N__58218));
    InMux I__14584 (
            .O(N__58224),
            .I(N__58215));
    Odrv4 I__14583 (
            .O(N__58221),
            .I(\comm_spi.n22676 ));
    Odrv4 I__14582 (
            .O(N__58218),
            .I(\comm_spi.n22676 ));
    LocalMux I__14581 (
            .O(N__58215),
            .I(\comm_spi.n22676 ));
    InMux I__14580 (
            .O(N__58208),
            .I(N__58204));
    InMux I__14579 (
            .O(N__58207),
            .I(N__58201));
    LocalMux I__14578 (
            .O(N__58204),
            .I(N__58198));
    LocalMux I__14577 (
            .O(N__58201),
            .I(\comm_spi.n14646 ));
    Odrv4 I__14576 (
            .O(N__58198),
            .I(\comm_spi.n14646 ));
    InMux I__14575 (
            .O(N__58193),
            .I(N__58189));
    InMux I__14574 (
            .O(N__58192),
            .I(N__58186));
    LocalMux I__14573 (
            .O(N__58189),
            .I(\comm_spi.n14647 ));
    LocalMux I__14572 (
            .O(N__58186),
            .I(\comm_spi.n14647 ));
    InMux I__14571 (
            .O(N__58181),
            .I(N__58178));
    LocalMux I__14570 (
            .O(N__58178),
            .I(N__58174));
    InMux I__14569 (
            .O(N__58177),
            .I(N__58171));
    Odrv4 I__14568 (
            .O(N__58174),
            .I(\comm_spi.n14650 ));
    LocalMux I__14567 (
            .O(N__58171),
            .I(\comm_spi.n14650 ));
    SRMux I__14566 (
            .O(N__58166),
            .I(N__58163));
    LocalMux I__14565 (
            .O(N__58163),
            .I(N__58160));
    Span4Mux_h I__14564 (
            .O(N__58160),
            .I(N__58157));
    Odrv4 I__14563 (
            .O(N__58157),
            .I(\comm_spi.data_tx_7__N_769 ));
    InMux I__14562 (
            .O(N__58154),
            .I(N__58149));
    InMux I__14561 (
            .O(N__58153),
            .I(N__58146));
    InMux I__14560 (
            .O(N__58152),
            .I(N__58143));
    LocalMux I__14559 (
            .O(N__58149),
            .I(N__58136));
    LocalMux I__14558 (
            .O(N__58146),
            .I(N__58136));
    LocalMux I__14557 (
            .O(N__58143),
            .I(N__58136));
    Span4Mux_v I__14556 (
            .O(N__58136),
            .I(N__58132));
    InMux I__14555 (
            .O(N__58135),
            .I(N__58129));
    Span4Mux_h I__14554 (
            .O(N__58132),
            .I(N__58125));
    LocalMux I__14553 (
            .O(N__58129),
            .I(N__58122));
    InMux I__14552 (
            .O(N__58128),
            .I(N__58119));
    Sp12to4 I__14551 (
            .O(N__58125),
            .I(N__58116));
    Span4Mux_h I__14550 (
            .O(N__58122),
            .I(N__58113));
    LocalMux I__14549 (
            .O(N__58119),
            .I(N__58110));
    Span12Mux_s6_h I__14548 (
            .O(N__58116),
            .I(N__58103));
    Sp12to4 I__14547 (
            .O(N__58113),
            .I(N__58103));
    Span12Mux_v I__14546 (
            .O(N__58110),
            .I(N__58103));
    Span12Mux_v I__14545 (
            .O(N__58103),
            .I(N__58100));
    Odrv12 I__14544 (
            .O(N__58100),
            .I(ICE_SPI_MOSI));
    SRMux I__14543 (
            .O(N__58097),
            .I(N__58094));
    LocalMux I__14542 (
            .O(N__58094),
            .I(N__58091));
    Span4Mux_h I__14541 (
            .O(N__58091),
            .I(N__58088));
    Odrv4 I__14540 (
            .O(N__58088),
            .I(\comm_spi.imosi_N_754 ));
    InMux I__14539 (
            .O(N__58085),
            .I(N__58081));
    InMux I__14538 (
            .O(N__58084),
            .I(N__58078));
    LocalMux I__14537 (
            .O(N__58081),
            .I(N__58073));
    LocalMux I__14536 (
            .O(N__58078),
            .I(N__58073));
    Span4Mux_h I__14535 (
            .O(N__58073),
            .I(N__58070));
    Odrv4 I__14534 (
            .O(N__58070),
            .I(\comm_spi.n14608 ));
    SRMux I__14533 (
            .O(N__58067),
            .I(N__58064));
    LocalMux I__14532 (
            .O(N__58064),
            .I(N__58061));
    Span4Mux_h I__14531 (
            .O(N__58061),
            .I(N__58058));
    Odrv4 I__14530 (
            .O(N__58058),
            .I(\comm_spi.data_tx_7__N_774 ));
    InMux I__14529 (
            .O(N__58055),
            .I(N__58051));
    InMux I__14528 (
            .O(N__58054),
            .I(N__58048));
    LocalMux I__14527 (
            .O(N__58051),
            .I(N__58045));
    LocalMux I__14526 (
            .O(N__58048),
            .I(N__58042));
    Span4Mux_v I__14525 (
            .O(N__58045),
            .I(N__58038));
    Span4Mux_v I__14524 (
            .O(N__58042),
            .I(N__58035));
    InMux I__14523 (
            .O(N__58041),
            .I(N__58032));
    Span4Mux_h I__14522 (
            .O(N__58038),
            .I(N__58025));
    Span4Mux_v I__14521 (
            .O(N__58035),
            .I(N__58025));
    LocalMux I__14520 (
            .O(N__58032),
            .I(N__58022));
    InMux I__14519 (
            .O(N__58031),
            .I(N__58019));
    InMux I__14518 (
            .O(N__58030),
            .I(N__58016));
    Sp12to4 I__14517 (
            .O(N__58025),
            .I(N__58013));
    Sp12to4 I__14516 (
            .O(N__58022),
            .I(N__58006));
    LocalMux I__14515 (
            .O(N__58019),
            .I(N__58006));
    LocalMux I__14514 (
            .O(N__58016),
            .I(N__58006));
    Span12Mux_s8_h I__14513 (
            .O(N__58013),
            .I(N__58001));
    Span12Mux_v I__14512 (
            .O(N__58006),
            .I(N__58001));
    Span12Mux_v I__14511 (
            .O(N__58001),
            .I(N__57998));
    Odrv12 I__14510 (
            .O(N__57998),
            .I(ICE_SPI_SCLK));
    InMux I__14509 (
            .O(N__57995),
            .I(N__57992));
    LocalMux I__14508 (
            .O(N__57992),
            .I(N__57989));
    Span4Mux_v I__14507 (
            .O(N__57989),
            .I(N__57986));
    Odrv4 I__14506 (
            .O(N__57986),
            .I(\comm_spi.n14613 ));
    ClkMux I__14505 (
            .O(N__57983),
            .I(N__57443));
    ClkMux I__14504 (
            .O(N__57982),
            .I(N__57443));
    ClkMux I__14503 (
            .O(N__57981),
            .I(N__57443));
    ClkMux I__14502 (
            .O(N__57980),
            .I(N__57443));
    ClkMux I__14501 (
            .O(N__57979),
            .I(N__57443));
    ClkMux I__14500 (
            .O(N__57978),
            .I(N__57443));
    ClkMux I__14499 (
            .O(N__57977),
            .I(N__57443));
    ClkMux I__14498 (
            .O(N__57976),
            .I(N__57443));
    ClkMux I__14497 (
            .O(N__57975),
            .I(N__57443));
    ClkMux I__14496 (
            .O(N__57974),
            .I(N__57443));
    ClkMux I__14495 (
            .O(N__57973),
            .I(N__57443));
    ClkMux I__14494 (
            .O(N__57972),
            .I(N__57443));
    ClkMux I__14493 (
            .O(N__57971),
            .I(N__57443));
    ClkMux I__14492 (
            .O(N__57970),
            .I(N__57443));
    ClkMux I__14491 (
            .O(N__57969),
            .I(N__57443));
    ClkMux I__14490 (
            .O(N__57968),
            .I(N__57443));
    ClkMux I__14489 (
            .O(N__57967),
            .I(N__57443));
    ClkMux I__14488 (
            .O(N__57966),
            .I(N__57443));
    ClkMux I__14487 (
            .O(N__57965),
            .I(N__57443));
    ClkMux I__14486 (
            .O(N__57964),
            .I(N__57443));
    ClkMux I__14485 (
            .O(N__57963),
            .I(N__57443));
    ClkMux I__14484 (
            .O(N__57962),
            .I(N__57443));
    ClkMux I__14483 (
            .O(N__57961),
            .I(N__57443));
    ClkMux I__14482 (
            .O(N__57960),
            .I(N__57443));
    ClkMux I__14481 (
            .O(N__57959),
            .I(N__57443));
    ClkMux I__14480 (
            .O(N__57958),
            .I(N__57443));
    ClkMux I__14479 (
            .O(N__57957),
            .I(N__57443));
    ClkMux I__14478 (
            .O(N__57956),
            .I(N__57443));
    ClkMux I__14477 (
            .O(N__57955),
            .I(N__57443));
    ClkMux I__14476 (
            .O(N__57954),
            .I(N__57443));
    ClkMux I__14475 (
            .O(N__57953),
            .I(N__57443));
    ClkMux I__14474 (
            .O(N__57952),
            .I(N__57443));
    ClkMux I__14473 (
            .O(N__57951),
            .I(N__57443));
    ClkMux I__14472 (
            .O(N__57950),
            .I(N__57443));
    ClkMux I__14471 (
            .O(N__57949),
            .I(N__57443));
    ClkMux I__14470 (
            .O(N__57948),
            .I(N__57443));
    ClkMux I__14469 (
            .O(N__57947),
            .I(N__57443));
    ClkMux I__14468 (
            .O(N__57946),
            .I(N__57443));
    ClkMux I__14467 (
            .O(N__57945),
            .I(N__57443));
    ClkMux I__14466 (
            .O(N__57944),
            .I(N__57443));
    ClkMux I__14465 (
            .O(N__57943),
            .I(N__57443));
    ClkMux I__14464 (
            .O(N__57942),
            .I(N__57443));
    ClkMux I__14463 (
            .O(N__57941),
            .I(N__57443));
    ClkMux I__14462 (
            .O(N__57940),
            .I(N__57443));
    ClkMux I__14461 (
            .O(N__57939),
            .I(N__57443));
    ClkMux I__14460 (
            .O(N__57938),
            .I(N__57443));
    ClkMux I__14459 (
            .O(N__57937),
            .I(N__57443));
    ClkMux I__14458 (
            .O(N__57936),
            .I(N__57443));
    ClkMux I__14457 (
            .O(N__57935),
            .I(N__57443));
    ClkMux I__14456 (
            .O(N__57934),
            .I(N__57443));
    ClkMux I__14455 (
            .O(N__57933),
            .I(N__57443));
    ClkMux I__14454 (
            .O(N__57932),
            .I(N__57443));
    ClkMux I__14453 (
            .O(N__57931),
            .I(N__57443));
    ClkMux I__14452 (
            .O(N__57930),
            .I(N__57443));
    ClkMux I__14451 (
            .O(N__57929),
            .I(N__57443));
    ClkMux I__14450 (
            .O(N__57928),
            .I(N__57443));
    ClkMux I__14449 (
            .O(N__57927),
            .I(N__57443));
    ClkMux I__14448 (
            .O(N__57926),
            .I(N__57443));
    ClkMux I__14447 (
            .O(N__57925),
            .I(N__57443));
    ClkMux I__14446 (
            .O(N__57924),
            .I(N__57443));
    ClkMux I__14445 (
            .O(N__57923),
            .I(N__57443));
    ClkMux I__14444 (
            .O(N__57922),
            .I(N__57443));
    ClkMux I__14443 (
            .O(N__57921),
            .I(N__57443));
    ClkMux I__14442 (
            .O(N__57920),
            .I(N__57443));
    ClkMux I__14441 (
            .O(N__57919),
            .I(N__57443));
    ClkMux I__14440 (
            .O(N__57918),
            .I(N__57443));
    ClkMux I__14439 (
            .O(N__57917),
            .I(N__57443));
    ClkMux I__14438 (
            .O(N__57916),
            .I(N__57443));
    ClkMux I__14437 (
            .O(N__57915),
            .I(N__57443));
    ClkMux I__14436 (
            .O(N__57914),
            .I(N__57443));
    ClkMux I__14435 (
            .O(N__57913),
            .I(N__57443));
    ClkMux I__14434 (
            .O(N__57912),
            .I(N__57443));
    ClkMux I__14433 (
            .O(N__57911),
            .I(N__57443));
    ClkMux I__14432 (
            .O(N__57910),
            .I(N__57443));
    ClkMux I__14431 (
            .O(N__57909),
            .I(N__57443));
    ClkMux I__14430 (
            .O(N__57908),
            .I(N__57443));
    ClkMux I__14429 (
            .O(N__57907),
            .I(N__57443));
    ClkMux I__14428 (
            .O(N__57906),
            .I(N__57443));
    ClkMux I__14427 (
            .O(N__57905),
            .I(N__57443));
    ClkMux I__14426 (
            .O(N__57904),
            .I(N__57443));
    ClkMux I__14425 (
            .O(N__57903),
            .I(N__57443));
    ClkMux I__14424 (
            .O(N__57902),
            .I(N__57443));
    ClkMux I__14423 (
            .O(N__57901),
            .I(N__57443));
    ClkMux I__14422 (
            .O(N__57900),
            .I(N__57443));
    ClkMux I__14421 (
            .O(N__57899),
            .I(N__57443));
    ClkMux I__14420 (
            .O(N__57898),
            .I(N__57443));
    ClkMux I__14419 (
            .O(N__57897),
            .I(N__57443));
    ClkMux I__14418 (
            .O(N__57896),
            .I(N__57443));
    ClkMux I__14417 (
            .O(N__57895),
            .I(N__57443));
    ClkMux I__14416 (
            .O(N__57894),
            .I(N__57443));
    ClkMux I__14415 (
            .O(N__57893),
            .I(N__57443));
    ClkMux I__14414 (
            .O(N__57892),
            .I(N__57443));
    ClkMux I__14413 (
            .O(N__57891),
            .I(N__57443));
    ClkMux I__14412 (
            .O(N__57890),
            .I(N__57443));
    ClkMux I__14411 (
            .O(N__57889),
            .I(N__57443));
    ClkMux I__14410 (
            .O(N__57888),
            .I(N__57443));
    ClkMux I__14409 (
            .O(N__57887),
            .I(N__57443));
    ClkMux I__14408 (
            .O(N__57886),
            .I(N__57443));
    ClkMux I__14407 (
            .O(N__57885),
            .I(N__57443));
    ClkMux I__14406 (
            .O(N__57884),
            .I(N__57443));
    ClkMux I__14405 (
            .O(N__57883),
            .I(N__57443));
    ClkMux I__14404 (
            .O(N__57882),
            .I(N__57443));
    ClkMux I__14403 (
            .O(N__57881),
            .I(N__57443));
    ClkMux I__14402 (
            .O(N__57880),
            .I(N__57443));
    ClkMux I__14401 (
            .O(N__57879),
            .I(N__57443));
    ClkMux I__14400 (
            .O(N__57878),
            .I(N__57443));
    ClkMux I__14399 (
            .O(N__57877),
            .I(N__57443));
    ClkMux I__14398 (
            .O(N__57876),
            .I(N__57443));
    ClkMux I__14397 (
            .O(N__57875),
            .I(N__57443));
    ClkMux I__14396 (
            .O(N__57874),
            .I(N__57443));
    ClkMux I__14395 (
            .O(N__57873),
            .I(N__57443));
    ClkMux I__14394 (
            .O(N__57872),
            .I(N__57443));
    ClkMux I__14393 (
            .O(N__57871),
            .I(N__57443));
    ClkMux I__14392 (
            .O(N__57870),
            .I(N__57443));
    ClkMux I__14391 (
            .O(N__57869),
            .I(N__57443));
    ClkMux I__14390 (
            .O(N__57868),
            .I(N__57443));
    ClkMux I__14389 (
            .O(N__57867),
            .I(N__57443));
    ClkMux I__14388 (
            .O(N__57866),
            .I(N__57443));
    ClkMux I__14387 (
            .O(N__57865),
            .I(N__57443));
    ClkMux I__14386 (
            .O(N__57864),
            .I(N__57443));
    ClkMux I__14385 (
            .O(N__57863),
            .I(N__57443));
    ClkMux I__14384 (
            .O(N__57862),
            .I(N__57443));
    ClkMux I__14383 (
            .O(N__57861),
            .I(N__57443));
    ClkMux I__14382 (
            .O(N__57860),
            .I(N__57443));
    ClkMux I__14381 (
            .O(N__57859),
            .I(N__57443));
    ClkMux I__14380 (
            .O(N__57858),
            .I(N__57443));
    ClkMux I__14379 (
            .O(N__57857),
            .I(N__57443));
    ClkMux I__14378 (
            .O(N__57856),
            .I(N__57443));
    ClkMux I__14377 (
            .O(N__57855),
            .I(N__57443));
    ClkMux I__14376 (
            .O(N__57854),
            .I(N__57443));
    ClkMux I__14375 (
            .O(N__57853),
            .I(N__57443));
    ClkMux I__14374 (
            .O(N__57852),
            .I(N__57443));
    ClkMux I__14373 (
            .O(N__57851),
            .I(N__57443));
    ClkMux I__14372 (
            .O(N__57850),
            .I(N__57443));
    ClkMux I__14371 (
            .O(N__57849),
            .I(N__57443));
    ClkMux I__14370 (
            .O(N__57848),
            .I(N__57443));
    ClkMux I__14369 (
            .O(N__57847),
            .I(N__57443));
    ClkMux I__14368 (
            .O(N__57846),
            .I(N__57443));
    ClkMux I__14367 (
            .O(N__57845),
            .I(N__57443));
    ClkMux I__14366 (
            .O(N__57844),
            .I(N__57443));
    ClkMux I__14365 (
            .O(N__57843),
            .I(N__57443));
    ClkMux I__14364 (
            .O(N__57842),
            .I(N__57443));
    ClkMux I__14363 (
            .O(N__57841),
            .I(N__57443));
    ClkMux I__14362 (
            .O(N__57840),
            .I(N__57443));
    ClkMux I__14361 (
            .O(N__57839),
            .I(N__57443));
    ClkMux I__14360 (
            .O(N__57838),
            .I(N__57443));
    ClkMux I__14359 (
            .O(N__57837),
            .I(N__57443));
    ClkMux I__14358 (
            .O(N__57836),
            .I(N__57443));
    ClkMux I__14357 (
            .O(N__57835),
            .I(N__57443));
    ClkMux I__14356 (
            .O(N__57834),
            .I(N__57443));
    ClkMux I__14355 (
            .O(N__57833),
            .I(N__57443));
    ClkMux I__14354 (
            .O(N__57832),
            .I(N__57443));
    ClkMux I__14353 (
            .O(N__57831),
            .I(N__57443));
    ClkMux I__14352 (
            .O(N__57830),
            .I(N__57443));
    ClkMux I__14351 (
            .O(N__57829),
            .I(N__57443));
    ClkMux I__14350 (
            .O(N__57828),
            .I(N__57443));
    ClkMux I__14349 (
            .O(N__57827),
            .I(N__57443));
    ClkMux I__14348 (
            .O(N__57826),
            .I(N__57443));
    ClkMux I__14347 (
            .O(N__57825),
            .I(N__57443));
    ClkMux I__14346 (
            .O(N__57824),
            .I(N__57443));
    ClkMux I__14345 (
            .O(N__57823),
            .I(N__57443));
    ClkMux I__14344 (
            .O(N__57822),
            .I(N__57443));
    ClkMux I__14343 (
            .O(N__57821),
            .I(N__57443));
    ClkMux I__14342 (
            .O(N__57820),
            .I(N__57443));
    ClkMux I__14341 (
            .O(N__57819),
            .I(N__57443));
    ClkMux I__14340 (
            .O(N__57818),
            .I(N__57443));
    ClkMux I__14339 (
            .O(N__57817),
            .I(N__57443));
    ClkMux I__14338 (
            .O(N__57816),
            .I(N__57443));
    ClkMux I__14337 (
            .O(N__57815),
            .I(N__57443));
    ClkMux I__14336 (
            .O(N__57814),
            .I(N__57443));
    ClkMux I__14335 (
            .O(N__57813),
            .I(N__57443));
    ClkMux I__14334 (
            .O(N__57812),
            .I(N__57443));
    ClkMux I__14333 (
            .O(N__57811),
            .I(N__57443));
    ClkMux I__14332 (
            .O(N__57810),
            .I(N__57443));
    ClkMux I__14331 (
            .O(N__57809),
            .I(N__57443));
    ClkMux I__14330 (
            .O(N__57808),
            .I(N__57443));
    ClkMux I__14329 (
            .O(N__57807),
            .I(N__57443));
    ClkMux I__14328 (
            .O(N__57806),
            .I(N__57443));
    ClkMux I__14327 (
            .O(N__57805),
            .I(N__57443));
    ClkMux I__14326 (
            .O(N__57804),
            .I(N__57443));
    GlobalMux I__14325 (
            .O(N__57443),
            .I(clk_32MHz));
    SRMux I__14324 (
            .O(N__57440),
            .I(N__57437));
    LocalMux I__14323 (
            .O(N__57437),
            .I(N__57434));
    Span4Mux_h I__14322 (
            .O(N__57434),
            .I(N__57431));
    Span4Mux_v I__14321 (
            .O(N__57431),
            .I(N__57428));
    Odrv4 I__14320 (
            .O(N__57428),
            .I(\comm_spi.iclk_N_764 ));
    CascadeMux I__14319 (
            .O(N__57425),
            .I(N__57419));
    CascadeMux I__14318 (
            .O(N__57424),
            .I(N__57415));
    CascadeMux I__14317 (
            .O(N__57423),
            .I(N__57411));
    InMux I__14316 (
            .O(N__57422),
            .I(N__57395));
    InMux I__14315 (
            .O(N__57419),
            .I(N__57395));
    InMux I__14314 (
            .O(N__57418),
            .I(N__57395));
    InMux I__14313 (
            .O(N__57415),
            .I(N__57395));
    InMux I__14312 (
            .O(N__57414),
            .I(N__57395));
    InMux I__14311 (
            .O(N__57411),
            .I(N__57395));
    InMux I__14310 (
            .O(N__57410),
            .I(N__57395));
    LocalMux I__14309 (
            .O(N__57395),
            .I(N__57385));
    CascadeMux I__14308 (
            .O(N__57394),
            .I(N__57376));
    CascadeMux I__14307 (
            .O(N__57393),
            .I(N__57370));
    CascadeMux I__14306 (
            .O(N__57392),
            .I(N__57366));
    CascadeMux I__14305 (
            .O(N__57391),
            .I(N__57362));
    CascadeMux I__14304 (
            .O(N__57390),
            .I(N__57358));
    CascadeMux I__14303 (
            .O(N__57389),
            .I(N__57354));
    CascadeMux I__14302 (
            .O(N__57388),
            .I(N__57350));
    Span4Mux_v I__14301 (
            .O(N__57385),
            .I(N__57347));
    CascadeMux I__14300 (
            .O(N__57384),
            .I(N__57343));
    CascadeMux I__14299 (
            .O(N__57383),
            .I(N__57339));
    CascadeMux I__14298 (
            .O(N__57382),
            .I(N__57335));
    CascadeMux I__14297 (
            .O(N__57381),
            .I(N__57331));
    SRMux I__14296 (
            .O(N__57380),
            .I(N__57328));
    SRMux I__14295 (
            .O(N__57379),
            .I(N__57321));
    InMux I__14294 (
            .O(N__57376),
            .I(N__57301));
    InMux I__14293 (
            .O(N__57375),
            .I(N__57301));
    InMux I__14292 (
            .O(N__57374),
            .I(N__57301));
    InMux I__14291 (
            .O(N__57373),
            .I(N__57301));
    InMux I__14290 (
            .O(N__57370),
            .I(N__57301));
    InMux I__14289 (
            .O(N__57369),
            .I(N__57301));
    InMux I__14288 (
            .O(N__57366),
            .I(N__57301));
    InMux I__14287 (
            .O(N__57365),
            .I(N__57301));
    InMux I__14286 (
            .O(N__57362),
            .I(N__57286));
    InMux I__14285 (
            .O(N__57361),
            .I(N__57286));
    InMux I__14284 (
            .O(N__57358),
            .I(N__57286));
    InMux I__14283 (
            .O(N__57357),
            .I(N__57286));
    InMux I__14282 (
            .O(N__57354),
            .I(N__57286));
    InMux I__14281 (
            .O(N__57353),
            .I(N__57286));
    InMux I__14280 (
            .O(N__57350),
            .I(N__57286));
    Span4Mux_v I__14279 (
            .O(N__57347),
            .I(N__57283));
    InMux I__14278 (
            .O(N__57346),
            .I(N__57266));
    InMux I__14277 (
            .O(N__57343),
            .I(N__57266));
    InMux I__14276 (
            .O(N__57342),
            .I(N__57266));
    InMux I__14275 (
            .O(N__57339),
            .I(N__57266));
    InMux I__14274 (
            .O(N__57338),
            .I(N__57266));
    InMux I__14273 (
            .O(N__57335),
            .I(N__57266));
    InMux I__14272 (
            .O(N__57334),
            .I(N__57266));
    InMux I__14271 (
            .O(N__57331),
            .I(N__57266));
    LocalMux I__14270 (
            .O(N__57328),
            .I(N__57263));
    CascadeMux I__14269 (
            .O(N__57327),
            .I(N__57260));
    CascadeMux I__14268 (
            .O(N__57326),
            .I(N__57256));
    CascadeMux I__14267 (
            .O(N__57325),
            .I(N__57252));
    CascadeMux I__14266 (
            .O(N__57324),
            .I(N__57248));
    LocalMux I__14265 (
            .O(N__57321),
            .I(N__57245));
    SRMux I__14264 (
            .O(N__57320),
            .I(N__57242));
    SRMux I__14263 (
            .O(N__57319),
            .I(N__57239));
    SRMux I__14262 (
            .O(N__57318),
            .I(N__57233));
    LocalMux I__14261 (
            .O(N__57301),
            .I(N__57227));
    LocalMux I__14260 (
            .O(N__57286),
            .I(N__57227));
    Span4Mux_v I__14259 (
            .O(N__57283),
            .I(N__57222));
    LocalMux I__14258 (
            .O(N__57266),
            .I(N__57222));
    Span4Mux_h I__14257 (
            .O(N__57263),
            .I(N__57219));
    InMux I__14256 (
            .O(N__57260),
            .I(N__57204));
    InMux I__14255 (
            .O(N__57259),
            .I(N__57204));
    InMux I__14254 (
            .O(N__57256),
            .I(N__57204));
    InMux I__14253 (
            .O(N__57255),
            .I(N__57204));
    InMux I__14252 (
            .O(N__57252),
            .I(N__57204));
    InMux I__14251 (
            .O(N__57251),
            .I(N__57204));
    InMux I__14250 (
            .O(N__57248),
            .I(N__57204));
    Span4Mux_v I__14249 (
            .O(N__57245),
            .I(N__57197));
    LocalMux I__14248 (
            .O(N__57242),
            .I(N__57197));
    LocalMux I__14247 (
            .O(N__57239),
            .I(N__57197));
    SRMux I__14246 (
            .O(N__57238),
            .I(N__57194));
    InMux I__14245 (
            .O(N__57237),
            .I(N__57191));
    SRMux I__14244 (
            .O(N__57236),
            .I(N__57188));
    LocalMux I__14243 (
            .O(N__57233),
            .I(N__57182));
    IoInMux I__14242 (
            .O(N__57232),
            .I(N__57179));
    Span4Mux_v I__14241 (
            .O(N__57227),
            .I(N__57174));
    Span4Mux_v I__14240 (
            .O(N__57222),
            .I(N__57174));
    Span4Mux_h I__14239 (
            .O(N__57219),
            .I(N__57171));
    LocalMux I__14238 (
            .O(N__57204),
            .I(N__57168));
    Span4Mux_v I__14237 (
            .O(N__57197),
            .I(N__57158));
    LocalMux I__14236 (
            .O(N__57194),
            .I(N__57158));
    LocalMux I__14235 (
            .O(N__57191),
            .I(N__57158));
    LocalMux I__14234 (
            .O(N__57188),
            .I(N__57158));
    SRMux I__14233 (
            .O(N__57187),
            .I(N__57155));
    InMux I__14232 (
            .O(N__57186),
            .I(N__57152));
    SRMux I__14231 (
            .O(N__57185),
            .I(N__57149));
    Span12Mux_h I__14230 (
            .O(N__57182),
            .I(N__57144));
    LocalMux I__14229 (
            .O(N__57179),
            .I(N__57141));
    Span4Mux_h I__14228 (
            .O(N__57174),
            .I(N__57138));
    Span4Mux_h I__14227 (
            .O(N__57171),
            .I(N__57133));
    Span4Mux_h I__14226 (
            .O(N__57168),
            .I(N__57133));
    SRMux I__14225 (
            .O(N__57167),
            .I(N__57130));
    Span4Mux_v I__14224 (
            .O(N__57158),
            .I(N__57121));
    LocalMux I__14223 (
            .O(N__57155),
            .I(N__57121));
    LocalMux I__14222 (
            .O(N__57152),
            .I(N__57121));
    LocalMux I__14221 (
            .O(N__57149),
            .I(N__57121));
    SRMux I__14220 (
            .O(N__57148),
            .I(N__57118));
    SRMux I__14219 (
            .O(N__57147),
            .I(N__57115));
    Span12Mux_h I__14218 (
            .O(N__57144),
            .I(N__57112));
    Span12Mux_s8_v I__14217 (
            .O(N__57141),
            .I(N__57109));
    Span4Mux_h I__14216 (
            .O(N__57138),
            .I(N__57106));
    Span4Mux_h I__14215 (
            .O(N__57133),
            .I(N__57103));
    LocalMux I__14214 (
            .O(N__57130),
            .I(N__57100));
    Span4Mux_v I__14213 (
            .O(N__57121),
            .I(N__57093));
    LocalMux I__14212 (
            .O(N__57118),
            .I(N__57093));
    LocalMux I__14211 (
            .O(N__57115),
            .I(N__57093));
    Odrv12 I__14210 (
            .O(N__57112),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__14209 (
            .O(N__57109),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__14208 (
            .O(N__57106),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__14207 (
            .O(N__57103),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__14206 (
            .O(N__57100),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__14205 (
            .O(N__57093),
            .I(CONSTANT_ONE_NET));
    InMux I__14204 (
            .O(N__57080),
            .I(N__57076));
    InMux I__14203 (
            .O(N__57079),
            .I(N__57073));
    LocalMux I__14202 (
            .O(N__57076),
            .I(N__57070));
    LocalMux I__14201 (
            .O(N__57073),
            .I(N__57067));
    Odrv12 I__14200 (
            .O(N__57070),
            .I(\comm_spi.n14609 ));
    Odrv4 I__14199 (
            .O(N__57067),
            .I(\comm_spi.n14609 ));
    ClkMux I__14198 (
            .O(N__57062),
            .I(N__57059));
    LocalMux I__14197 (
            .O(N__57059),
            .I(N__57055));
    ClkMux I__14196 (
            .O(N__57058),
            .I(N__57052));
    Span4Mux_h I__14195 (
            .O(N__57055),
            .I(N__57044));
    LocalMux I__14194 (
            .O(N__57052),
            .I(N__57044));
    ClkMux I__14193 (
            .O(N__57051),
            .I(N__57041));
    ClkMux I__14192 (
            .O(N__57050),
            .I(N__57037));
    ClkMux I__14191 (
            .O(N__57049),
            .I(N__57032));
    Span4Mux_v I__14190 (
            .O(N__57044),
            .I(N__57027));
    LocalMux I__14189 (
            .O(N__57041),
            .I(N__57027));
    ClkMux I__14188 (
            .O(N__57040),
            .I(N__57024));
    LocalMux I__14187 (
            .O(N__57037),
            .I(N__57021));
    ClkMux I__14186 (
            .O(N__57036),
            .I(N__57018));
    ClkMux I__14185 (
            .O(N__57035),
            .I(N__57013));
    LocalMux I__14184 (
            .O(N__57032),
            .I(N__57009));
    Span4Mux_h I__14183 (
            .O(N__57027),
            .I(N__57004));
    LocalMux I__14182 (
            .O(N__57024),
            .I(N__57004));
    Span4Mux_v I__14181 (
            .O(N__57021),
            .I(N__56999));
    LocalMux I__14180 (
            .O(N__57018),
            .I(N__56999));
    ClkMux I__14179 (
            .O(N__57017),
            .I(N__56992));
    ClkMux I__14178 (
            .O(N__57016),
            .I(N__56988));
    LocalMux I__14177 (
            .O(N__57013),
            .I(N__56984));
    ClkMux I__14176 (
            .O(N__57012),
            .I(N__56980));
    Span4Mux_v I__14175 (
            .O(N__57009),
            .I(N__56975));
    Span4Mux_v I__14174 (
            .O(N__57004),
            .I(N__56975));
    Span4Mux_h I__14173 (
            .O(N__56999),
            .I(N__56972));
    ClkMux I__14172 (
            .O(N__56998),
            .I(N__56969));
    ClkMux I__14171 (
            .O(N__56997),
            .I(N__56966));
    ClkMux I__14170 (
            .O(N__56996),
            .I(N__56963));
    ClkMux I__14169 (
            .O(N__56995),
            .I(N__56960));
    LocalMux I__14168 (
            .O(N__56992),
            .I(N__56957));
    ClkMux I__14167 (
            .O(N__56991),
            .I(N__56954));
    LocalMux I__14166 (
            .O(N__56988),
            .I(N__56951));
    ClkMux I__14165 (
            .O(N__56987),
            .I(N__56948));
    Span4Mux_v I__14164 (
            .O(N__56984),
            .I(N__56945));
    ClkMux I__14163 (
            .O(N__56983),
            .I(N__56942));
    LocalMux I__14162 (
            .O(N__56980),
            .I(N__56939));
    Span4Mux_h I__14161 (
            .O(N__56975),
            .I(N__56936));
    Span4Mux_v I__14160 (
            .O(N__56972),
            .I(N__56931));
    LocalMux I__14159 (
            .O(N__56969),
            .I(N__56931));
    LocalMux I__14158 (
            .O(N__56966),
            .I(N__56926));
    LocalMux I__14157 (
            .O(N__56963),
            .I(N__56926));
    LocalMux I__14156 (
            .O(N__56960),
            .I(N__56919));
    Span4Mux_h I__14155 (
            .O(N__56957),
            .I(N__56919));
    LocalMux I__14154 (
            .O(N__56954),
            .I(N__56919));
    Span4Mux_h I__14153 (
            .O(N__56951),
            .I(N__56912));
    LocalMux I__14152 (
            .O(N__56948),
            .I(N__56912));
    Span4Mux_h I__14151 (
            .O(N__56945),
            .I(N__56907));
    LocalMux I__14150 (
            .O(N__56942),
            .I(N__56904));
    Span4Mux_v I__14149 (
            .O(N__56939),
            .I(N__56899));
    Span4Mux_v I__14148 (
            .O(N__56936),
            .I(N__56899));
    Span4Mux_v I__14147 (
            .O(N__56931),
            .I(N__56892));
    Span4Mux_v I__14146 (
            .O(N__56926),
            .I(N__56892));
    Span4Mux_v I__14145 (
            .O(N__56919),
            .I(N__56892));
    ClkMux I__14144 (
            .O(N__56918),
            .I(N__56889));
    ClkMux I__14143 (
            .O(N__56917),
            .I(N__56886));
    Span4Mux_v I__14142 (
            .O(N__56912),
            .I(N__56883));
    ClkMux I__14141 (
            .O(N__56911),
            .I(N__56880));
    ClkMux I__14140 (
            .O(N__56910),
            .I(N__56877));
    Odrv4 I__14139 (
            .O(N__56907),
            .I(\comm_spi.iclk ));
    Odrv12 I__14138 (
            .O(N__56904),
            .I(\comm_spi.iclk ));
    Odrv4 I__14137 (
            .O(N__56899),
            .I(\comm_spi.iclk ));
    Odrv4 I__14136 (
            .O(N__56892),
            .I(\comm_spi.iclk ));
    LocalMux I__14135 (
            .O(N__56889),
            .I(\comm_spi.iclk ));
    LocalMux I__14134 (
            .O(N__56886),
            .I(\comm_spi.iclk ));
    Odrv4 I__14133 (
            .O(N__56883),
            .I(\comm_spi.iclk ));
    LocalMux I__14132 (
            .O(N__56880),
            .I(\comm_spi.iclk ));
    LocalMux I__14131 (
            .O(N__56877),
            .I(\comm_spi.iclk ));
    SRMux I__14130 (
            .O(N__56858),
            .I(N__56855));
    LocalMux I__14129 (
            .O(N__56855),
            .I(N__56849));
    SRMux I__14128 (
            .O(N__56854),
            .I(N__56846));
    CascadeMux I__14127 (
            .O(N__56853),
            .I(N__56838));
    InMux I__14126 (
            .O(N__56852),
            .I(N__56829));
    Span4Mux_v I__14125 (
            .O(N__56849),
            .I(N__56824));
    LocalMux I__14124 (
            .O(N__56846),
            .I(N__56824));
    InMux I__14123 (
            .O(N__56845),
            .I(N__56818));
    InMux I__14122 (
            .O(N__56844),
            .I(N__56818));
    InMux I__14121 (
            .O(N__56843),
            .I(N__56811));
    InMux I__14120 (
            .O(N__56842),
            .I(N__56811));
    InMux I__14119 (
            .O(N__56841),
            .I(N__56804));
    InMux I__14118 (
            .O(N__56838),
            .I(N__56795));
    InMux I__14117 (
            .O(N__56837),
            .I(N__56795));
    InMux I__14116 (
            .O(N__56836),
            .I(N__56795));
    InMux I__14115 (
            .O(N__56835),
            .I(N__56795));
    InMux I__14114 (
            .O(N__56834),
            .I(N__56792));
    InMux I__14113 (
            .O(N__56833),
            .I(N__56787));
    InMux I__14112 (
            .O(N__56832),
            .I(N__56787));
    LocalMux I__14111 (
            .O(N__56829),
            .I(N__56784));
    Span4Mux_v I__14110 (
            .O(N__56824),
            .I(N__56781));
    SRMux I__14109 (
            .O(N__56823),
            .I(N__56778));
    LocalMux I__14108 (
            .O(N__56818),
            .I(N__56772));
    InMux I__14107 (
            .O(N__56817),
            .I(N__56767));
    InMux I__14106 (
            .O(N__56816),
            .I(N__56767));
    LocalMux I__14105 (
            .O(N__56811),
            .I(N__56764));
    InMux I__14104 (
            .O(N__56810),
            .I(N__56761));
    InMux I__14103 (
            .O(N__56809),
            .I(N__56755));
    InMux I__14102 (
            .O(N__56808),
            .I(N__56755));
    InMux I__14101 (
            .O(N__56807),
            .I(N__56752));
    LocalMux I__14100 (
            .O(N__56804),
            .I(N__56737));
    LocalMux I__14099 (
            .O(N__56795),
            .I(N__56737));
    LocalMux I__14098 (
            .O(N__56792),
            .I(N__56732));
    LocalMux I__14097 (
            .O(N__56787),
            .I(N__56732));
    Span4Mux_v I__14096 (
            .O(N__56784),
            .I(N__56727));
    Span4Mux_v I__14095 (
            .O(N__56781),
            .I(N__56727));
    LocalMux I__14094 (
            .O(N__56778),
            .I(N__56724));
    InMux I__14093 (
            .O(N__56777),
            .I(N__56719));
    InMux I__14092 (
            .O(N__56776),
            .I(N__56719));
    InMux I__14091 (
            .O(N__56775),
            .I(N__56716));
    Span4Mux_h I__14090 (
            .O(N__56772),
            .I(N__56713));
    LocalMux I__14089 (
            .O(N__56767),
            .I(N__56706));
    Span4Mux_v I__14088 (
            .O(N__56764),
            .I(N__56706));
    LocalMux I__14087 (
            .O(N__56761),
            .I(N__56706));
    InMux I__14086 (
            .O(N__56760),
            .I(N__56703));
    LocalMux I__14085 (
            .O(N__56755),
            .I(N__56698));
    LocalMux I__14084 (
            .O(N__56752),
            .I(N__56698));
    InMux I__14083 (
            .O(N__56751),
            .I(N__56695));
    InMux I__14082 (
            .O(N__56750),
            .I(N__56684));
    InMux I__14081 (
            .O(N__56749),
            .I(N__56684));
    InMux I__14080 (
            .O(N__56748),
            .I(N__56684));
    InMux I__14079 (
            .O(N__56747),
            .I(N__56684));
    InMux I__14078 (
            .O(N__56746),
            .I(N__56684));
    InMux I__14077 (
            .O(N__56745),
            .I(N__56675));
    InMux I__14076 (
            .O(N__56744),
            .I(N__56675));
    InMux I__14075 (
            .O(N__56743),
            .I(N__56675));
    InMux I__14074 (
            .O(N__56742),
            .I(N__56675));
    Span4Mux_v I__14073 (
            .O(N__56737),
            .I(N__56672));
    Span4Mux_h I__14072 (
            .O(N__56732),
            .I(N__56667));
    Span4Mux_h I__14071 (
            .O(N__56727),
            .I(N__56667));
    Span12Mux_h I__14070 (
            .O(N__56724),
            .I(N__56662));
    LocalMux I__14069 (
            .O(N__56719),
            .I(N__56662));
    LocalMux I__14068 (
            .O(N__56716),
            .I(N__56655));
    Span4Mux_v I__14067 (
            .O(N__56713),
            .I(N__56655));
    Span4Mux_h I__14066 (
            .O(N__56706),
            .I(N__56655));
    LocalMux I__14065 (
            .O(N__56703),
            .I(N__56650));
    Span4Mux_v I__14064 (
            .O(N__56698),
            .I(N__56650));
    LocalMux I__14063 (
            .O(N__56695),
            .I(comm_clear));
    LocalMux I__14062 (
            .O(N__56684),
            .I(comm_clear));
    LocalMux I__14061 (
            .O(N__56675),
            .I(comm_clear));
    Odrv4 I__14060 (
            .O(N__56672),
            .I(comm_clear));
    Odrv4 I__14059 (
            .O(N__56667),
            .I(comm_clear));
    Odrv12 I__14058 (
            .O(N__56662),
            .I(comm_clear));
    Odrv4 I__14057 (
            .O(N__56655),
            .I(comm_clear));
    Odrv4 I__14056 (
            .O(N__56650),
            .I(comm_clear));
    InMux I__14055 (
            .O(N__56633),
            .I(N__56629));
    InMux I__14054 (
            .O(N__56632),
            .I(N__56625));
    LocalMux I__14053 (
            .O(N__56629),
            .I(N__56622));
    InMux I__14052 (
            .O(N__56628),
            .I(N__56619));
    LocalMux I__14051 (
            .O(N__56625),
            .I(N__56616));
    Span4Mux_v I__14050 (
            .O(N__56622),
            .I(N__56611));
    LocalMux I__14049 (
            .O(N__56619),
            .I(N__56611));
    Sp12to4 I__14048 (
            .O(N__56616),
            .I(N__56608));
    Span4Mux_v I__14047 (
            .O(N__56611),
            .I(N__56605));
    Span12Mux_v I__14046 (
            .O(N__56608),
            .I(N__56600));
    Sp12to4 I__14045 (
            .O(N__56605),
            .I(N__56600));
    Odrv12 I__14044 (
            .O(N__56600),
            .I(comm_tx_buf_0));
    SRMux I__14043 (
            .O(N__56597),
            .I(N__56594));
    LocalMux I__14042 (
            .O(N__56594),
            .I(N__56591));
    Span4Mux_h I__14041 (
            .O(N__56591),
            .I(N__56588));
    Odrv4 I__14040 (
            .O(N__56588),
            .I(\comm_spi.data_tx_7__N_796 ));
    InMux I__14039 (
            .O(N__56585),
            .I(N__56581));
    InMux I__14038 (
            .O(N__56584),
            .I(N__56578));
    LocalMux I__14037 (
            .O(N__56581),
            .I(N__56572));
    LocalMux I__14036 (
            .O(N__56578),
            .I(N__56572));
    InMux I__14035 (
            .O(N__56577),
            .I(N__56569));
    Odrv4 I__14034 (
            .O(N__56572),
            .I(\comm_spi.n22661 ));
    LocalMux I__14033 (
            .O(N__56569),
            .I(\comm_spi.n22661 ));
    InMux I__14032 (
            .O(N__56564),
            .I(N__56560));
    InMux I__14031 (
            .O(N__56563),
            .I(N__56557));
    LocalMux I__14030 (
            .O(N__56560),
            .I(N__56554));
    LocalMux I__14029 (
            .O(N__56557),
            .I(\comm_spi.n14623 ));
    Odrv4 I__14028 (
            .O(N__56554),
            .I(\comm_spi.n14623 ));
    SRMux I__14027 (
            .O(N__56549),
            .I(N__56546));
    LocalMux I__14026 (
            .O(N__56546),
            .I(N__56543));
    Span4Mux_v I__14025 (
            .O(N__56543),
            .I(N__56539));
    SRMux I__14024 (
            .O(N__56542),
            .I(N__56536));
    Span4Mux_v I__14023 (
            .O(N__56539),
            .I(N__56530));
    LocalMux I__14022 (
            .O(N__56536),
            .I(N__56530));
    SRMux I__14021 (
            .O(N__56535),
            .I(N__56527));
    Span4Mux_h I__14020 (
            .O(N__56530),
            .I(N__56524));
    LocalMux I__14019 (
            .O(N__56527),
            .I(N__56521));
    Span4Mux_v I__14018 (
            .O(N__56524),
            .I(N__56516));
    Span4Mux_v I__14017 (
            .O(N__56521),
            .I(N__56516));
    Odrv4 I__14016 (
            .O(N__56516),
            .I(\comm_spi.data_tx_7__N_767 ));
    InMux I__14015 (
            .O(N__56513),
            .I(N__56510));
    LocalMux I__14014 (
            .O(N__56510),
            .I(N__56507));
    Span4Mux_h I__14013 (
            .O(N__56507),
            .I(N__56502));
    InMux I__14012 (
            .O(N__56506),
            .I(N__56499));
    InMux I__14011 (
            .O(N__56505),
            .I(N__56496));
    Odrv4 I__14010 (
            .O(N__56502),
            .I(comm_tx_buf_7));
    LocalMux I__14009 (
            .O(N__56499),
            .I(comm_tx_buf_7));
    LocalMux I__14008 (
            .O(N__56496),
            .I(comm_tx_buf_7));
    SRMux I__14007 (
            .O(N__56489),
            .I(N__56484));
    SRMux I__14006 (
            .O(N__56488),
            .I(N__56481));
    SRMux I__14005 (
            .O(N__56487),
            .I(N__56478));
    LocalMux I__14004 (
            .O(N__56484),
            .I(N__56475));
    LocalMux I__14003 (
            .O(N__56481),
            .I(N__56470));
    LocalMux I__14002 (
            .O(N__56478),
            .I(N__56470));
    Span4Mux_v I__14001 (
            .O(N__56475),
            .I(N__56467));
    Span4Mux_v I__14000 (
            .O(N__56470),
            .I(N__56464));
    Odrv4 I__13999 (
            .O(N__56467),
            .I(\comm_spi.data_tx_7__N_775 ));
    Odrv4 I__13998 (
            .O(N__56464),
            .I(\comm_spi.data_tx_7__N_775 ));
    InMux I__13997 (
            .O(N__56459),
            .I(N__56456));
    LocalMux I__13996 (
            .O(N__56456),
            .I(N__56452));
    InMux I__13995 (
            .O(N__56455),
            .I(N__56449));
    Odrv4 I__13994 (
            .O(N__56452),
            .I(\comm_spi.n14635 ));
    LocalMux I__13993 (
            .O(N__56449),
            .I(\comm_spi.n14635 ));
    SRMux I__13992 (
            .O(N__56444),
            .I(N__56441));
    LocalMux I__13991 (
            .O(N__56441),
            .I(N__56438));
    Span4Mux_v I__13990 (
            .O(N__56438),
            .I(N__56435));
    Odrv4 I__13989 (
            .O(N__56435),
            .I(\comm_spi.data_tx_7__N_793 ));
    InMux I__13988 (
            .O(N__56432),
            .I(N__56429));
    LocalMux I__13987 (
            .O(N__56429),
            .I(N__56426));
    Span4Mux_h I__13986 (
            .O(N__56426),
            .I(N__56422));
    InMux I__13985 (
            .O(N__56425),
            .I(N__56419));
    Odrv4 I__13984 (
            .O(N__56422),
            .I(\comm_spi.n22664 ));
    LocalMux I__13983 (
            .O(N__56419),
            .I(\comm_spi.n22664 ));
    InMux I__13982 (
            .O(N__56414),
            .I(N__56411));
    LocalMux I__13981 (
            .O(N__56411),
            .I(\comm_spi.n14612 ));
    SRMux I__13980 (
            .O(N__56408),
            .I(N__56405));
    LocalMux I__13979 (
            .O(N__56405),
            .I(N__56402));
    Sp12to4 I__13978 (
            .O(N__56402),
            .I(N__56399));
    Odrv12 I__13977 (
            .O(N__56399),
            .I(\comm_spi.iclk_N_763 ));
    InMux I__13976 (
            .O(N__56396),
            .I(N__56391));
    InMux I__13975 (
            .O(N__56395),
            .I(N__56388));
    InMux I__13974 (
            .O(N__56394),
            .I(N__56385));
    LocalMux I__13973 (
            .O(N__56391),
            .I(\comm_spi.n22688 ));
    LocalMux I__13972 (
            .O(N__56388),
            .I(\comm_spi.n22688 ));
    LocalMux I__13971 (
            .O(N__56385),
            .I(\comm_spi.n22688 ));
    CascadeMux I__13970 (
            .O(N__56378),
            .I(N__56374));
    InMux I__13969 (
            .O(N__56377),
            .I(N__56364));
    InMux I__13968 (
            .O(N__56374),
            .I(N__56348));
    InMux I__13967 (
            .O(N__56373),
            .I(N__56348));
    InMux I__13966 (
            .O(N__56372),
            .I(N__56348));
    InMux I__13965 (
            .O(N__56371),
            .I(N__56348));
    InMux I__13964 (
            .O(N__56370),
            .I(N__56345));
    InMux I__13963 (
            .O(N__56369),
            .I(N__56342));
    InMux I__13962 (
            .O(N__56368),
            .I(N__56326));
    InMux I__13961 (
            .O(N__56367),
            .I(N__56314));
    LocalMux I__13960 (
            .O(N__56364),
            .I(N__56310));
    InMux I__13959 (
            .O(N__56363),
            .I(N__56306));
    InMux I__13958 (
            .O(N__56362),
            .I(N__56292));
    InMux I__13957 (
            .O(N__56361),
            .I(N__56288));
    InMux I__13956 (
            .O(N__56360),
            .I(N__56283));
    InMux I__13955 (
            .O(N__56359),
            .I(N__56278));
    InMux I__13954 (
            .O(N__56358),
            .I(N__56275));
    InMux I__13953 (
            .O(N__56357),
            .I(N__56272));
    LocalMux I__13952 (
            .O(N__56348),
            .I(N__56265));
    LocalMux I__13951 (
            .O(N__56345),
            .I(N__56260));
    LocalMux I__13950 (
            .O(N__56342),
            .I(N__56257));
    InMux I__13949 (
            .O(N__56341),
            .I(N__56254));
    InMux I__13948 (
            .O(N__56340),
            .I(N__56241));
    InMux I__13947 (
            .O(N__56339),
            .I(N__56238));
    InMux I__13946 (
            .O(N__56338),
            .I(N__56231));
    InMux I__13945 (
            .O(N__56337),
            .I(N__56231));
    InMux I__13944 (
            .O(N__56336),
            .I(N__56226));
    InMux I__13943 (
            .O(N__56335),
            .I(N__56226));
    InMux I__13942 (
            .O(N__56334),
            .I(N__56223));
    InMux I__13941 (
            .O(N__56333),
            .I(N__56216));
    InMux I__13940 (
            .O(N__56332),
            .I(N__56216));
    InMux I__13939 (
            .O(N__56331),
            .I(N__56216));
    InMux I__13938 (
            .O(N__56330),
            .I(N__56213));
    InMux I__13937 (
            .O(N__56329),
            .I(N__56210));
    LocalMux I__13936 (
            .O(N__56326),
            .I(N__56207));
    InMux I__13935 (
            .O(N__56325),
            .I(N__56204));
    InMux I__13934 (
            .O(N__56324),
            .I(N__56197));
    InMux I__13933 (
            .O(N__56323),
            .I(N__56197));
    InMux I__13932 (
            .O(N__56322),
            .I(N__56197));
    InMux I__13931 (
            .O(N__56321),
            .I(N__56188));
    InMux I__13930 (
            .O(N__56320),
            .I(N__56188));
    InMux I__13929 (
            .O(N__56319),
            .I(N__56188));
    InMux I__13928 (
            .O(N__56318),
            .I(N__56188));
    InMux I__13927 (
            .O(N__56317),
            .I(N__56177));
    LocalMux I__13926 (
            .O(N__56314),
            .I(N__56174));
    InMux I__13925 (
            .O(N__56313),
            .I(N__56171));
    Span4Mux_h I__13924 (
            .O(N__56310),
            .I(N__56168));
    InMux I__13923 (
            .O(N__56309),
            .I(N__56163));
    LocalMux I__13922 (
            .O(N__56306),
            .I(N__56160));
    InMux I__13921 (
            .O(N__56305),
            .I(N__56154));
    InMux I__13920 (
            .O(N__56304),
            .I(N__56154));
    InMux I__13919 (
            .O(N__56303),
            .I(N__56145));
    InMux I__13918 (
            .O(N__56302),
            .I(N__56145));
    InMux I__13917 (
            .O(N__56301),
            .I(N__56145));
    InMux I__13916 (
            .O(N__56300),
            .I(N__56145));
    InMux I__13915 (
            .O(N__56299),
            .I(N__56140));
    InMux I__13914 (
            .O(N__56298),
            .I(N__56137));
    InMux I__13913 (
            .O(N__56297),
            .I(N__56132));
    InMux I__13912 (
            .O(N__56296),
            .I(N__56132));
    InMux I__13911 (
            .O(N__56295),
            .I(N__56129));
    LocalMux I__13910 (
            .O(N__56292),
            .I(N__56126));
    InMux I__13909 (
            .O(N__56291),
            .I(N__56123));
    LocalMux I__13908 (
            .O(N__56288),
            .I(N__56120));
    InMux I__13907 (
            .O(N__56287),
            .I(N__56115));
    InMux I__13906 (
            .O(N__56286),
            .I(N__56115));
    LocalMux I__13905 (
            .O(N__56283),
            .I(N__56112));
    InMux I__13904 (
            .O(N__56282),
            .I(N__56107));
    InMux I__13903 (
            .O(N__56281),
            .I(N__56107));
    LocalMux I__13902 (
            .O(N__56278),
            .I(N__56103));
    LocalMux I__13901 (
            .O(N__56275),
            .I(N__56100));
    LocalMux I__13900 (
            .O(N__56272),
            .I(N__56097));
    InMux I__13899 (
            .O(N__56271),
            .I(N__56094));
    InMux I__13898 (
            .O(N__56270),
            .I(N__56087));
    InMux I__13897 (
            .O(N__56269),
            .I(N__56087));
    InMux I__13896 (
            .O(N__56268),
            .I(N__56087));
    Span4Mux_h I__13895 (
            .O(N__56265),
            .I(N__56084));
    InMux I__13894 (
            .O(N__56264),
            .I(N__56079));
    InMux I__13893 (
            .O(N__56263),
            .I(N__56079));
    Span4Mux_v I__13892 (
            .O(N__56260),
            .I(N__56074));
    Span4Mux_h I__13891 (
            .O(N__56257),
            .I(N__56074));
    LocalMux I__13890 (
            .O(N__56254),
            .I(N__56068));
    InMux I__13889 (
            .O(N__56253),
            .I(N__56061));
    InMux I__13888 (
            .O(N__56252),
            .I(N__56061));
    InMux I__13887 (
            .O(N__56251),
            .I(N__56061));
    InMux I__13886 (
            .O(N__56250),
            .I(N__56056));
    InMux I__13885 (
            .O(N__56249),
            .I(N__56056));
    InMux I__13884 (
            .O(N__56248),
            .I(N__56051));
    InMux I__13883 (
            .O(N__56247),
            .I(N__56051));
    InMux I__13882 (
            .O(N__56246),
            .I(N__56046));
    InMux I__13881 (
            .O(N__56245),
            .I(N__56046));
    InMux I__13880 (
            .O(N__56244),
            .I(N__56043));
    LocalMux I__13879 (
            .O(N__56241),
            .I(N__56040));
    LocalMux I__13878 (
            .O(N__56238),
            .I(N__56037));
    InMux I__13877 (
            .O(N__56237),
            .I(N__56032));
    InMux I__13876 (
            .O(N__56236),
            .I(N__56032));
    LocalMux I__13875 (
            .O(N__56231),
            .I(N__56029));
    LocalMux I__13874 (
            .O(N__56226),
            .I(N__56020));
    LocalMux I__13873 (
            .O(N__56223),
            .I(N__56020));
    LocalMux I__13872 (
            .O(N__56216),
            .I(N__56020));
    LocalMux I__13871 (
            .O(N__56213),
            .I(N__56020));
    LocalMux I__13870 (
            .O(N__56210),
            .I(N__56009));
    Span4Mux_v I__13869 (
            .O(N__56207),
            .I(N__56009));
    LocalMux I__13868 (
            .O(N__56204),
            .I(N__56009));
    LocalMux I__13867 (
            .O(N__56197),
            .I(N__56009));
    LocalMux I__13866 (
            .O(N__56188),
            .I(N__56009));
    InMux I__13865 (
            .O(N__56187),
            .I(N__55999));
    InMux I__13864 (
            .O(N__56186),
            .I(N__55999));
    InMux I__13863 (
            .O(N__56185),
            .I(N__55999));
    InMux I__13862 (
            .O(N__56184),
            .I(N__55996));
    InMux I__13861 (
            .O(N__56183),
            .I(N__55993));
    InMux I__13860 (
            .O(N__56182),
            .I(N__55988));
    InMux I__13859 (
            .O(N__56181),
            .I(N__55988));
    InMux I__13858 (
            .O(N__56180),
            .I(N__55985));
    LocalMux I__13857 (
            .O(N__56177),
            .I(N__55978));
    Span4Mux_h I__13856 (
            .O(N__56174),
            .I(N__55978));
    LocalMux I__13855 (
            .O(N__56171),
            .I(N__55978));
    Span4Mux_v I__13854 (
            .O(N__56168),
            .I(N__55975));
    InMux I__13853 (
            .O(N__56167),
            .I(N__55970));
    InMux I__13852 (
            .O(N__56166),
            .I(N__55970));
    LocalMux I__13851 (
            .O(N__56163),
            .I(N__55967));
    Span4Mux_h I__13850 (
            .O(N__56160),
            .I(N__55964));
    InMux I__13849 (
            .O(N__56159),
            .I(N__55961));
    LocalMux I__13848 (
            .O(N__56154),
            .I(N__55956));
    LocalMux I__13847 (
            .O(N__56145),
            .I(N__55956));
    InMux I__13846 (
            .O(N__56144),
            .I(N__55953));
    InMux I__13845 (
            .O(N__56143),
            .I(N__55950));
    LocalMux I__13844 (
            .O(N__56140),
            .I(N__55940));
    LocalMux I__13843 (
            .O(N__56137),
            .I(N__55935));
    LocalMux I__13842 (
            .O(N__56132),
            .I(N__55935));
    LocalMux I__13841 (
            .O(N__56129),
            .I(N__55932));
    Span4Mux_h I__13840 (
            .O(N__56126),
            .I(N__55929));
    LocalMux I__13839 (
            .O(N__56123),
            .I(N__55924));
    Span4Mux_h I__13838 (
            .O(N__56120),
            .I(N__55924));
    LocalMux I__13837 (
            .O(N__56115),
            .I(N__55917));
    Span4Mux_v I__13836 (
            .O(N__56112),
            .I(N__55917));
    LocalMux I__13835 (
            .O(N__56107),
            .I(N__55917));
    InMux I__13834 (
            .O(N__56106),
            .I(N__55914));
    Span4Mux_h I__13833 (
            .O(N__56103),
            .I(N__55909));
    Span4Mux_h I__13832 (
            .O(N__56100),
            .I(N__55909));
    Span4Mux_h I__13831 (
            .O(N__56097),
            .I(N__55900));
    LocalMux I__13830 (
            .O(N__56094),
            .I(N__55900));
    LocalMux I__13829 (
            .O(N__56087),
            .I(N__55900));
    Span4Mux_v I__13828 (
            .O(N__56084),
            .I(N__55900));
    LocalMux I__13827 (
            .O(N__56079),
            .I(N__55897));
    Span4Mux_v I__13826 (
            .O(N__56074),
            .I(N__55894));
    InMux I__13825 (
            .O(N__56073),
            .I(N__55891));
    InMux I__13824 (
            .O(N__56072),
            .I(N__55886));
    InMux I__13823 (
            .O(N__56071),
            .I(N__55886));
    Span4Mux_v I__13822 (
            .O(N__56068),
            .I(N__55881));
    LocalMux I__13821 (
            .O(N__56061),
            .I(N__55881));
    LocalMux I__13820 (
            .O(N__56056),
            .I(N__55876));
    LocalMux I__13819 (
            .O(N__56051),
            .I(N__55876));
    LocalMux I__13818 (
            .O(N__56046),
            .I(N__55873));
    LocalMux I__13817 (
            .O(N__56043),
            .I(N__55864));
    Span4Mux_h I__13816 (
            .O(N__56040),
            .I(N__55864));
    Span4Mux_h I__13815 (
            .O(N__56037),
            .I(N__55864));
    LocalMux I__13814 (
            .O(N__56032),
            .I(N__55864));
    Span4Mux_h I__13813 (
            .O(N__56029),
            .I(N__55857));
    Span4Mux_v I__13812 (
            .O(N__56020),
            .I(N__55857));
    Span4Mux_v I__13811 (
            .O(N__56009),
            .I(N__55857));
    InMux I__13810 (
            .O(N__56008),
            .I(N__55850));
    InMux I__13809 (
            .O(N__56007),
            .I(N__55850));
    InMux I__13808 (
            .O(N__56006),
            .I(N__55850));
    LocalMux I__13807 (
            .O(N__55999),
            .I(N__55847));
    LocalMux I__13806 (
            .O(N__55996),
            .I(N__55842));
    LocalMux I__13805 (
            .O(N__55993),
            .I(N__55842));
    LocalMux I__13804 (
            .O(N__55988),
            .I(N__55839));
    LocalMux I__13803 (
            .O(N__55985),
            .I(N__55836));
    Span4Mux_v I__13802 (
            .O(N__55978),
            .I(N__55831));
    Span4Mux_v I__13801 (
            .O(N__55975),
            .I(N__55831));
    LocalMux I__13800 (
            .O(N__55970),
            .I(N__55818));
    Span4Mux_v I__13799 (
            .O(N__55967),
            .I(N__55818));
    Span4Mux_v I__13798 (
            .O(N__55964),
            .I(N__55818));
    LocalMux I__13797 (
            .O(N__55961),
            .I(N__55818));
    Span4Mux_h I__13796 (
            .O(N__55956),
            .I(N__55818));
    LocalMux I__13795 (
            .O(N__55953),
            .I(N__55818));
    LocalMux I__13794 (
            .O(N__55950),
            .I(N__55813));
    InMux I__13793 (
            .O(N__55949),
            .I(N__55810));
    InMux I__13792 (
            .O(N__55948),
            .I(N__55803));
    InMux I__13791 (
            .O(N__55947),
            .I(N__55803));
    InMux I__13790 (
            .O(N__55946),
            .I(N__55803));
    InMux I__13789 (
            .O(N__55945),
            .I(N__55798));
    InMux I__13788 (
            .O(N__55944),
            .I(N__55798));
    InMux I__13787 (
            .O(N__55943),
            .I(N__55795));
    Span12Mux_h I__13786 (
            .O(N__55940),
            .I(N__55788));
    Span12Mux_h I__13785 (
            .O(N__55935),
            .I(N__55788));
    Span12Mux_h I__13784 (
            .O(N__55932),
            .I(N__55788));
    Span4Mux_h I__13783 (
            .O(N__55929),
            .I(N__55781));
    Span4Mux_v I__13782 (
            .O(N__55924),
            .I(N__55781));
    Span4Mux_h I__13781 (
            .O(N__55917),
            .I(N__55781));
    LocalMux I__13780 (
            .O(N__55914),
            .I(N__55770));
    Span4Mux_v I__13779 (
            .O(N__55909),
            .I(N__55770));
    Span4Mux_h I__13778 (
            .O(N__55900),
            .I(N__55770));
    Span4Mux_h I__13777 (
            .O(N__55897),
            .I(N__55770));
    Span4Mux_h I__13776 (
            .O(N__55894),
            .I(N__55770));
    LocalMux I__13775 (
            .O(N__55891),
            .I(N__55755));
    LocalMux I__13774 (
            .O(N__55886),
            .I(N__55755));
    Span4Mux_v I__13773 (
            .O(N__55881),
            .I(N__55755));
    Span4Mux_h I__13772 (
            .O(N__55876),
            .I(N__55755));
    Span4Mux_h I__13771 (
            .O(N__55873),
            .I(N__55755));
    Span4Mux_v I__13770 (
            .O(N__55864),
            .I(N__55755));
    Span4Mux_h I__13769 (
            .O(N__55857),
            .I(N__55755));
    LocalMux I__13768 (
            .O(N__55850),
            .I(N__55740));
    Span4Mux_v I__13767 (
            .O(N__55847),
            .I(N__55740));
    Span4Mux_v I__13766 (
            .O(N__55842),
            .I(N__55740));
    Span4Mux_h I__13765 (
            .O(N__55839),
            .I(N__55740));
    Span4Mux_h I__13764 (
            .O(N__55836),
            .I(N__55740));
    Span4Mux_h I__13763 (
            .O(N__55831),
            .I(N__55740));
    Span4Mux_v I__13762 (
            .O(N__55818),
            .I(N__55740));
    InMux I__13761 (
            .O(N__55817),
            .I(N__55735));
    InMux I__13760 (
            .O(N__55816),
            .I(N__55735));
    Odrv4 I__13759 (
            .O(N__55813),
            .I(comm_cmd_0));
    LocalMux I__13758 (
            .O(N__55810),
            .I(comm_cmd_0));
    LocalMux I__13757 (
            .O(N__55803),
            .I(comm_cmd_0));
    LocalMux I__13756 (
            .O(N__55798),
            .I(comm_cmd_0));
    LocalMux I__13755 (
            .O(N__55795),
            .I(comm_cmd_0));
    Odrv12 I__13754 (
            .O(N__55788),
            .I(comm_cmd_0));
    Odrv4 I__13753 (
            .O(N__55781),
            .I(comm_cmd_0));
    Odrv4 I__13752 (
            .O(N__55770),
            .I(comm_cmd_0));
    Odrv4 I__13751 (
            .O(N__55755),
            .I(comm_cmd_0));
    Odrv4 I__13750 (
            .O(N__55740),
            .I(comm_cmd_0));
    LocalMux I__13749 (
            .O(N__55735),
            .I(comm_cmd_0));
    InMux I__13748 (
            .O(N__55712),
            .I(N__55709));
    LocalMux I__13747 (
            .O(N__55709),
            .I(N__55706));
    Span4Mux_h I__13746 (
            .O(N__55706),
            .I(N__55703));
    Odrv4 I__13745 (
            .O(N__55703),
            .I(buf_data_iac_10));
    CascadeMux I__13744 (
            .O(N__55700),
            .I(N__55697));
    InMux I__13743 (
            .O(N__55697),
            .I(N__55694));
    LocalMux I__13742 (
            .O(N__55694),
            .I(N__55691));
    Span4Mux_h I__13741 (
            .O(N__55691),
            .I(N__55688));
    Odrv4 I__13740 (
            .O(N__55688),
            .I(n21320));
    InMux I__13739 (
            .O(N__55685),
            .I(N__55681));
    InMux I__13738 (
            .O(N__55684),
            .I(N__55678));
    LocalMux I__13737 (
            .O(N__55681),
            .I(N__55673));
    LocalMux I__13736 (
            .O(N__55678),
            .I(N__55673));
    Odrv12 I__13735 (
            .O(N__55673),
            .I(\comm_spi.n14655 ));
    SRMux I__13734 (
            .O(N__55670),
            .I(N__55667));
    LocalMux I__13733 (
            .O(N__55667),
            .I(N__55664));
    Span4Mux_h I__13732 (
            .O(N__55664),
            .I(N__55661));
    Span4Mux_v I__13731 (
            .O(N__55661),
            .I(N__55658));
    Odrv4 I__13730 (
            .O(N__55658),
            .I(\comm_spi.data_tx_7__N_778 ));
    InMux I__13729 (
            .O(N__55655),
            .I(N__55650));
    InMux I__13728 (
            .O(N__55654),
            .I(N__55647));
    InMux I__13727 (
            .O(N__55653),
            .I(N__55644));
    LocalMux I__13726 (
            .O(N__55650),
            .I(\comm_spi.n22673 ));
    LocalMux I__13725 (
            .O(N__55647),
            .I(\comm_spi.n22673 ));
    LocalMux I__13724 (
            .O(N__55644),
            .I(\comm_spi.n22673 ));
    InMux I__13723 (
            .O(N__55637),
            .I(N__55633));
    InMux I__13722 (
            .O(N__55636),
            .I(N__55630));
    LocalMux I__13721 (
            .O(N__55633),
            .I(N__55627));
    LocalMux I__13720 (
            .O(N__55630),
            .I(N__55624));
    Odrv4 I__13719 (
            .O(N__55627),
            .I(\comm_spi.n14651 ));
    Odrv4 I__13718 (
            .O(N__55624),
            .I(\comm_spi.n14651 ));
    InMux I__13717 (
            .O(N__55619),
            .I(N__55615));
    InMux I__13716 (
            .O(N__55618),
            .I(N__55612));
    LocalMux I__13715 (
            .O(N__55615),
            .I(N__55607));
    LocalMux I__13714 (
            .O(N__55612),
            .I(N__55607));
    Odrv12 I__13713 (
            .O(N__55607),
            .I(\comm_spi.n14654 ));
    SRMux I__13712 (
            .O(N__55604),
            .I(N__55601));
    LocalMux I__13711 (
            .O(N__55601),
            .I(N__55598));
    Span4Mux_h I__13710 (
            .O(N__55598),
            .I(N__55595));
    Odrv4 I__13709 (
            .O(N__55595),
            .I(\comm_spi.data_tx_7__N_781 ));
    InMux I__13708 (
            .O(N__55592),
            .I(N__55589));
    LocalMux I__13707 (
            .O(N__55589),
            .I(buf_data_iac_23));
    InMux I__13706 (
            .O(N__55586),
            .I(N__55583));
    LocalMux I__13705 (
            .O(N__55583),
            .I(N__55580));
    Span4Mux_v I__13704 (
            .O(N__55580),
            .I(N__55577));
    Span4Mux_h I__13703 (
            .O(N__55577),
            .I(N__55574));
    Span4Mux_h I__13702 (
            .O(N__55574),
            .I(N__55571));
    Sp12to4 I__13701 (
            .O(N__55571),
            .I(N__55568));
    Odrv12 I__13700 (
            .O(N__55568),
            .I(n21204));
    IoInMux I__13699 (
            .O(N__55565),
            .I(N__55562));
    LocalMux I__13698 (
            .O(N__55562),
            .I(N__55559));
    Span4Mux_s3_h I__13697 (
            .O(N__55559),
            .I(N__55556));
    Span4Mux_v I__13696 (
            .O(N__55556),
            .I(N__55553));
    Span4Mux_v I__13695 (
            .O(N__55553),
            .I(N__55550));
    Span4Mux_h I__13694 (
            .O(N__55550),
            .I(N__55547));
    Odrv4 I__13693 (
            .O(N__55547),
            .I(ICE_SPI_MISO));
    InMux I__13692 (
            .O(N__55544),
            .I(N__55541));
    LocalMux I__13691 (
            .O(N__55541),
            .I(\comm_spi.n14621 ));
    InMux I__13690 (
            .O(N__55538),
            .I(N__55535));
    LocalMux I__13689 (
            .O(N__55535),
            .I(N__55531));
    InMux I__13688 (
            .O(N__55534),
            .I(N__55528));
    Span4Mux_h I__13687 (
            .O(N__55531),
            .I(N__55523));
    LocalMux I__13686 (
            .O(N__55528),
            .I(N__55523));
    Odrv4 I__13685 (
            .O(N__55523),
            .I(\comm_spi.n14626 ));
    InMux I__13684 (
            .O(N__55520),
            .I(N__55517));
    LocalMux I__13683 (
            .O(N__55517),
            .I(N__55514));
    Odrv4 I__13682 (
            .O(N__55514),
            .I(\comm_spi.n14620 ));
    InMux I__13681 (
            .O(N__55511),
            .I(N__55507));
    InMux I__13680 (
            .O(N__55510),
            .I(N__55504));
    LocalMux I__13679 (
            .O(N__55507),
            .I(N__55501));
    LocalMux I__13678 (
            .O(N__55504),
            .I(N__55498));
    Span4Mux_v I__13677 (
            .O(N__55501),
            .I(N__55492));
    Span4Mux_h I__13676 (
            .O(N__55498),
            .I(N__55492));
    InMux I__13675 (
            .O(N__55497),
            .I(N__55489));
    Span4Mux_v I__13674 (
            .O(N__55492),
            .I(N__55484));
    LocalMux I__13673 (
            .O(N__55489),
            .I(N__55484));
    Span4Mux_v I__13672 (
            .O(N__55484),
            .I(N__55481));
    Odrv4 I__13671 (
            .O(N__55481),
            .I(comm_tx_buf_6));
    InMux I__13670 (
            .O(N__55478),
            .I(N__55473));
    InMux I__13669 (
            .O(N__55477),
            .I(N__55470));
    InMux I__13668 (
            .O(N__55476),
            .I(N__55466));
    LocalMux I__13667 (
            .O(N__55473),
            .I(N__55460));
    LocalMux I__13666 (
            .O(N__55470),
            .I(N__55460));
    InMux I__13665 (
            .O(N__55469),
            .I(N__55457));
    LocalMux I__13664 (
            .O(N__55466),
            .I(N__55454));
    InMux I__13663 (
            .O(N__55465),
            .I(N__55451));
    Span4Mux_v I__13662 (
            .O(N__55460),
            .I(N__55445));
    LocalMux I__13661 (
            .O(N__55457),
            .I(N__55445));
    Span4Mux_v I__13660 (
            .O(N__55454),
            .I(N__55440));
    LocalMux I__13659 (
            .O(N__55451),
            .I(N__55440));
    InMux I__13658 (
            .O(N__55450),
            .I(N__55437));
    Span4Mux_h I__13657 (
            .O(N__55445),
            .I(N__55434));
    Odrv4 I__13656 (
            .O(N__55440),
            .I(\comm_spi.n14619 ));
    LocalMux I__13655 (
            .O(N__55437),
            .I(\comm_spi.n14619 ));
    Odrv4 I__13654 (
            .O(N__55434),
            .I(\comm_spi.n14619 ));
    InMux I__13653 (
            .O(N__55427),
            .I(N__55424));
    LocalMux I__13652 (
            .O(N__55424),
            .I(N__55420));
    InMux I__13651 (
            .O(N__55423),
            .I(N__55417));
    Odrv4 I__13650 (
            .O(N__55420),
            .I(\comm_spi.n14627 ));
    LocalMux I__13649 (
            .O(N__55417),
            .I(\comm_spi.n14627 ));
    InMux I__13648 (
            .O(N__55412),
            .I(N__55408));
    InMux I__13647 (
            .O(N__55411),
            .I(N__55405));
    LocalMux I__13646 (
            .O(N__55408),
            .I(\comm_spi.n14624 ));
    LocalMux I__13645 (
            .O(N__55405),
            .I(\comm_spi.n14624 ));
    InMux I__13644 (
            .O(N__55400),
            .I(N__55397));
    LocalMux I__13643 (
            .O(N__55397),
            .I(N__55394));
    Span4Mux_v I__13642 (
            .O(N__55394),
            .I(N__55390));
    InMux I__13641 (
            .O(N__55393),
            .I(N__55387));
    Span4Mux_h I__13640 (
            .O(N__55390),
            .I(N__55381));
    LocalMux I__13639 (
            .O(N__55387),
            .I(N__55381));
    InMux I__13638 (
            .O(N__55386),
            .I(N__55378));
    Odrv4 I__13637 (
            .O(N__55381),
            .I(\comm_spi.n22682 ));
    LocalMux I__13636 (
            .O(N__55378),
            .I(\comm_spi.n22682 ));
    InMux I__13635 (
            .O(N__55373),
            .I(N__55370));
    LocalMux I__13634 (
            .O(N__55370),
            .I(N__55367));
    Sp12to4 I__13633 (
            .O(N__55367),
            .I(N__55363));
    InMux I__13632 (
            .O(N__55366),
            .I(N__55360));
    Span12Mux_h I__13631 (
            .O(N__55363),
            .I(N__55357));
    LocalMux I__13630 (
            .O(N__55360),
            .I(N__55354));
    Odrv12 I__13629 (
            .O(N__55357),
            .I(\comm_spi.n14638 ));
    Odrv4 I__13628 (
            .O(N__55354),
            .I(\comm_spi.n14638 ));
    InMux I__13627 (
            .O(N__55349),
            .I(N__55346));
    LocalMux I__13626 (
            .O(N__55346),
            .I(N__55343));
    Span4Mux_h I__13625 (
            .O(N__55343),
            .I(N__55340));
    Span4Mux_h I__13624 (
            .O(N__55340),
            .I(N__55336));
    InMux I__13623 (
            .O(N__55339),
            .I(N__55333));
    Sp12to4 I__13622 (
            .O(N__55336),
            .I(N__55328));
    LocalMux I__13621 (
            .O(N__55333),
            .I(N__55328));
    Odrv12 I__13620 (
            .O(N__55328),
            .I(\comm_spi.n14639 ));
    SRMux I__13619 (
            .O(N__55325),
            .I(N__55322));
    LocalMux I__13618 (
            .O(N__55322),
            .I(\comm_spi.data_tx_7__N_787 ));
    InMux I__13617 (
            .O(N__55319),
            .I(N__55315));
    InMux I__13616 (
            .O(N__55318),
            .I(N__55312));
    LocalMux I__13615 (
            .O(N__55315),
            .I(N__55308));
    LocalMux I__13614 (
            .O(N__55312),
            .I(N__55305));
    InMux I__13613 (
            .O(N__55311),
            .I(N__55302));
    Span4Mux_v I__13612 (
            .O(N__55308),
            .I(N__55299));
    Span4Mux_v I__13611 (
            .O(N__55305),
            .I(N__55294));
    LocalMux I__13610 (
            .O(N__55302),
            .I(N__55294));
    Sp12to4 I__13609 (
            .O(N__55299),
            .I(N__55291));
    Span4Mux_h I__13608 (
            .O(N__55294),
            .I(N__55288));
    Span12Mux_h I__13607 (
            .O(N__55291),
            .I(N__55283));
    Sp12to4 I__13606 (
            .O(N__55288),
            .I(N__55283));
    Odrv12 I__13605 (
            .O(N__55283),
            .I(comm_tx_buf_3));
    InMux I__13604 (
            .O(N__55280),
            .I(N__55276));
    InMux I__13603 (
            .O(N__55279),
            .I(N__55273));
    LocalMux I__13602 (
            .O(N__55276),
            .I(N__55267));
    LocalMux I__13601 (
            .O(N__55273),
            .I(N__55267));
    InMux I__13600 (
            .O(N__55272),
            .I(N__55264));
    Span4Mux_v I__13599 (
            .O(N__55267),
            .I(N__55259));
    LocalMux I__13598 (
            .O(N__55264),
            .I(N__55259));
    Span4Mux_v I__13597 (
            .O(N__55259),
            .I(N__55256));
    Span4Mux_v I__13596 (
            .O(N__55256),
            .I(N__55253));
    Span4Mux_h I__13595 (
            .O(N__55253),
            .I(N__55250));
    Odrv4 I__13594 (
            .O(N__55250),
            .I(comm_tx_buf_4));
    InMux I__13593 (
            .O(N__55247),
            .I(N__55241));
    InMux I__13592 (
            .O(N__55246),
            .I(N__55241));
    LocalMux I__13591 (
            .O(N__55241),
            .I(N__55238));
    Span4Mux_h I__13590 (
            .O(N__55238),
            .I(N__55234));
    InMux I__13589 (
            .O(N__55237),
            .I(N__55231));
    Sp12to4 I__13588 (
            .O(N__55234),
            .I(N__55226));
    LocalMux I__13587 (
            .O(N__55231),
            .I(N__55226));
    Span12Mux_v I__13586 (
            .O(N__55226),
            .I(N__55223));
    Odrv12 I__13585 (
            .O(N__55223),
            .I(comm_tx_buf_5));
    InMux I__13584 (
            .O(N__55220),
            .I(N__55215));
    InMux I__13583 (
            .O(N__55219),
            .I(N__55212));
    InMux I__13582 (
            .O(N__55218),
            .I(N__55209));
    LocalMux I__13581 (
            .O(N__55215),
            .I(\comm_spi.n22679 ));
    LocalMux I__13580 (
            .O(N__55212),
            .I(\comm_spi.n22679 ));
    LocalMux I__13579 (
            .O(N__55209),
            .I(\comm_spi.n22679 ));
    InMux I__13578 (
            .O(N__55202),
            .I(N__55198));
    InMux I__13577 (
            .O(N__55201),
            .I(N__55195));
    LocalMux I__13576 (
            .O(N__55198),
            .I(N__55190));
    LocalMux I__13575 (
            .O(N__55195),
            .I(N__55190));
    Odrv12 I__13574 (
            .O(N__55190),
            .I(\comm_spi.n14642 ));
    InMux I__13573 (
            .O(N__55187),
            .I(N__55183));
    InMux I__13572 (
            .O(N__55186),
            .I(N__55180));
    LocalMux I__13571 (
            .O(N__55183),
            .I(N__55175));
    LocalMux I__13570 (
            .O(N__55180),
            .I(N__55175));
    Odrv4 I__13569 (
            .O(N__55175),
            .I(\comm_spi.n14643 ));
    SRMux I__13568 (
            .O(N__55172),
            .I(N__55169));
    LocalMux I__13567 (
            .O(N__55169),
            .I(N__55166));
    Span4Mux_v I__13566 (
            .O(N__55166),
            .I(N__55163));
    Odrv4 I__13565 (
            .O(N__55163),
            .I(\comm_spi.data_tx_7__N_784 ));
    InMux I__13564 (
            .O(N__55160),
            .I(N__55157));
    LocalMux I__13563 (
            .O(N__55157),
            .I(N__55154));
    Span4Mux_v I__13562 (
            .O(N__55154),
            .I(N__55149));
    InMux I__13561 (
            .O(N__55153),
            .I(N__55144));
    InMux I__13560 (
            .O(N__55152),
            .I(N__55144));
    Span4Mux_v I__13559 (
            .O(N__55149),
            .I(N__55141));
    LocalMux I__13558 (
            .O(N__55144),
            .I(N__55138));
    Sp12to4 I__13557 (
            .O(N__55141),
            .I(N__55135));
    Span4Mux_h I__13556 (
            .O(N__55138),
            .I(N__55132));
    Odrv12 I__13555 (
            .O(N__55135),
            .I(comm_tx_buf_2));
    Odrv4 I__13554 (
            .O(N__55132),
            .I(comm_tx_buf_2));
    InMux I__13553 (
            .O(N__55127),
            .I(N__55124));
    LocalMux I__13552 (
            .O(N__55124),
            .I(N__55120));
    InMux I__13551 (
            .O(N__55123),
            .I(N__55117));
    Span4Mux_v I__13550 (
            .O(N__55120),
            .I(N__55112));
    LocalMux I__13549 (
            .O(N__55117),
            .I(N__55112));
    Span4Mux_v I__13548 (
            .O(N__55112),
            .I(N__55109));
    Odrv4 I__13547 (
            .O(N__55109),
            .I(\comm_spi.imosi ));
    SRMux I__13546 (
            .O(N__55106),
            .I(N__55103));
    LocalMux I__13545 (
            .O(N__55103),
            .I(N__55100));
    Span4Mux_v I__13544 (
            .O(N__55100),
            .I(N__55097));
    Odrv4 I__13543 (
            .O(N__55097),
            .I(\comm_spi.DOUT_7__N_748 ));
    SRMux I__13542 (
            .O(N__55094),
            .I(N__55091));
    LocalMux I__13541 (
            .O(N__55091),
            .I(N__55088));
    Span4Mux_h I__13540 (
            .O(N__55088),
            .I(N__55085));
    Odrv4 I__13539 (
            .O(N__55085),
            .I(\comm_spi.imosi_N_753 ));
    SRMux I__13538 (
            .O(N__55082),
            .I(N__55079));
    LocalMux I__13537 (
            .O(N__55079),
            .I(N__55076));
    Span4Mux_v I__13536 (
            .O(N__55076),
            .I(N__55073));
    Odrv4 I__13535 (
            .O(N__55073),
            .I(\comm_spi.data_tx_7__N_790 ));
    InMux I__13534 (
            .O(N__55070),
            .I(N__55065));
    InMux I__13533 (
            .O(N__55069),
            .I(N__55062));
    InMux I__13532 (
            .O(N__55068),
            .I(N__55059));
    LocalMux I__13531 (
            .O(N__55065),
            .I(\comm_spi.n22685 ));
    LocalMux I__13530 (
            .O(N__55062),
            .I(\comm_spi.n22685 ));
    LocalMux I__13529 (
            .O(N__55059),
            .I(\comm_spi.n22685 ));
    SRMux I__13528 (
            .O(N__55052),
            .I(N__55049));
    LocalMux I__13527 (
            .O(N__55049),
            .I(N__55046));
    Odrv4 I__13526 (
            .O(N__55046),
            .I(\comm_spi.data_tx_7__N_772 ));
    InMux I__13525 (
            .O(N__55043),
            .I(N__55040));
    LocalMux I__13524 (
            .O(N__55040),
            .I(N__55036));
    InMux I__13523 (
            .O(N__55039),
            .I(N__55033));
    Odrv4 I__13522 (
            .O(N__55036),
            .I(\comm_spi.n14634 ));
    LocalMux I__13521 (
            .O(N__55033),
            .I(\comm_spi.n14634 ));
    InMux I__13520 (
            .O(N__55028),
            .I(N__55024));
    InMux I__13519 (
            .O(N__55027),
            .I(N__55021));
    LocalMux I__13518 (
            .O(N__55024),
            .I(N__55017));
    LocalMux I__13517 (
            .O(N__55021),
            .I(N__55014));
    InMux I__13516 (
            .O(N__55020),
            .I(N__55011));
    Span4Mux_v I__13515 (
            .O(N__55017),
            .I(N__55008));
    Span4Mux_v I__13514 (
            .O(N__55014),
            .I(N__55003));
    LocalMux I__13513 (
            .O(N__55011),
            .I(N__55003));
    Span4Mux_v I__13512 (
            .O(N__55008),
            .I(N__55000));
    Span4Mux_v I__13511 (
            .O(N__55003),
            .I(N__54997));
    Odrv4 I__13510 (
            .O(N__55000),
            .I(comm_tx_buf_1));
    Odrv4 I__13509 (
            .O(N__54997),
            .I(comm_tx_buf_1));
    SRMux I__13508 (
            .O(N__54992),
            .I(N__54989));
    LocalMux I__13507 (
            .O(N__54989),
            .I(N__54986));
    Odrv4 I__13506 (
            .O(N__54986),
            .I(\comm_spi.data_tx_7__N_773 ));
    CascadeMux I__13505 (
            .O(N__54983),
            .I(N__54978));
    InMux I__13504 (
            .O(N__54982),
            .I(N__54968));
    InMux I__13503 (
            .O(N__54981),
            .I(N__54955));
    InMux I__13502 (
            .O(N__54978),
            .I(N__54955));
    CascadeMux I__13501 (
            .O(N__54977),
            .I(N__54950));
    InMux I__13500 (
            .O(N__54976),
            .I(N__54932));
    InMux I__13499 (
            .O(N__54975),
            .I(N__54932));
    InMux I__13498 (
            .O(N__54974),
            .I(N__54932));
    InMux I__13497 (
            .O(N__54973),
            .I(N__54932));
    InMux I__13496 (
            .O(N__54972),
            .I(N__54932));
    InMux I__13495 (
            .O(N__54971),
            .I(N__54932));
    LocalMux I__13494 (
            .O(N__54968),
            .I(N__54929));
    InMux I__13493 (
            .O(N__54967),
            .I(N__54924));
    InMux I__13492 (
            .O(N__54966),
            .I(N__54924));
    InMux I__13491 (
            .O(N__54965),
            .I(N__54917));
    InMux I__13490 (
            .O(N__54964),
            .I(N__54917));
    InMux I__13489 (
            .O(N__54963),
            .I(N__54914));
    CascadeMux I__13488 (
            .O(N__54962),
            .I(N__54908));
    CascadeMux I__13487 (
            .O(N__54961),
            .I(N__54904));
    CascadeMux I__13486 (
            .O(N__54960),
            .I(N__54896));
    LocalMux I__13485 (
            .O(N__54955),
            .I(N__54884));
    InMux I__13484 (
            .O(N__54954),
            .I(N__54879));
    InMux I__13483 (
            .O(N__54953),
            .I(N__54879));
    InMux I__13482 (
            .O(N__54950),
            .I(N__54872));
    InMux I__13481 (
            .O(N__54949),
            .I(N__54872));
    InMux I__13480 (
            .O(N__54948),
            .I(N__54872));
    InMux I__13479 (
            .O(N__54947),
            .I(N__54864));
    InMux I__13478 (
            .O(N__54946),
            .I(N__54859));
    InMux I__13477 (
            .O(N__54945),
            .I(N__54859));
    LocalMux I__13476 (
            .O(N__54932),
            .I(N__54854));
    Span4Mux_v I__13475 (
            .O(N__54929),
            .I(N__54854));
    LocalMux I__13474 (
            .O(N__54924),
            .I(N__54851));
    InMux I__13473 (
            .O(N__54923),
            .I(N__54848));
    InMux I__13472 (
            .O(N__54922),
            .I(N__54843));
    LocalMux I__13471 (
            .O(N__54917),
            .I(N__54838));
    LocalMux I__13470 (
            .O(N__54914),
            .I(N__54838));
    InMux I__13469 (
            .O(N__54913),
            .I(N__54833));
    InMux I__13468 (
            .O(N__54912),
            .I(N__54830));
    InMux I__13467 (
            .O(N__54911),
            .I(N__54825));
    InMux I__13466 (
            .O(N__54908),
            .I(N__54818));
    InMux I__13465 (
            .O(N__54907),
            .I(N__54818));
    InMux I__13464 (
            .O(N__54904),
            .I(N__54811));
    InMux I__13463 (
            .O(N__54903),
            .I(N__54811));
    InMux I__13462 (
            .O(N__54902),
            .I(N__54811));
    InMux I__13461 (
            .O(N__54901),
            .I(N__54796));
    InMux I__13460 (
            .O(N__54900),
            .I(N__54796));
    InMux I__13459 (
            .O(N__54899),
            .I(N__54796));
    InMux I__13458 (
            .O(N__54896),
            .I(N__54785));
    InMux I__13457 (
            .O(N__54895),
            .I(N__54785));
    InMux I__13456 (
            .O(N__54894),
            .I(N__54785));
    InMux I__13455 (
            .O(N__54893),
            .I(N__54785));
    InMux I__13454 (
            .O(N__54892),
            .I(N__54785));
    InMux I__13453 (
            .O(N__54891),
            .I(N__54776));
    InMux I__13452 (
            .O(N__54890),
            .I(N__54776));
    InMux I__13451 (
            .O(N__54889),
            .I(N__54776));
    InMux I__13450 (
            .O(N__54888),
            .I(N__54776));
    InMux I__13449 (
            .O(N__54887),
            .I(N__54773));
    Span4Mux_v I__13448 (
            .O(N__54884),
            .I(N__54766));
    LocalMux I__13447 (
            .O(N__54879),
            .I(N__54766));
    LocalMux I__13446 (
            .O(N__54872),
            .I(N__54766));
    InMux I__13445 (
            .O(N__54871),
            .I(N__54758));
    InMux I__13444 (
            .O(N__54870),
            .I(N__54758));
    InMux I__13443 (
            .O(N__54869),
            .I(N__54751));
    InMux I__13442 (
            .O(N__54868),
            .I(N__54751));
    InMux I__13441 (
            .O(N__54867),
            .I(N__54751));
    LocalMux I__13440 (
            .O(N__54864),
            .I(N__54740));
    LocalMux I__13439 (
            .O(N__54859),
            .I(N__54740));
    Span4Mux_v I__13438 (
            .O(N__54854),
            .I(N__54740));
    Span4Mux_h I__13437 (
            .O(N__54851),
            .I(N__54740));
    LocalMux I__13436 (
            .O(N__54848),
            .I(N__54740));
    InMux I__13435 (
            .O(N__54847),
            .I(N__54737));
    InMux I__13434 (
            .O(N__54846),
            .I(N__54732));
    LocalMux I__13433 (
            .O(N__54843),
            .I(N__54727));
    Span4Mux_v I__13432 (
            .O(N__54838),
            .I(N__54727));
    CascadeMux I__13431 (
            .O(N__54837),
            .I(N__54724));
    SRMux I__13430 (
            .O(N__54836),
            .I(N__54719));
    LocalMux I__13429 (
            .O(N__54833),
            .I(N__54714));
    LocalMux I__13428 (
            .O(N__54830),
            .I(N__54711));
    InMux I__13427 (
            .O(N__54829),
            .I(N__54700));
    InMux I__13426 (
            .O(N__54828),
            .I(N__54700));
    LocalMux I__13425 (
            .O(N__54825),
            .I(N__54697));
    InMux I__13424 (
            .O(N__54824),
            .I(N__54694));
    InMux I__13423 (
            .O(N__54823),
            .I(N__54691));
    LocalMux I__13422 (
            .O(N__54818),
            .I(N__54686));
    LocalMux I__13421 (
            .O(N__54811),
            .I(N__54686));
    InMux I__13420 (
            .O(N__54810),
            .I(N__54677));
    InMux I__13419 (
            .O(N__54809),
            .I(N__54677));
    InMux I__13418 (
            .O(N__54808),
            .I(N__54677));
    InMux I__13417 (
            .O(N__54807),
            .I(N__54677));
    InMux I__13416 (
            .O(N__54806),
            .I(N__54668));
    InMux I__13415 (
            .O(N__54805),
            .I(N__54668));
    InMux I__13414 (
            .O(N__54804),
            .I(N__54668));
    InMux I__13413 (
            .O(N__54803),
            .I(N__54668));
    LocalMux I__13412 (
            .O(N__54796),
            .I(N__54661));
    LocalMux I__13411 (
            .O(N__54785),
            .I(N__54661));
    LocalMux I__13410 (
            .O(N__54776),
            .I(N__54661));
    LocalMux I__13409 (
            .O(N__54773),
            .I(N__54656));
    Span4Mux_h I__13408 (
            .O(N__54766),
            .I(N__54656));
    InMux I__13407 (
            .O(N__54765),
            .I(N__54649));
    InMux I__13406 (
            .O(N__54764),
            .I(N__54649));
    InMux I__13405 (
            .O(N__54763),
            .I(N__54646));
    LocalMux I__13404 (
            .O(N__54758),
            .I(N__54641));
    LocalMux I__13403 (
            .O(N__54751),
            .I(N__54641));
    Span4Mux_v I__13402 (
            .O(N__54740),
            .I(N__54638));
    LocalMux I__13401 (
            .O(N__54737),
            .I(N__54632));
    InMux I__13400 (
            .O(N__54736),
            .I(N__54629));
    InMux I__13399 (
            .O(N__54735),
            .I(N__54626));
    LocalMux I__13398 (
            .O(N__54732),
            .I(N__54621));
    Span4Mux_v I__13397 (
            .O(N__54727),
            .I(N__54621));
    InMux I__13396 (
            .O(N__54724),
            .I(N__54616));
    InMux I__13395 (
            .O(N__54723),
            .I(N__54616));
    InMux I__13394 (
            .O(N__54722),
            .I(N__54613));
    LocalMux I__13393 (
            .O(N__54719),
            .I(N__54610));
    InMux I__13392 (
            .O(N__54718),
            .I(N__54605));
    InMux I__13391 (
            .O(N__54717),
            .I(N__54605));
    Span4Mux_v I__13390 (
            .O(N__54714),
            .I(N__54600));
    Span4Mux_v I__13389 (
            .O(N__54711),
            .I(N__54600));
    InMux I__13388 (
            .O(N__54710),
            .I(N__54593));
    InMux I__13387 (
            .O(N__54709),
            .I(N__54593));
    InMux I__13386 (
            .O(N__54708),
            .I(N__54593));
    InMux I__13385 (
            .O(N__54707),
            .I(N__54588));
    InMux I__13384 (
            .O(N__54706),
            .I(N__54588));
    InMux I__13383 (
            .O(N__54705),
            .I(N__54585));
    LocalMux I__13382 (
            .O(N__54700),
            .I(N__54580));
    Span4Mux_v I__13381 (
            .O(N__54697),
            .I(N__54580));
    LocalMux I__13380 (
            .O(N__54694),
            .I(N__54577));
    LocalMux I__13379 (
            .O(N__54691),
            .I(N__54566));
    Span4Mux_v I__13378 (
            .O(N__54686),
            .I(N__54566));
    LocalMux I__13377 (
            .O(N__54677),
            .I(N__54566));
    LocalMux I__13376 (
            .O(N__54668),
            .I(N__54566));
    Span4Mux_v I__13375 (
            .O(N__54661),
            .I(N__54566));
    Span4Mux_h I__13374 (
            .O(N__54656),
            .I(N__54563));
    InMux I__13373 (
            .O(N__54655),
            .I(N__54560));
    InMux I__13372 (
            .O(N__54654),
            .I(N__54555));
    LocalMux I__13371 (
            .O(N__54649),
            .I(N__54548));
    LocalMux I__13370 (
            .O(N__54646),
            .I(N__54548));
    Span4Mux_v I__13369 (
            .O(N__54641),
            .I(N__54548));
    Span4Mux_h I__13368 (
            .O(N__54638),
            .I(N__54545));
    InMux I__13367 (
            .O(N__54637),
            .I(N__54538));
    InMux I__13366 (
            .O(N__54636),
            .I(N__54538));
    InMux I__13365 (
            .O(N__54635),
            .I(N__54538));
    Span4Mux_h I__13364 (
            .O(N__54632),
            .I(N__54534));
    LocalMux I__13363 (
            .O(N__54629),
            .I(N__54531));
    LocalMux I__13362 (
            .O(N__54626),
            .I(N__54525));
    Span4Mux_v I__13361 (
            .O(N__54621),
            .I(N__54522));
    LocalMux I__13360 (
            .O(N__54616),
            .I(N__54507));
    LocalMux I__13359 (
            .O(N__54613),
            .I(N__54507));
    Span4Mux_v I__13358 (
            .O(N__54610),
            .I(N__54507));
    LocalMux I__13357 (
            .O(N__54605),
            .I(N__54507));
    Span4Mux_v I__13356 (
            .O(N__54600),
            .I(N__54507));
    LocalMux I__13355 (
            .O(N__54593),
            .I(N__54507));
    LocalMux I__13354 (
            .O(N__54588),
            .I(N__54507));
    LocalMux I__13353 (
            .O(N__54585),
            .I(N__54496));
    Span4Mux_h I__13352 (
            .O(N__54580),
            .I(N__54496));
    Span4Mux_h I__13351 (
            .O(N__54577),
            .I(N__54496));
    Span4Mux_h I__13350 (
            .O(N__54566),
            .I(N__54496));
    Span4Mux_v I__13349 (
            .O(N__54563),
            .I(N__54496));
    LocalMux I__13348 (
            .O(N__54560),
            .I(N__54493));
    InMux I__13347 (
            .O(N__54559),
            .I(N__54488));
    InMux I__13346 (
            .O(N__54558),
            .I(N__54488));
    LocalMux I__13345 (
            .O(N__54555),
            .I(N__54479));
    Span4Mux_v I__13344 (
            .O(N__54548),
            .I(N__54479));
    Span4Mux_h I__13343 (
            .O(N__54545),
            .I(N__54479));
    LocalMux I__13342 (
            .O(N__54538),
            .I(N__54479));
    InMux I__13341 (
            .O(N__54537),
            .I(N__54476));
    Sp12to4 I__13340 (
            .O(N__54534),
            .I(N__54471));
    Span12Mux_s11_v I__13339 (
            .O(N__54531),
            .I(N__54471));
    InMux I__13338 (
            .O(N__54530),
            .I(N__54468));
    InMux I__13337 (
            .O(N__54529),
            .I(N__54463));
    InMux I__13336 (
            .O(N__54528),
            .I(N__54463));
    Span4Mux_v I__13335 (
            .O(N__54525),
            .I(N__54456));
    Span4Mux_h I__13334 (
            .O(N__54522),
            .I(N__54456));
    Span4Mux_v I__13333 (
            .O(N__54507),
            .I(N__54456));
    Span4Mux_v I__13332 (
            .O(N__54496),
            .I(N__54453));
    Span4Mux_v I__13331 (
            .O(N__54493),
            .I(N__54446));
    LocalMux I__13330 (
            .O(N__54488),
            .I(N__54446));
    Span4Mux_v I__13329 (
            .O(N__54479),
            .I(N__54446));
    LocalMux I__13328 (
            .O(N__54476),
            .I(comm_state_3));
    Odrv12 I__13327 (
            .O(N__54471),
            .I(comm_state_3));
    LocalMux I__13326 (
            .O(N__54468),
            .I(comm_state_3));
    LocalMux I__13325 (
            .O(N__54463),
            .I(comm_state_3));
    Odrv4 I__13324 (
            .O(N__54456),
            .I(comm_state_3));
    Odrv4 I__13323 (
            .O(N__54453),
            .I(comm_state_3));
    Odrv4 I__13322 (
            .O(N__54446),
            .I(comm_state_3));
    CEMux I__13321 (
            .O(N__54431),
            .I(N__54428));
    LocalMux I__13320 (
            .O(N__54428),
            .I(N__54425));
    Span4Mux_h I__13319 (
            .O(N__54425),
            .I(N__54422));
    Span4Mux_h I__13318 (
            .O(N__54422),
            .I(N__54419));
    Odrv4 I__13317 (
            .O(N__54419),
            .I(n11377));
    SRMux I__13316 (
            .O(N__54416),
            .I(N__54413));
    LocalMux I__13315 (
            .O(N__54413),
            .I(N__54410));
    Odrv4 I__13314 (
            .O(N__54410),
            .I(\comm_spi.data_tx_7__N_770 ));
    InMux I__13313 (
            .O(N__54407),
            .I(N__54404));
    LocalMux I__13312 (
            .O(N__54404),
            .I(N__54401));
    Sp12to4 I__13311 (
            .O(N__54401),
            .I(N__54398));
    Odrv12 I__13310 (
            .O(N__54398),
            .I(comm_buf_5_6));
    InMux I__13309 (
            .O(N__54395),
            .I(N__54392));
    LocalMux I__13308 (
            .O(N__54392),
            .I(N__54389));
    Span12Mux_h I__13307 (
            .O(N__54389),
            .I(N__54386));
    Odrv12 I__13306 (
            .O(N__54386),
            .I(comm_buf_4_6));
    CascadeMux I__13305 (
            .O(N__54383),
            .I(N__54375));
    InMux I__13304 (
            .O(N__54382),
            .I(N__54356));
    InMux I__13303 (
            .O(N__54381),
            .I(N__54356));
    InMux I__13302 (
            .O(N__54380),
            .I(N__54356));
    InMux I__13301 (
            .O(N__54379),
            .I(N__54356));
    InMux I__13300 (
            .O(N__54378),
            .I(N__54356));
    InMux I__13299 (
            .O(N__54375),
            .I(N__54353));
    CascadeMux I__13298 (
            .O(N__54374),
            .I(N__54348));
    InMux I__13297 (
            .O(N__54373),
            .I(N__54332));
    InMux I__13296 (
            .O(N__54372),
            .I(N__54332));
    InMux I__13295 (
            .O(N__54371),
            .I(N__54332));
    InMux I__13294 (
            .O(N__54370),
            .I(N__54332));
    InMux I__13293 (
            .O(N__54369),
            .I(N__54332));
    InMux I__13292 (
            .O(N__54368),
            .I(N__54324));
    CascadeMux I__13291 (
            .O(N__54367),
            .I(N__54321));
    LocalMux I__13290 (
            .O(N__54356),
            .I(N__54315));
    LocalMux I__13289 (
            .O(N__54353),
            .I(N__54312));
    InMux I__13288 (
            .O(N__54352),
            .I(N__54309));
    InMux I__13287 (
            .O(N__54351),
            .I(N__54303));
    InMux I__13286 (
            .O(N__54348),
            .I(N__54303));
    InMux I__13285 (
            .O(N__54347),
            .I(N__54298));
    InMux I__13284 (
            .O(N__54346),
            .I(N__54298));
    InMux I__13283 (
            .O(N__54345),
            .I(N__54291));
    InMux I__13282 (
            .O(N__54344),
            .I(N__54291));
    InMux I__13281 (
            .O(N__54343),
            .I(N__54291));
    LocalMux I__13280 (
            .O(N__54332),
            .I(N__54284));
    InMux I__13279 (
            .O(N__54331),
            .I(N__54273));
    InMux I__13278 (
            .O(N__54330),
            .I(N__54273));
    InMux I__13277 (
            .O(N__54329),
            .I(N__54273));
    InMux I__13276 (
            .O(N__54328),
            .I(N__54273));
    InMux I__13275 (
            .O(N__54327),
            .I(N__54273));
    LocalMux I__13274 (
            .O(N__54324),
            .I(N__54266));
    InMux I__13273 (
            .O(N__54321),
            .I(N__54257));
    InMux I__13272 (
            .O(N__54320),
            .I(N__54257));
    InMux I__13271 (
            .O(N__54319),
            .I(N__54257));
    InMux I__13270 (
            .O(N__54318),
            .I(N__54257));
    Span4Mux_v I__13269 (
            .O(N__54315),
            .I(N__54254));
    Span4Mux_h I__13268 (
            .O(N__54312),
            .I(N__54249));
    LocalMux I__13267 (
            .O(N__54309),
            .I(N__54249));
    InMux I__13266 (
            .O(N__54308),
            .I(N__54246));
    LocalMux I__13265 (
            .O(N__54303),
            .I(N__54239));
    LocalMux I__13264 (
            .O(N__54298),
            .I(N__54239));
    LocalMux I__13263 (
            .O(N__54291),
            .I(N__54239));
    InMux I__13262 (
            .O(N__54290),
            .I(N__54230));
    InMux I__13261 (
            .O(N__54289),
            .I(N__54230));
    InMux I__13260 (
            .O(N__54288),
            .I(N__54230));
    InMux I__13259 (
            .O(N__54287),
            .I(N__54230));
    Span4Mux_v I__13258 (
            .O(N__54284),
            .I(N__54225));
    LocalMux I__13257 (
            .O(N__54273),
            .I(N__54225));
    InMux I__13256 (
            .O(N__54272),
            .I(N__54216));
    InMux I__13255 (
            .O(N__54271),
            .I(N__54216));
    InMux I__13254 (
            .O(N__54270),
            .I(N__54216));
    InMux I__13253 (
            .O(N__54269),
            .I(N__54216));
    Span4Mux_v I__13252 (
            .O(N__54266),
            .I(N__54207));
    LocalMux I__13251 (
            .O(N__54257),
            .I(N__54207));
    Span4Mux_h I__13250 (
            .O(N__54254),
            .I(N__54207));
    Span4Mux_v I__13249 (
            .O(N__54249),
            .I(N__54207));
    LocalMux I__13248 (
            .O(N__54246),
            .I(N__54204));
    Odrv4 I__13247 (
            .O(N__54239),
            .I(comm_index_0));
    LocalMux I__13246 (
            .O(N__54230),
            .I(comm_index_0));
    Odrv4 I__13245 (
            .O(N__54225),
            .I(comm_index_0));
    LocalMux I__13244 (
            .O(N__54216),
            .I(comm_index_0));
    Odrv4 I__13243 (
            .O(N__54207),
            .I(comm_index_0));
    Odrv12 I__13242 (
            .O(N__54204),
            .I(comm_index_0));
    InMux I__13241 (
            .O(N__54191),
            .I(N__54188));
    LocalMux I__13240 (
            .O(N__54188),
            .I(N__54185));
    Span4Mux_h I__13239 (
            .O(N__54185),
            .I(N__54182));
    Odrv4 I__13238 (
            .O(N__54182),
            .I(n4_adj_1585));
    InMux I__13237 (
            .O(N__54179),
            .I(N__54151));
    InMux I__13236 (
            .O(N__54178),
            .I(N__54151));
    InMux I__13235 (
            .O(N__54177),
            .I(N__54151));
    InMux I__13234 (
            .O(N__54176),
            .I(N__54151));
    InMux I__13233 (
            .O(N__54175),
            .I(N__54151));
    InMux I__13232 (
            .O(N__54174),
            .I(N__54151));
    CascadeMux I__13231 (
            .O(N__54173),
            .I(N__54146));
    CascadeMux I__13230 (
            .O(N__54172),
            .I(N__54142));
    InMux I__13229 (
            .O(N__54171),
            .I(N__54133));
    InMux I__13228 (
            .O(N__54170),
            .I(N__54130));
    InMux I__13227 (
            .O(N__54169),
            .I(N__54125));
    InMux I__13226 (
            .O(N__54168),
            .I(N__54113));
    InMux I__13225 (
            .O(N__54167),
            .I(N__54113));
    InMux I__13224 (
            .O(N__54166),
            .I(N__54113));
    InMux I__13223 (
            .O(N__54165),
            .I(N__54113));
    InMux I__13222 (
            .O(N__54164),
            .I(N__54113));
    LocalMux I__13221 (
            .O(N__54151),
            .I(N__54110));
    InMux I__13220 (
            .O(N__54150),
            .I(N__54107));
    InMux I__13219 (
            .O(N__54149),
            .I(N__54095));
    InMux I__13218 (
            .O(N__54146),
            .I(N__54095));
    InMux I__13217 (
            .O(N__54145),
            .I(N__54095));
    InMux I__13216 (
            .O(N__54142),
            .I(N__54095));
    InMux I__13215 (
            .O(N__54141),
            .I(N__54095));
    CascadeMux I__13214 (
            .O(N__54140),
            .I(N__54092));
    InMux I__13213 (
            .O(N__54139),
            .I(N__54064));
    InMux I__13212 (
            .O(N__54138),
            .I(N__54057));
    InMux I__13211 (
            .O(N__54137),
            .I(N__54057));
    InMux I__13210 (
            .O(N__54136),
            .I(N__54057));
    LocalMux I__13209 (
            .O(N__54133),
            .I(N__54048));
    LocalMux I__13208 (
            .O(N__54130),
            .I(N__54045));
    InMux I__13207 (
            .O(N__54129),
            .I(N__54040));
    InMux I__13206 (
            .O(N__54128),
            .I(N__54040));
    LocalMux I__13205 (
            .O(N__54125),
            .I(N__54037));
    InMux I__13204 (
            .O(N__54124),
            .I(N__54023));
    LocalMux I__13203 (
            .O(N__54113),
            .I(N__54015));
    Span4Mux_h I__13202 (
            .O(N__54110),
            .I(N__54015));
    LocalMux I__13201 (
            .O(N__54107),
            .I(N__54015));
    InMux I__13200 (
            .O(N__54106),
            .I(N__54012));
    LocalMux I__13199 (
            .O(N__54095),
            .I(N__54009));
    InMux I__13198 (
            .O(N__54092),
            .I(N__53998));
    InMux I__13197 (
            .O(N__54091),
            .I(N__53998));
    InMux I__13196 (
            .O(N__54090),
            .I(N__53998));
    InMux I__13195 (
            .O(N__54089),
            .I(N__53991));
    InMux I__13194 (
            .O(N__54088),
            .I(N__53988));
    InMux I__13193 (
            .O(N__54087),
            .I(N__53985));
    InMux I__13192 (
            .O(N__54086),
            .I(N__53982));
    InMux I__13191 (
            .O(N__54085),
            .I(N__53965));
    InMux I__13190 (
            .O(N__54084),
            .I(N__53965));
    InMux I__13189 (
            .O(N__54083),
            .I(N__53965));
    InMux I__13188 (
            .O(N__54082),
            .I(N__53965));
    InMux I__13187 (
            .O(N__54081),
            .I(N__53965));
    InMux I__13186 (
            .O(N__54080),
            .I(N__53965));
    InMux I__13185 (
            .O(N__54079),
            .I(N__53965));
    InMux I__13184 (
            .O(N__54078),
            .I(N__53965));
    InMux I__13183 (
            .O(N__54077),
            .I(N__53960));
    InMux I__13182 (
            .O(N__54076),
            .I(N__53952));
    InMux I__13181 (
            .O(N__54075),
            .I(N__53947));
    InMux I__13180 (
            .O(N__54074),
            .I(N__53930));
    InMux I__13179 (
            .O(N__54073),
            .I(N__53930));
    InMux I__13178 (
            .O(N__54072),
            .I(N__53930));
    InMux I__13177 (
            .O(N__54071),
            .I(N__53930));
    InMux I__13176 (
            .O(N__54070),
            .I(N__53930));
    InMux I__13175 (
            .O(N__54069),
            .I(N__53930));
    InMux I__13174 (
            .O(N__54068),
            .I(N__53930));
    InMux I__13173 (
            .O(N__54067),
            .I(N__53930));
    LocalMux I__13172 (
            .O(N__54064),
            .I(N__53925));
    LocalMux I__13171 (
            .O(N__54057),
            .I(N__53925));
    CascadeMux I__13170 (
            .O(N__54056),
            .I(N__53922));
    InMux I__13169 (
            .O(N__54055),
            .I(N__53918));
    InMux I__13168 (
            .O(N__54054),
            .I(N__53914));
    InMux I__13167 (
            .O(N__54053),
            .I(N__53911));
    InMux I__13166 (
            .O(N__54052),
            .I(N__53908));
    InMux I__13165 (
            .O(N__54051),
            .I(N__53905));
    Span4Mux_h I__13164 (
            .O(N__54048),
            .I(N__53902));
    Span4Mux_h I__13163 (
            .O(N__54045),
            .I(N__53895));
    LocalMux I__13162 (
            .O(N__54040),
            .I(N__53895));
    Span4Mux_h I__13161 (
            .O(N__54037),
            .I(N__53895));
    InMux I__13160 (
            .O(N__54036),
            .I(N__53892));
    InMux I__13159 (
            .O(N__54035),
            .I(N__53885));
    InMux I__13158 (
            .O(N__54034),
            .I(N__53885));
    InMux I__13157 (
            .O(N__54033),
            .I(N__53885));
    InMux I__13156 (
            .O(N__54032),
            .I(N__53878));
    InMux I__13155 (
            .O(N__54031),
            .I(N__53878));
    InMux I__13154 (
            .O(N__54030),
            .I(N__53878));
    InMux I__13153 (
            .O(N__54029),
            .I(N__53875));
    InMux I__13152 (
            .O(N__54028),
            .I(N__53872));
    InMux I__13151 (
            .O(N__54027),
            .I(N__53869));
    InMux I__13150 (
            .O(N__54026),
            .I(N__53866));
    LocalMux I__13149 (
            .O(N__54023),
            .I(N__53863));
    InMux I__13148 (
            .O(N__54022),
            .I(N__53859));
    Span4Mux_v I__13147 (
            .O(N__54015),
            .I(N__53856));
    LocalMux I__13146 (
            .O(N__54012),
            .I(N__53851));
    Span4Mux_v I__13145 (
            .O(N__54009),
            .I(N__53851));
    InMux I__13144 (
            .O(N__54008),
            .I(N__53844));
    InMux I__13143 (
            .O(N__54007),
            .I(N__53844));
    InMux I__13142 (
            .O(N__54006),
            .I(N__53844));
    InMux I__13141 (
            .O(N__54005),
            .I(N__53839));
    LocalMux I__13140 (
            .O(N__53998),
            .I(N__53836));
    InMux I__13139 (
            .O(N__53997),
            .I(N__53829));
    InMux I__13138 (
            .O(N__53996),
            .I(N__53829));
    InMux I__13137 (
            .O(N__53995),
            .I(N__53829));
    InMux I__13136 (
            .O(N__53994),
            .I(N__53826));
    LocalMux I__13135 (
            .O(N__53991),
            .I(N__53817));
    LocalMux I__13134 (
            .O(N__53988),
            .I(N__53817));
    LocalMux I__13133 (
            .O(N__53985),
            .I(N__53817));
    LocalMux I__13132 (
            .O(N__53982),
            .I(N__53817));
    LocalMux I__13131 (
            .O(N__53965),
            .I(N__53814));
    InMux I__13130 (
            .O(N__53964),
            .I(N__53807));
    InMux I__13129 (
            .O(N__53963),
            .I(N__53807));
    LocalMux I__13128 (
            .O(N__53960),
            .I(N__53801));
    InMux I__13127 (
            .O(N__53959),
            .I(N__53794));
    InMux I__13126 (
            .O(N__53958),
            .I(N__53794));
    InMux I__13125 (
            .O(N__53957),
            .I(N__53794));
    InMux I__13124 (
            .O(N__53956),
            .I(N__53789));
    InMux I__13123 (
            .O(N__53955),
            .I(N__53789));
    LocalMux I__13122 (
            .O(N__53952),
            .I(N__53783));
    InMux I__13121 (
            .O(N__53951),
            .I(N__53778));
    InMux I__13120 (
            .O(N__53950),
            .I(N__53778));
    LocalMux I__13119 (
            .O(N__53947),
            .I(N__53775));
    LocalMux I__13118 (
            .O(N__53930),
            .I(N__53765));
    Span4Mux_v I__13117 (
            .O(N__53925),
            .I(N__53765));
    InMux I__13116 (
            .O(N__53922),
            .I(N__53760));
    InMux I__13115 (
            .O(N__53921),
            .I(N__53760));
    LocalMux I__13114 (
            .O(N__53918),
            .I(N__53757));
    InMux I__13113 (
            .O(N__53917),
            .I(N__53754));
    LocalMux I__13112 (
            .O(N__53914),
            .I(N__53741));
    LocalMux I__13111 (
            .O(N__53911),
            .I(N__53741));
    LocalMux I__13110 (
            .O(N__53908),
            .I(N__53741));
    LocalMux I__13109 (
            .O(N__53905),
            .I(N__53741));
    Span4Mux_h I__13108 (
            .O(N__53902),
            .I(N__53741));
    Span4Mux_v I__13107 (
            .O(N__53895),
            .I(N__53741));
    LocalMux I__13106 (
            .O(N__53892),
            .I(N__53732));
    LocalMux I__13105 (
            .O(N__53885),
            .I(N__53732));
    LocalMux I__13104 (
            .O(N__53878),
            .I(N__53732));
    LocalMux I__13103 (
            .O(N__53875),
            .I(N__53732));
    LocalMux I__13102 (
            .O(N__53872),
            .I(N__53729));
    LocalMux I__13101 (
            .O(N__53869),
            .I(N__53722));
    LocalMux I__13100 (
            .O(N__53866),
            .I(N__53722));
    Span4Mux_h I__13099 (
            .O(N__53863),
            .I(N__53722));
    InMux I__13098 (
            .O(N__53862),
            .I(N__53719));
    LocalMux I__13097 (
            .O(N__53859),
            .I(N__53710));
    Span4Mux_h I__13096 (
            .O(N__53856),
            .I(N__53710));
    Span4Mux_h I__13095 (
            .O(N__53851),
            .I(N__53710));
    LocalMux I__13094 (
            .O(N__53844),
            .I(N__53710));
    InMux I__13093 (
            .O(N__53843),
            .I(N__53705));
    InMux I__13092 (
            .O(N__53842),
            .I(N__53705));
    LocalMux I__13091 (
            .O(N__53839),
            .I(N__53698));
    Sp12to4 I__13090 (
            .O(N__53836),
            .I(N__53698));
    LocalMux I__13089 (
            .O(N__53829),
            .I(N__53698));
    LocalMux I__13088 (
            .O(N__53826),
            .I(N__53691));
    Span4Mux_v I__13087 (
            .O(N__53817),
            .I(N__53691));
    Span4Mux_v I__13086 (
            .O(N__53814),
            .I(N__53691));
    InMux I__13085 (
            .O(N__53813),
            .I(N__53686));
    InMux I__13084 (
            .O(N__53812),
            .I(N__53686));
    LocalMux I__13083 (
            .O(N__53807),
            .I(N__53683));
    InMux I__13082 (
            .O(N__53806),
            .I(N__53676));
    InMux I__13081 (
            .O(N__53805),
            .I(N__53676));
    InMux I__13080 (
            .O(N__53804),
            .I(N__53676));
    Span4Mux_h I__13079 (
            .O(N__53801),
            .I(N__53669));
    LocalMux I__13078 (
            .O(N__53794),
            .I(N__53669));
    LocalMux I__13077 (
            .O(N__53789),
            .I(N__53669));
    InMux I__13076 (
            .O(N__53788),
            .I(N__53662));
    InMux I__13075 (
            .O(N__53787),
            .I(N__53662));
    InMux I__13074 (
            .O(N__53786),
            .I(N__53662));
    Span4Mux_v I__13073 (
            .O(N__53783),
            .I(N__53655));
    LocalMux I__13072 (
            .O(N__53778),
            .I(N__53655));
    Span4Mux_h I__13071 (
            .O(N__53775),
            .I(N__53655));
    InMux I__13070 (
            .O(N__53774),
            .I(N__53650));
    InMux I__13069 (
            .O(N__53773),
            .I(N__53650));
    InMux I__13068 (
            .O(N__53772),
            .I(N__53643));
    InMux I__13067 (
            .O(N__53771),
            .I(N__53643));
    InMux I__13066 (
            .O(N__53770),
            .I(N__53643));
    Span4Mux_h I__13065 (
            .O(N__53765),
            .I(N__53628));
    LocalMux I__13064 (
            .O(N__53760),
            .I(N__53628));
    Span4Mux_v I__13063 (
            .O(N__53757),
            .I(N__53628));
    LocalMux I__13062 (
            .O(N__53754),
            .I(N__53628));
    Span4Mux_v I__13061 (
            .O(N__53741),
            .I(N__53628));
    Span4Mux_v I__13060 (
            .O(N__53732),
            .I(N__53628));
    Span4Mux_v I__13059 (
            .O(N__53729),
            .I(N__53628));
    Span4Mux_v I__13058 (
            .O(N__53722),
            .I(N__53621));
    LocalMux I__13057 (
            .O(N__53719),
            .I(N__53621));
    Span4Mux_h I__13056 (
            .O(N__53710),
            .I(N__53621));
    LocalMux I__13055 (
            .O(N__53705),
            .I(N__53616));
    Span12Mux_v I__13054 (
            .O(N__53698),
            .I(N__53616));
    Odrv4 I__13053 (
            .O(N__53691),
            .I(comm_state_1));
    LocalMux I__13052 (
            .O(N__53686),
            .I(comm_state_1));
    Odrv4 I__13051 (
            .O(N__53683),
            .I(comm_state_1));
    LocalMux I__13050 (
            .O(N__53676),
            .I(comm_state_1));
    Odrv4 I__13049 (
            .O(N__53669),
            .I(comm_state_1));
    LocalMux I__13048 (
            .O(N__53662),
            .I(comm_state_1));
    Odrv4 I__13047 (
            .O(N__53655),
            .I(comm_state_1));
    LocalMux I__13046 (
            .O(N__53650),
            .I(comm_state_1));
    LocalMux I__13045 (
            .O(N__53643),
            .I(comm_state_1));
    Odrv4 I__13044 (
            .O(N__53628),
            .I(comm_state_1));
    Odrv4 I__13043 (
            .O(N__53621),
            .I(comm_state_1));
    Odrv12 I__13042 (
            .O(N__53616),
            .I(comm_state_1));
    InMux I__13041 (
            .O(N__53591),
            .I(N__53583));
    InMux I__13040 (
            .O(N__53590),
            .I(N__53572));
    InMux I__13039 (
            .O(N__53589),
            .I(N__53572));
    InMux I__13038 (
            .O(N__53588),
            .I(N__53572));
    InMux I__13037 (
            .O(N__53587),
            .I(N__53572));
    InMux I__13036 (
            .O(N__53586),
            .I(N__53569));
    LocalMux I__13035 (
            .O(N__53583),
            .I(N__53558));
    InMux I__13034 (
            .O(N__53582),
            .I(N__53555));
    InMux I__13033 (
            .O(N__53581),
            .I(N__53550));
    LocalMux I__13032 (
            .O(N__53572),
            .I(N__53545));
    LocalMux I__13031 (
            .O(N__53569),
            .I(N__53542));
    InMux I__13030 (
            .O(N__53568),
            .I(N__53539));
    InMux I__13029 (
            .O(N__53567),
            .I(N__53534));
    InMux I__13028 (
            .O(N__53566),
            .I(N__53531));
    InMux I__13027 (
            .O(N__53565),
            .I(N__53524));
    InMux I__13026 (
            .O(N__53564),
            .I(N__53524));
    InMux I__13025 (
            .O(N__53563),
            .I(N__53524));
    InMux I__13024 (
            .O(N__53562),
            .I(N__53521));
    InMux I__13023 (
            .O(N__53561),
            .I(N__53513));
    Span4Mux_v I__13022 (
            .O(N__53558),
            .I(N__53510));
    LocalMux I__13021 (
            .O(N__53555),
            .I(N__53507));
    InMux I__13020 (
            .O(N__53554),
            .I(N__53498));
    InMux I__13019 (
            .O(N__53553),
            .I(N__53498));
    LocalMux I__13018 (
            .O(N__53550),
            .I(N__53492));
    InMux I__13017 (
            .O(N__53549),
            .I(N__53489));
    InMux I__13016 (
            .O(N__53548),
            .I(N__53486));
    Span4Mux_v I__13015 (
            .O(N__53545),
            .I(N__53479));
    Span4Mux_v I__13014 (
            .O(N__53542),
            .I(N__53479));
    LocalMux I__13013 (
            .O(N__53539),
            .I(N__53479));
    InMux I__13012 (
            .O(N__53538),
            .I(N__53474));
    InMux I__13011 (
            .O(N__53537),
            .I(N__53474));
    LocalMux I__13010 (
            .O(N__53534),
            .I(N__53471));
    LocalMux I__13009 (
            .O(N__53531),
            .I(N__53468));
    LocalMux I__13008 (
            .O(N__53524),
            .I(N__53460));
    LocalMux I__13007 (
            .O(N__53521),
            .I(N__53460));
    InMux I__13006 (
            .O(N__53520),
            .I(N__53455));
    InMux I__13005 (
            .O(N__53519),
            .I(N__53455));
    InMux I__13004 (
            .O(N__53518),
            .I(N__53448));
    InMux I__13003 (
            .O(N__53517),
            .I(N__53448));
    InMux I__13002 (
            .O(N__53516),
            .I(N__53448));
    LocalMux I__13001 (
            .O(N__53513),
            .I(N__53443));
    Span4Mux_h I__13000 (
            .O(N__53510),
            .I(N__53443));
    Span4Mux_v I__12999 (
            .O(N__53507),
            .I(N__53440));
    InMux I__12998 (
            .O(N__53506),
            .I(N__53435));
    InMux I__12997 (
            .O(N__53505),
            .I(N__53435));
    InMux I__12996 (
            .O(N__53504),
            .I(N__53430));
    InMux I__12995 (
            .O(N__53503),
            .I(N__53430));
    LocalMux I__12994 (
            .O(N__53498),
            .I(N__53427));
    InMux I__12993 (
            .O(N__53497),
            .I(N__53420));
    InMux I__12992 (
            .O(N__53496),
            .I(N__53420));
    InMux I__12991 (
            .O(N__53495),
            .I(N__53420));
    Span4Mux_v I__12990 (
            .O(N__53492),
            .I(N__53417));
    LocalMux I__12989 (
            .O(N__53489),
            .I(N__53414));
    LocalMux I__12988 (
            .O(N__53486),
            .I(N__53411));
    Span4Mux_v I__12987 (
            .O(N__53479),
            .I(N__53408));
    LocalMux I__12986 (
            .O(N__53474),
            .I(N__53405));
    Span4Mux_v I__12985 (
            .O(N__53471),
            .I(N__53400));
    Span4Mux_v I__12984 (
            .O(N__53468),
            .I(N__53400));
    InMux I__12983 (
            .O(N__53467),
            .I(N__53393));
    InMux I__12982 (
            .O(N__53466),
            .I(N__53393));
    InMux I__12981 (
            .O(N__53465),
            .I(N__53393));
    Span4Mux_h I__12980 (
            .O(N__53460),
            .I(N__53386));
    LocalMux I__12979 (
            .O(N__53455),
            .I(N__53386));
    LocalMux I__12978 (
            .O(N__53448),
            .I(N__53386));
    Span4Mux_h I__12977 (
            .O(N__53443),
            .I(N__53383));
    Span4Mux_v I__12976 (
            .O(N__53440),
            .I(N__53364));
    LocalMux I__12975 (
            .O(N__53435),
            .I(N__53364));
    LocalMux I__12974 (
            .O(N__53430),
            .I(N__53364));
    Span4Mux_v I__12973 (
            .O(N__53427),
            .I(N__53364));
    LocalMux I__12972 (
            .O(N__53420),
            .I(N__53364));
    Span4Mux_v I__12971 (
            .O(N__53417),
            .I(N__53364));
    Span4Mux_v I__12970 (
            .O(N__53414),
            .I(N__53364));
    Span4Mux_v I__12969 (
            .O(N__53411),
            .I(N__53364));
    Span4Mux_h I__12968 (
            .O(N__53408),
            .I(N__53364));
    Odrv4 I__12967 (
            .O(N__53405),
            .I(comm_state_0));
    Odrv4 I__12966 (
            .O(N__53400),
            .I(comm_state_0));
    LocalMux I__12965 (
            .O(N__53393),
            .I(comm_state_0));
    Odrv4 I__12964 (
            .O(N__53386),
            .I(comm_state_0));
    Odrv4 I__12963 (
            .O(N__53383),
            .I(comm_state_0));
    Odrv4 I__12962 (
            .O(N__53364),
            .I(comm_state_0));
    CascadeMux I__12961 (
            .O(N__53351),
            .I(N__53347));
    InMux I__12960 (
            .O(N__53350),
            .I(N__53341));
    InMux I__12959 (
            .O(N__53347),
            .I(N__53341));
    InMux I__12958 (
            .O(N__53346),
            .I(N__53338));
    LocalMux I__12957 (
            .O(N__53341),
            .I(N__53333));
    LocalMux I__12956 (
            .O(N__53338),
            .I(N__53333));
    Span4Mux_h I__12955 (
            .O(N__53333),
            .I(N__53330));
    Odrv4 I__12954 (
            .O(N__53330),
            .I(n9270));
    InMux I__12953 (
            .O(N__53327),
            .I(N__53321));
    InMux I__12952 (
            .O(N__53326),
            .I(N__53318));
    InMux I__12951 (
            .O(N__53325),
            .I(N__53313));
    InMux I__12950 (
            .O(N__53324),
            .I(N__53313));
    LocalMux I__12949 (
            .O(N__53321),
            .I(\comm_spi.n22670 ));
    LocalMux I__12948 (
            .O(N__53318),
            .I(\comm_spi.n22670 ));
    LocalMux I__12947 (
            .O(N__53313),
            .I(\comm_spi.n22670 ));
    InMux I__12946 (
            .O(N__53306),
            .I(N__53303));
    LocalMux I__12945 (
            .O(N__53303),
            .I(\comm_spi.n14631 ));
    InMux I__12944 (
            .O(N__53300),
            .I(N__53297));
    LocalMux I__12943 (
            .O(N__53297),
            .I(N__53292));
    InMux I__12942 (
            .O(N__53296),
            .I(N__53289));
    InMux I__12941 (
            .O(N__53295),
            .I(N__53286));
    Odrv4 I__12940 (
            .O(N__53292),
            .I(\comm_spi.n14616 ));
    LocalMux I__12939 (
            .O(N__53289),
            .I(\comm_spi.n14616 ));
    LocalMux I__12938 (
            .O(N__53286),
            .I(\comm_spi.n14616 ));
    InMux I__12937 (
            .O(N__53279),
            .I(N__53274));
    InMux I__12936 (
            .O(N__53278),
            .I(N__53271));
    InMux I__12935 (
            .O(N__53277),
            .I(N__53268));
    LocalMux I__12934 (
            .O(N__53274),
            .I(N__53265));
    LocalMux I__12933 (
            .O(N__53271),
            .I(N__53260));
    LocalMux I__12932 (
            .O(N__53268),
            .I(N__53260));
    Odrv4 I__12931 (
            .O(N__53265),
            .I(\comm_spi.n14617 ));
    Odrv4 I__12930 (
            .O(N__53260),
            .I(\comm_spi.n14617 ));
    CascadeMux I__12929 (
            .O(N__53255),
            .I(N__53251));
    InMux I__12928 (
            .O(N__53254),
            .I(N__53247));
    InMux I__12927 (
            .O(N__53251),
            .I(N__53242));
    InMux I__12926 (
            .O(N__53250),
            .I(N__53242));
    LocalMux I__12925 (
            .O(N__53247),
            .I(cmd_rdadctmp_19_adj_1431));
    LocalMux I__12924 (
            .O(N__53242),
            .I(cmd_rdadctmp_19_adj_1431));
    InMux I__12923 (
            .O(N__53237),
            .I(N__53234));
    LocalMux I__12922 (
            .O(N__53234),
            .I(N__53231));
    Span4Mux_v I__12921 (
            .O(N__53231),
            .I(N__53226));
    InMux I__12920 (
            .O(N__53230),
            .I(N__53223));
    InMux I__12919 (
            .O(N__53229),
            .I(N__53220));
    Span4Mux_h I__12918 (
            .O(N__53226),
            .I(N__53217));
    LocalMux I__12917 (
            .O(N__53223),
            .I(N__53214));
    LocalMux I__12916 (
            .O(N__53220),
            .I(buf_adcdata_iac_11));
    Odrv4 I__12915 (
            .O(N__53217),
            .I(buf_adcdata_iac_11));
    Odrv12 I__12914 (
            .O(N__53214),
            .I(buf_adcdata_iac_11));
    InMux I__12913 (
            .O(N__53207),
            .I(N__53201));
    InMux I__12912 (
            .O(N__53206),
            .I(N__53201));
    LocalMux I__12911 (
            .O(N__53201),
            .I(N__53195));
    InMux I__12910 (
            .O(N__53200),
            .I(N__53192));
    InMux I__12909 (
            .O(N__53199),
            .I(N__53189));
    InMux I__12908 (
            .O(N__53198),
            .I(N__53186));
    Span4Mux_h I__12907 (
            .O(N__53195),
            .I(N__53180));
    LocalMux I__12906 (
            .O(N__53192),
            .I(N__53172));
    LocalMux I__12905 (
            .O(N__53189),
            .I(N__53167));
    LocalMux I__12904 (
            .O(N__53186),
            .I(N__53167));
    InMux I__12903 (
            .O(N__53185),
            .I(N__53163));
    InMux I__12902 (
            .O(N__53184),
            .I(N__53160));
    InMux I__12901 (
            .O(N__53183),
            .I(N__53157));
    Span4Mux_h I__12900 (
            .O(N__53180),
            .I(N__53153));
    InMux I__12899 (
            .O(N__53179),
            .I(N__53146));
    InMux I__12898 (
            .O(N__53178),
            .I(N__53146));
    InMux I__12897 (
            .O(N__53177),
            .I(N__53146));
    InMux I__12896 (
            .O(N__53176),
            .I(N__53143));
    InMux I__12895 (
            .O(N__53175),
            .I(N__53140));
    Span4Mux_h I__12894 (
            .O(N__53172),
            .I(N__53135));
    Span4Mux_v I__12893 (
            .O(N__53167),
            .I(N__53135));
    InMux I__12892 (
            .O(N__53166),
            .I(N__53132));
    LocalMux I__12891 (
            .O(N__53163),
            .I(N__53124));
    LocalMux I__12890 (
            .O(N__53160),
            .I(N__53121));
    LocalMux I__12889 (
            .O(N__53157),
            .I(N__53118));
    CascadeMux I__12888 (
            .O(N__53156),
            .I(N__53113));
    Sp12to4 I__12887 (
            .O(N__53153),
            .I(N__53110));
    LocalMux I__12886 (
            .O(N__53146),
            .I(N__53105));
    LocalMux I__12885 (
            .O(N__53143),
            .I(N__53105));
    LocalMux I__12884 (
            .O(N__53140),
            .I(N__53102));
    Span4Mux_v I__12883 (
            .O(N__53135),
            .I(N__53097));
    LocalMux I__12882 (
            .O(N__53132),
            .I(N__53097));
    InMux I__12881 (
            .O(N__53131),
            .I(N__53092));
    InMux I__12880 (
            .O(N__53130),
            .I(N__53092));
    InMux I__12879 (
            .O(N__53129),
            .I(N__53085));
    InMux I__12878 (
            .O(N__53128),
            .I(N__53085));
    InMux I__12877 (
            .O(N__53127),
            .I(N__53085));
    Span4Mux_v I__12876 (
            .O(N__53124),
            .I(N__53080));
    Span4Mux_v I__12875 (
            .O(N__53121),
            .I(N__53080));
    Span4Mux_v I__12874 (
            .O(N__53118),
            .I(N__53077));
    InMux I__12873 (
            .O(N__53117),
            .I(N__53070));
    InMux I__12872 (
            .O(N__53116),
            .I(N__53070));
    InMux I__12871 (
            .O(N__53113),
            .I(N__53070));
    Span12Mux_v I__12870 (
            .O(N__53110),
            .I(N__53063));
    Span12Mux_v I__12869 (
            .O(N__53105),
            .I(N__53063));
    Span4Mux_h I__12868 (
            .O(N__53102),
            .I(N__53060));
    Span4Mux_v I__12867 (
            .O(N__53097),
            .I(N__53053));
    LocalMux I__12866 (
            .O(N__53092),
            .I(N__53053));
    LocalMux I__12865 (
            .O(N__53085),
            .I(N__53053));
    Span4Mux_v I__12864 (
            .O(N__53080),
            .I(N__53050));
    Span4Mux_v I__12863 (
            .O(N__53077),
            .I(N__53047));
    LocalMux I__12862 (
            .O(N__53070),
            .I(N__53044));
    InMux I__12861 (
            .O(N__53069),
            .I(N__53039));
    InMux I__12860 (
            .O(N__53068),
            .I(N__53039));
    Span12Mux_h I__12859 (
            .O(N__53063),
            .I(N__53036));
    Span4Mux_h I__12858 (
            .O(N__53060),
            .I(N__53033));
    Span4Mux_h I__12857 (
            .O(N__53053),
            .I(N__53030));
    Span4Mux_v I__12856 (
            .O(N__53050),
            .I(N__53021));
    Span4Mux_h I__12855 (
            .O(N__53047),
            .I(N__53021));
    Span4Mux_h I__12854 (
            .O(N__53044),
            .I(N__53021));
    LocalMux I__12853 (
            .O(N__53039),
            .I(N__53021));
    Odrv12 I__12852 (
            .O(N__53036),
            .I(n20584));
    Odrv4 I__12851 (
            .O(N__53033),
            .I(n20584));
    Odrv4 I__12850 (
            .O(N__53030),
            .I(n20584));
    Odrv4 I__12849 (
            .O(N__53021),
            .I(n20584));
    InMux I__12848 (
            .O(N__53012),
            .I(N__53008));
    InMux I__12847 (
            .O(N__53011),
            .I(N__52986));
    LocalMux I__12846 (
            .O(N__53008),
            .I(N__52983));
    InMux I__12845 (
            .O(N__53007),
            .I(N__52970));
    InMux I__12844 (
            .O(N__53006),
            .I(N__52970));
    InMux I__12843 (
            .O(N__53005),
            .I(N__52970));
    InMux I__12842 (
            .O(N__53004),
            .I(N__52970));
    InMux I__12841 (
            .O(N__53003),
            .I(N__52970));
    InMux I__12840 (
            .O(N__53002),
            .I(N__52970));
    CascadeMux I__12839 (
            .O(N__53001),
            .I(N__52967));
    InMux I__12838 (
            .O(N__53000),
            .I(N__52960));
    InMux I__12837 (
            .O(N__52999),
            .I(N__52960));
    InMux I__12836 (
            .O(N__52998),
            .I(N__52960));
    CascadeMux I__12835 (
            .O(N__52997),
            .I(N__52955));
    InMux I__12834 (
            .O(N__52996),
            .I(N__52948));
    InMux I__12833 (
            .O(N__52995),
            .I(N__52945));
    InMux I__12832 (
            .O(N__52994),
            .I(N__52942));
    InMux I__12831 (
            .O(N__52993),
            .I(N__52937));
    InMux I__12830 (
            .O(N__52992),
            .I(N__52937));
    InMux I__12829 (
            .O(N__52991),
            .I(N__52930));
    InMux I__12828 (
            .O(N__52990),
            .I(N__52927));
    InMux I__12827 (
            .O(N__52989),
            .I(N__52924));
    LocalMux I__12826 (
            .O(N__52986),
            .I(N__52917));
    Span4Mux_h I__12825 (
            .O(N__52983),
            .I(N__52917));
    LocalMux I__12824 (
            .O(N__52970),
            .I(N__52917));
    InMux I__12823 (
            .O(N__52967),
            .I(N__52912));
    LocalMux I__12822 (
            .O(N__52960),
            .I(N__52908));
    InMux I__12821 (
            .O(N__52959),
            .I(N__52903));
    InMux I__12820 (
            .O(N__52958),
            .I(N__52903));
    InMux I__12819 (
            .O(N__52955),
            .I(N__52900));
    InMux I__12818 (
            .O(N__52954),
            .I(N__52891));
    InMux I__12817 (
            .O(N__52953),
            .I(N__52891));
    InMux I__12816 (
            .O(N__52952),
            .I(N__52891));
    InMux I__12815 (
            .O(N__52951),
            .I(N__52891));
    LocalMux I__12814 (
            .O(N__52948),
            .I(N__52886));
    LocalMux I__12813 (
            .O(N__52945),
            .I(N__52886));
    LocalMux I__12812 (
            .O(N__52942),
            .I(N__52881));
    LocalMux I__12811 (
            .O(N__52937),
            .I(N__52881));
    InMux I__12810 (
            .O(N__52936),
            .I(N__52866));
    InMux I__12809 (
            .O(N__52935),
            .I(N__52866));
    InMux I__12808 (
            .O(N__52934),
            .I(N__52866));
    InMux I__12807 (
            .O(N__52933),
            .I(N__52866));
    LocalMux I__12806 (
            .O(N__52930),
            .I(N__52863));
    LocalMux I__12805 (
            .O(N__52927),
            .I(N__52858));
    LocalMux I__12804 (
            .O(N__52924),
            .I(N__52858));
    Span4Mux_v I__12803 (
            .O(N__52917),
            .I(N__52855));
    CascadeMux I__12802 (
            .O(N__52916),
            .I(N__52851));
    InMux I__12801 (
            .O(N__52915),
            .I(N__52841));
    LocalMux I__12800 (
            .O(N__52912),
            .I(N__52838));
    InMux I__12799 (
            .O(N__52911),
            .I(N__52835));
    Span4Mux_h I__12798 (
            .O(N__52908),
            .I(N__52832));
    LocalMux I__12797 (
            .O(N__52903),
            .I(N__52829));
    LocalMux I__12796 (
            .O(N__52900),
            .I(N__52820));
    LocalMux I__12795 (
            .O(N__52891),
            .I(N__52820));
    Span4Mux_h I__12794 (
            .O(N__52886),
            .I(N__52820));
    Span4Mux_h I__12793 (
            .O(N__52881),
            .I(N__52820));
    InMux I__12792 (
            .O(N__52880),
            .I(N__52806));
    InMux I__12791 (
            .O(N__52879),
            .I(N__52806));
    InMux I__12790 (
            .O(N__52878),
            .I(N__52806));
    InMux I__12789 (
            .O(N__52877),
            .I(N__52806));
    InMux I__12788 (
            .O(N__52876),
            .I(N__52806));
    InMux I__12787 (
            .O(N__52875),
            .I(N__52806));
    LocalMux I__12786 (
            .O(N__52866),
            .I(N__52801));
    Span4Mux_v I__12785 (
            .O(N__52863),
            .I(N__52801));
    Span4Mux_v I__12784 (
            .O(N__52858),
            .I(N__52796));
    Span4Mux_h I__12783 (
            .O(N__52855),
            .I(N__52796));
    InMux I__12782 (
            .O(N__52854),
            .I(N__52793));
    InMux I__12781 (
            .O(N__52851),
            .I(N__52788));
    InMux I__12780 (
            .O(N__52850),
            .I(N__52788));
    InMux I__12779 (
            .O(N__52849),
            .I(N__52779));
    InMux I__12778 (
            .O(N__52848),
            .I(N__52779));
    InMux I__12777 (
            .O(N__52847),
            .I(N__52779));
    InMux I__12776 (
            .O(N__52846),
            .I(N__52779));
    InMux I__12775 (
            .O(N__52845),
            .I(N__52774));
    InMux I__12774 (
            .O(N__52844),
            .I(N__52774));
    LocalMux I__12773 (
            .O(N__52841),
            .I(N__52769));
    Span4Mux_v I__12772 (
            .O(N__52838),
            .I(N__52769));
    LocalMux I__12771 (
            .O(N__52835),
            .I(N__52764));
    Span4Mux_v I__12770 (
            .O(N__52832),
            .I(N__52764));
    Span4Mux_h I__12769 (
            .O(N__52829),
            .I(N__52759));
    Span4Mux_v I__12768 (
            .O(N__52820),
            .I(N__52759));
    InMux I__12767 (
            .O(N__52819),
            .I(N__52743));
    LocalMux I__12766 (
            .O(N__52806),
            .I(N__52740));
    Span4Mux_v I__12765 (
            .O(N__52801),
            .I(N__52735));
    Span4Mux_h I__12764 (
            .O(N__52796),
            .I(N__52735));
    LocalMux I__12763 (
            .O(N__52793),
            .I(N__52722));
    LocalMux I__12762 (
            .O(N__52788),
            .I(N__52722));
    LocalMux I__12761 (
            .O(N__52779),
            .I(N__52722));
    LocalMux I__12760 (
            .O(N__52774),
            .I(N__52722));
    Span4Mux_h I__12759 (
            .O(N__52769),
            .I(N__52722));
    Span4Mux_v I__12758 (
            .O(N__52764),
            .I(N__52722));
    Span4Mux_v I__12757 (
            .O(N__52759),
            .I(N__52717));
    InMux I__12756 (
            .O(N__52758),
            .I(N__52710));
    InMux I__12755 (
            .O(N__52757),
            .I(N__52710));
    InMux I__12754 (
            .O(N__52756),
            .I(N__52710));
    InMux I__12753 (
            .O(N__52755),
            .I(N__52703));
    InMux I__12752 (
            .O(N__52754),
            .I(N__52696));
    InMux I__12751 (
            .O(N__52753),
            .I(N__52696));
    InMux I__12750 (
            .O(N__52752),
            .I(N__52696));
    InMux I__12749 (
            .O(N__52751),
            .I(N__52683));
    InMux I__12748 (
            .O(N__52750),
            .I(N__52683));
    InMux I__12747 (
            .O(N__52749),
            .I(N__52683));
    InMux I__12746 (
            .O(N__52748),
            .I(N__52683));
    InMux I__12745 (
            .O(N__52747),
            .I(N__52683));
    InMux I__12744 (
            .O(N__52746),
            .I(N__52683));
    LocalMux I__12743 (
            .O(N__52743),
            .I(N__52680));
    Span4Mux_v I__12742 (
            .O(N__52740),
            .I(N__52675));
    Span4Mux_h I__12741 (
            .O(N__52735),
            .I(N__52675));
    Span4Mux_h I__12740 (
            .O(N__52722),
            .I(N__52672));
    InMux I__12739 (
            .O(N__52721),
            .I(N__52667));
    InMux I__12738 (
            .O(N__52720),
            .I(N__52667));
    Span4Mux_h I__12737 (
            .O(N__52717),
            .I(N__52662));
    LocalMux I__12736 (
            .O(N__52710),
            .I(N__52662));
    InMux I__12735 (
            .O(N__52709),
            .I(N__52653));
    InMux I__12734 (
            .O(N__52708),
            .I(N__52653));
    InMux I__12733 (
            .O(N__52707),
            .I(N__52653));
    InMux I__12732 (
            .O(N__52706),
            .I(N__52653));
    LocalMux I__12731 (
            .O(N__52703),
            .I(adc_state_0_adj_1418));
    LocalMux I__12730 (
            .O(N__52696),
            .I(adc_state_0_adj_1418));
    LocalMux I__12729 (
            .O(N__52683),
            .I(adc_state_0_adj_1418));
    Odrv4 I__12728 (
            .O(N__52680),
            .I(adc_state_0_adj_1418));
    Odrv4 I__12727 (
            .O(N__52675),
            .I(adc_state_0_adj_1418));
    Odrv4 I__12726 (
            .O(N__52672),
            .I(adc_state_0_adj_1418));
    LocalMux I__12725 (
            .O(N__52667),
            .I(adc_state_0_adj_1418));
    Odrv4 I__12724 (
            .O(N__52662),
            .I(adc_state_0_adj_1418));
    LocalMux I__12723 (
            .O(N__52653),
            .I(adc_state_0_adj_1418));
    CascadeMux I__12722 (
            .O(N__52634),
            .I(N__52630));
    CascadeMux I__12721 (
            .O(N__52633),
            .I(N__52627));
    InMux I__12720 (
            .O(N__52630),
            .I(N__52623));
    InMux I__12719 (
            .O(N__52627),
            .I(N__52618));
    InMux I__12718 (
            .O(N__52626),
            .I(N__52618));
    LocalMux I__12717 (
            .O(N__52623),
            .I(cmd_rdadctmp_17_adj_1433));
    LocalMux I__12716 (
            .O(N__52618),
            .I(cmd_rdadctmp_17_adj_1433));
    InMux I__12715 (
            .O(N__52613),
            .I(N__52610));
    LocalMux I__12714 (
            .O(N__52610),
            .I(N__52606));
    InMux I__12713 (
            .O(N__52609),
            .I(N__52603));
    Span4Mux_h I__12712 (
            .O(N__52606),
            .I(N__52599));
    LocalMux I__12711 (
            .O(N__52603),
            .I(N__52596));
    InMux I__12710 (
            .O(N__52602),
            .I(N__52593));
    Span4Mux_v I__12709 (
            .O(N__52599),
            .I(N__52588));
    Span4Mux_h I__12708 (
            .O(N__52596),
            .I(N__52588));
    LocalMux I__12707 (
            .O(N__52593),
            .I(buf_adcdata_iac_9));
    Odrv4 I__12706 (
            .O(N__52588),
            .I(buf_adcdata_iac_9));
    InMux I__12705 (
            .O(N__52583),
            .I(N__52580));
    LocalMux I__12704 (
            .O(N__52580),
            .I(N__52577));
    Span4Mux_h I__12703 (
            .O(N__52577),
            .I(N__52574));
    Odrv4 I__12702 (
            .O(N__52574),
            .I(buf_data_iac_12));
    CascadeMux I__12701 (
            .O(N__52571),
            .I(N__52568));
    InMux I__12700 (
            .O(N__52568),
            .I(N__52565));
    LocalMux I__12699 (
            .O(N__52565),
            .I(N__52562));
    Span4Mux_h I__12698 (
            .O(N__52562),
            .I(N__52559));
    Span4Mux_h I__12697 (
            .O(N__52559),
            .I(N__52556));
    Odrv4 I__12696 (
            .O(N__52556),
            .I(n21230));
    InMux I__12695 (
            .O(N__52553),
            .I(N__52550));
    LocalMux I__12694 (
            .O(N__52550),
            .I(N__52547));
    Span4Mux_h I__12693 (
            .O(N__52547),
            .I(N__52544));
    Odrv4 I__12692 (
            .O(N__52544),
            .I(buf_data_iac_13));
    InMux I__12691 (
            .O(N__52541),
            .I(N__52538));
    LocalMux I__12690 (
            .O(N__52538),
            .I(N__52535));
    Span4Mux_v I__12689 (
            .O(N__52535),
            .I(N__52532));
    Span4Mux_h I__12688 (
            .O(N__52532),
            .I(N__52529));
    Odrv4 I__12687 (
            .O(N__52529),
            .I(n21297));
    SRMux I__12686 (
            .O(N__52526),
            .I(N__52523));
    LocalMux I__12685 (
            .O(N__52523),
            .I(N__52520));
    Span4Mux_h I__12684 (
            .O(N__52520),
            .I(N__52517));
    Span4Mux_v I__12683 (
            .O(N__52517),
            .I(N__52514));
    Odrv4 I__12682 (
            .O(N__52514),
            .I(\comm_spi.DOUT_7__N_747 ));
    CascadeMux I__12681 (
            .O(N__52511),
            .I(N__52508));
    InMux I__12680 (
            .O(N__52508),
            .I(N__52500));
    InMux I__12679 (
            .O(N__52507),
            .I(N__52500));
    CascadeMux I__12678 (
            .O(N__52506),
            .I(N__52497));
    InMux I__12677 (
            .O(N__52505),
            .I(N__52494));
    LocalMux I__12676 (
            .O(N__52500),
            .I(N__52490));
    InMux I__12675 (
            .O(N__52497),
            .I(N__52486));
    LocalMux I__12674 (
            .O(N__52494),
            .I(N__52483));
    InMux I__12673 (
            .O(N__52493),
            .I(N__52480));
    Span4Mux_v I__12672 (
            .O(N__52490),
            .I(N__52477));
    InMux I__12671 (
            .O(N__52489),
            .I(N__52474));
    LocalMux I__12670 (
            .O(N__52486),
            .I(N__52471));
    Span4Mux_v I__12669 (
            .O(N__52483),
            .I(N__52468));
    LocalMux I__12668 (
            .O(N__52480),
            .I(N__52465));
    Span4Mux_h I__12667 (
            .O(N__52477),
            .I(N__52460));
    LocalMux I__12666 (
            .O(N__52474),
            .I(N__52460));
    Span4Mux_v I__12665 (
            .O(N__52471),
            .I(N__52457));
    Sp12to4 I__12664 (
            .O(N__52468),
            .I(N__52454));
    Span4Mux_v I__12663 (
            .O(N__52465),
            .I(N__52451));
    Span4Mux_v I__12662 (
            .O(N__52460),
            .I(N__52448));
    Odrv4 I__12661 (
            .O(N__52457),
            .I(comm_buf_1_6));
    Odrv12 I__12660 (
            .O(N__52454),
            .I(comm_buf_1_6));
    Odrv4 I__12659 (
            .O(N__52451),
            .I(comm_buf_1_6));
    Odrv4 I__12658 (
            .O(N__52448),
            .I(comm_buf_1_6));
    InMux I__12657 (
            .O(N__52439),
            .I(N__52421));
    InMux I__12656 (
            .O(N__52438),
            .I(N__52421));
    InMux I__12655 (
            .O(N__52437),
            .I(N__52421));
    InMux I__12654 (
            .O(N__52436),
            .I(N__52421));
    InMux I__12653 (
            .O(N__52435),
            .I(N__52421));
    InMux I__12652 (
            .O(N__52434),
            .I(N__52417));
    InMux I__12651 (
            .O(N__52433),
            .I(N__52413));
    InMux I__12650 (
            .O(N__52432),
            .I(N__52403));
    LocalMux I__12649 (
            .O(N__52421),
            .I(N__52400));
    InMux I__12648 (
            .O(N__52420),
            .I(N__52397));
    LocalMux I__12647 (
            .O(N__52417),
            .I(N__52394));
    InMux I__12646 (
            .O(N__52416),
            .I(N__52384));
    LocalMux I__12645 (
            .O(N__52413),
            .I(N__52381));
    InMux I__12644 (
            .O(N__52412),
            .I(N__52371));
    InMux I__12643 (
            .O(N__52411),
            .I(N__52371));
    InMux I__12642 (
            .O(N__52410),
            .I(N__52361));
    InMux I__12641 (
            .O(N__52409),
            .I(N__52356));
    InMux I__12640 (
            .O(N__52408),
            .I(N__52356));
    InMux I__12639 (
            .O(N__52407),
            .I(N__52353));
    CascadeMux I__12638 (
            .O(N__52406),
            .I(N__52350));
    LocalMux I__12637 (
            .O(N__52403),
            .I(N__52345));
    Span4Mux_v I__12636 (
            .O(N__52400),
            .I(N__52342));
    LocalMux I__12635 (
            .O(N__52397),
            .I(N__52339));
    Span4Mux_h I__12634 (
            .O(N__52394),
            .I(N__52336));
    InMux I__12633 (
            .O(N__52393),
            .I(N__52327));
    InMux I__12632 (
            .O(N__52392),
            .I(N__52327));
    InMux I__12631 (
            .O(N__52391),
            .I(N__52327));
    InMux I__12630 (
            .O(N__52390),
            .I(N__52327));
    InMux I__12629 (
            .O(N__52389),
            .I(N__52319));
    InMux I__12628 (
            .O(N__52388),
            .I(N__52319));
    InMux I__12627 (
            .O(N__52387),
            .I(N__52319));
    LocalMux I__12626 (
            .O(N__52384),
            .I(N__52314));
    Span4Mux_h I__12625 (
            .O(N__52381),
            .I(N__52314));
    InMux I__12624 (
            .O(N__52380),
            .I(N__52307));
    InMux I__12623 (
            .O(N__52379),
            .I(N__52307));
    InMux I__12622 (
            .O(N__52378),
            .I(N__52307));
    InMux I__12621 (
            .O(N__52377),
            .I(N__52297));
    InMux I__12620 (
            .O(N__52376),
            .I(N__52297));
    LocalMux I__12619 (
            .O(N__52371),
            .I(N__52294));
    InMux I__12618 (
            .O(N__52370),
            .I(N__52289));
    InMux I__12617 (
            .O(N__52369),
            .I(N__52289));
    InMux I__12616 (
            .O(N__52368),
            .I(N__52286));
    InMux I__12615 (
            .O(N__52367),
            .I(N__52283));
    InMux I__12614 (
            .O(N__52366),
            .I(N__52280));
    InMux I__12613 (
            .O(N__52365),
            .I(N__52275));
    InMux I__12612 (
            .O(N__52364),
            .I(N__52275));
    LocalMux I__12611 (
            .O(N__52361),
            .I(N__52270));
    LocalMux I__12610 (
            .O(N__52356),
            .I(N__52270));
    LocalMux I__12609 (
            .O(N__52353),
            .I(N__52267));
    InMux I__12608 (
            .O(N__52350),
            .I(N__52260));
    InMux I__12607 (
            .O(N__52349),
            .I(N__52260));
    InMux I__12606 (
            .O(N__52348),
            .I(N__52260));
    Span4Mux_v I__12605 (
            .O(N__52345),
            .I(N__52254));
    Span4Mux_h I__12604 (
            .O(N__52342),
            .I(N__52254));
    Span4Mux_h I__12603 (
            .O(N__52339),
            .I(N__52247));
    Span4Mux_v I__12602 (
            .O(N__52336),
            .I(N__52247));
    LocalMux I__12601 (
            .O(N__52327),
            .I(N__52247));
    InMux I__12600 (
            .O(N__52326),
            .I(N__52244));
    LocalMux I__12599 (
            .O(N__52319),
            .I(N__52237));
    Sp12to4 I__12598 (
            .O(N__52314),
            .I(N__52237));
    LocalMux I__12597 (
            .O(N__52307),
            .I(N__52237));
    InMux I__12596 (
            .O(N__52306),
            .I(N__52232));
    InMux I__12595 (
            .O(N__52305),
            .I(N__52232));
    InMux I__12594 (
            .O(N__52304),
            .I(N__52225));
    InMux I__12593 (
            .O(N__52303),
            .I(N__52225));
    InMux I__12592 (
            .O(N__52302),
            .I(N__52225));
    LocalMux I__12591 (
            .O(N__52297),
            .I(N__52216));
    Span4Mux_v I__12590 (
            .O(N__52294),
            .I(N__52216));
    LocalMux I__12589 (
            .O(N__52289),
            .I(N__52216));
    LocalMux I__12588 (
            .O(N__52286),
            .I(N__52216));
    LocalMux I__12587 (
            .O(N__52283),
            .I(N__52203));
    LocalMux I__12586 (
            .O(N__52280),
            .I(N__52203));
    LocalMux I__12585 (
            .O(N__52275),
            .I(N__52203));
    Sp12to4 I__12584 (
            .O(N__52270),
            .I(N__52203));
    Span12Mux_h I__12583 (
            .O(N__52267),
            .I(N__52203));
    LocalMux I__12582 (
            .O(N__52260),
            .I(N__52203));
    InMux I__12581 (
            .O(N__52259),
            .I(N__52200));
    Span4Mux_h I__12580 (
            .O(N__52254),
            .I(N__52195));
    Span4Mux_v I__12579 (
            .O(N__52247),
            .I(N__52195));
    LocalMux I__12578 (
            .O(N__52244),
            .I(N__52190));
    Span12Mux_v I__12577 (
            .O(N__52237),
            .I(N__52190));
    LocalMux I__12576 (
            .O(N__52232),
            .I(comm_state_2));
    LocalMux I__12575 (
            .O(N__52225),
            .I(comm_state_2));
    Odrv4 I__12574 (
            .O(N__52216),
            .I(comm_state_2));
    Odrv12 I__12573 (
            .O(N__52203),
            .I(comm_state_2));
    LocalMux I__12572 (
            .O(N__52200),
            .I(comm_state_2));
    Odrv4 I__12571 (
            .O(N__52195),
            .I(comm_state_2));
    Odrv12 I__12570 (
            .O(N__52190),
            .I(comm_state_2));
    InMux I__12569 (
            .O(N__52175),
            .I(N__52171));
    InMux I__12568 (
            .O(N__52174),
            .I(N__52168));
    LocalMux I__12567 (
            .O(N__52171),
            .I(N__52165));
    LocalMux I__12566 (
            .O(N__52168),
            .I(N__52160));
    Span4Mux_h I__12565 (
            .O(N__52165),
            .I(N__52160));
    Odrv4 I__12564 (
            .O(N__52160),
            .I(n14_adj_1547));
    CascadeMux I__12563 (
            .O(N__52157),
            .I(N__52154));
    InMux I__12562 (
            .O(N__52154),
            .I(N__52150));
    InMux I__12561 (
            .O(N__52153),
            .I(N__52147));
    LocalMux I__12560 (
            .O(N__52150),
            .I(N__52144));
    LocalMux I__12559 (
            .O(N__52147),
            .I(N__52140));
    Span4Mux_v I__12558 (
            .O(N__52144),
            .I(N__52137));
    InMux I__12557 (
            .O(N__52143),
            .I(N__52134));
    Span12Mux_s10_h I__12556 (
            .O(N__52140),
            .I(N__52131));
    Span4Mux_h I__12555 (
            .O(N__52137),
            .I(N__52128));
    LocalMux I__12554 (
            .O(N__52134),
            .I(buf_adcdata_iac_8));
    Odrv12 I__12553 (
            .O(N__52131),
            .I(buf_adcdata_iac_8));
    Odrv4 I__12552 (
            .O(N__52128),
            .I(buf_adcdata_iac_8));
    CascadeMux I__12551 (
            .O(N__52121),
            .I(N__52117));
    CascadeMux I__12550 (
            .O(N__52120),
            .I(N__52114));
    InMux I__12549 (
            .O(N__52117),
            .I(N__52109));
    InMux I__12548 (
            .O(N__52114),
            .I(N__52109));
    LocalMux I__12547 (
            .O(N__52109),
            .I(N__52106));
    Span12Mux_v I__12546 (
            .O(N__52106),
            .I(N__52102));
    InMux I__12545 (
            .O(N__52105),
            .I(N__52099));
    Odrv12 I__12544 (
            .O(N__52102),
            .I(cmd_rdadctmp_16_adj_1434));
    LocalMux I__12543 (
            .O(N__52099),
            .I(cmd_rdadctmp_16_adj_1434));
    InMux I__12542 (
            .O(N__52094),
            .I(N__52091));
    LocalMux I__12541 (
            .O(N__52091),
            .I(N__52082));
    InMux I__12540 (
            .O(N__52090),
            .I(N__52079));
    InMux I__12539 (
            .O(N__52089),
            .I(N__52068));
    InMux I__12538 (
            .O(N__52088),
            .I(N__52065));
    InMux I__12537 (
            .O(N__52087),
            .I(N__52058));
    InMux I__12536 (
            .O(N__52086),
            .I(N__52058));
    InMux I__12535 (
            .O(N__52085),
            .I(N__52058));
    Span4Mux_h I__12534 (
            .O(N__52082),
            .I(N__52053));
    LocalMux I__12533 (
            .O(N__52079),
            .I(N__52053));
    InMux I__12532 (
            .O(N__52078),
            .I(N__52048));
    InMux I__12531 (
            .O(N__52077),
            .I(N__52048));
    InMux I__12530 (
            .O(N__52076),
            .I(N__52043));
    InMux I__12529 (
            .O(N__52075),
            .I(N__52040));
    InMux I__12528 (
            .O(N__52074),
            .I(N__52031));
    InMux I__12527 (
            .O(N__52073),
            .I(N__52031));
    InMux I__12526 (
            .O(N__52072),
            .I(N__52031));
    InMux I__12525 (
            .O(N__52071),
            .I(N__52031));
    LocalMux I__12524 (
            .O(N__52068),
            .I(N__52028));
    LocalMux I__12523 (
            .O(N__52065),
            .I(N__52023));
    LocalMux I__12522 (
            .O(N__52058),
            .I(N__52023));
    Span4Mux_v I__12521 (
            .O(N__52053),
            .I(N__52020));
    LocalMux I__12520 (
            .O(N__52048),
            .I(N__52017));
    InMux I__12519 (
            .O(N__52047),
            .I(N__52009));
    InMux I__12518 (
            .O(N__52046),
            .I(N__52009));
    LocalMux I__12517 (
            .O(N__52043),
            .I(N__52006));
    LocalMux I__12516 (
            .O(N__52040),
            .I(N__51999));
    LocalMux I__12515 (
            .O(N__52031),
            .I(N__51994));
    Sp12to4 I__12514 (
            .O(N__52028),
            .I(N__51994));
    Span4Mux_v I__12513 (
            .O(N__52023),
            .I(N__51991));
    Span4Mux_h I__12512 (
            .O(N__52020),
            .I(N__51988));
    Span4Mux_v I__12511 (
            .O(N__52017),
            .I(N__51985));
    InMux I__12510 (
            .O(N__52016),
            .I(N__51974));
    InMux I__12509 (
            .O(N__52015),
            .I(N__51969));
    InMux I__12508 (
            .O(N__52014),
            .I(N__51969));
    LocalMux I__12507 (
            .O(N__52009),
            .I(N__51964));
    Span4Mux_h I__12506 (
            .O(N__52006),
            .I(N__51964));
    InMux I__12505 (
            .O(N__52005),
            .I(N__51959));
    InMux I__12504 (
            .O(N__52004),
            .I(N__51959));
    InMux I__12503 (
            .O(N__52003),
            .I(N__51954));
    InMux I__12502 (
            .O(N__52002),
            .I(N__51954));
    Sp12to4 I__12501 (
            .O(N__51999),
            .I(N__51947));
    Span12Mux_v I__12500 (
            .O(N__51994),
            .I(N__51947));
    Sp12to4 I__12499 (
            .O(N__51991),
            .I(N__51947));
    Sp12to4 I__12498 (
            .O(N__51988),
            .I(N__51942));
    Sp12to4 I__12497 (
            .O(N__51985),
            .I(N__51942));
    InMux I__12496 (
            .O(N__51984),
            .I(N__51937));
    InMux I__12495 (
            .O(N__51983),
            .I(N__51937));
    InMux I__12494 (
            .O(N__51982),
            .I(N__51932));
    InMux I__12493 (
            .O(N__51981),
            .I(N__51932));
    InMux I__12492 (
            .O(N__51980),
            .I(N__51923));
    InMux I__12491 (
            .O(N__51979),
            .I(N__51923));
    InMux I__12490 (
            .O(N__51978),
            .I(N__51923));
    InMux I__12489 (
            .O(N__51977),
            .I(N__51923));
    LocalMux I__12488 (
            .O(N__51974),
            .I(N__51920));
    LocalMux I__12487 (
            .O(N__51969),
            .I(N__51915));
    Span4Mux_h I__12486 (
            .O(N__51964),
            .I(N__51915));
    LocalMux I__12485 (
            .O(N__51959),
            .I(N__51908));
    LocalMux I__12484 (
            .O(N__51954),
            .I(N__51908));
    Span12Mux_h I__12483 (
            .O(N__51947),
            .I(N__51908));
    Span12Mux_h I__12482 (
            .O(N__51942),
            .I(N__51905));
    LocalMux I__12481 (
            .O(N__51937),
            .I(n12663));
    LocalMux I__12480 (
            .O(N__51932),
            .I(n12663));
    LocalMux I__12479 (
            .O(N__51923),
            .I(n12663));
    Odrv4 I__12478 (
            .O(N__51920),
            .I(n12663));
    Odrv4 I__12477 (
            .O(N__51915),
            .I(n12663));
    Odrv12 I__12476 (
            .O(N__51908),
            .I(n12663));
    Odrv12 I__12475 (
            .O(N__51905),
            .I(n12663));
    CascadeMux I__12474 (
            .O(N__51890),
            .I(N__51886));
    InMux I__12473 (
            .O(N__51889),
            .I(N__51878));
    InMux I__12472 (
            .O(N__51886),
            .I(N__51878));
    InMux I__12471 (
            .O(N__51885),
            .I(N__51878));
    LocalMux I__12470 (
            .O(N__51878),
            .I(cmd_rdadctmp_18_adj_1432));
    InMux I__12469 (
            .O(N__51875),
            .I(N__51870));
    CascadeMux I__12468 (
            .O(N__51874),
            .I(N__51867));
    CascadeMux I__12467 (
            .O(N__51873),
            .I(N__51864));
    LocalMux I__12466 (
            .O(N__51870),
            .I(N__51861));
    InMux I__12465 (
            .O(N__51867),
            .I(N__51858));
    InMux I__12464 (
            .O(N__51864),
            .I(N__51855));
    Span12Mux_v I__12463 (
            .O(N__51861),
            .I(N__51852));
    LocalMux I__12462 (
            .O(N__51858),
            .I(buf_adcdata_iac_10));
    LocalMux I__12461 (
            .O(N__51855),
            .I(buf_adcdata_iac_10));
    Odrv12 I__12460 (
            .O(N__51852),
            .I(buf_adcdata_iac_10));
    CascadeMux I__12459 (
            .O(N__51845),
            .I(N__51835));
    CascadeMux I__12458 (
            .O(N__51844),
            .I(N__51832));
    CascadeMux I__12457 (
            .O(N__51843),
            .I(N__51829));
    InMux I__12456 (
            .O(N__51842),
            .I(N__51820));
    InMux I__12455 (
            .O(N__51841),
            .I(N__51820));
    InMux I__12454 (
            .O(N__51840),
            .I(N__51817));
    InMux I__12453 (
            .O(N__51839),
            .I(N__51814));
    CascadeMux I__12452 (
            .O(N__51838),
            .I(N__51811));
    InMux I__12451 (
            .O(N__51835),
            .I(N__51804));
    InMux I__12450 (
            .O(N__51832),
            .I(N__51804));
    InMux I__12449 (
            .O(N__51829),
            .I(N__51804));
    InMux I__12448 (
            .O(N__51828),
            .I(N__51801));
    InMux I__12447 (
            .O(N__51827),
            .I(N__51794));
    InMux I__12446 (
            .O(N__51826),
            .I(N__51794));
    InMux I__12445 (
            .O(N__51825),
            .I(N__51794));
    LocalMux I__12444 (
            .O(N__51820),
            .I(N__51789));
    LocalMux I__12443 (
            .O(N__51817),
            .I(N__51789));
    LocalMux I__12442 (
            .O(N__51814),
            .I(N__51786));
    InMux I__12441 (
            .O(N__51811),
            .I(N__51783));
    LocalMux I__12440 (
            .O(N__51804),
            .I(N__51777));
    LocalMux I__12439 (
            .O(N__51801),
            .I(N__51777));
    LocalMux I__12438 (
            .O(N__51794),
            .I(N__51774));
    Span4Mux_v I__12437 (
            .O(N__51789),
            .I(N__51767));
    Span4Mux_h I__12436 (
            .O(N__51786),
            .I(N__51767));
    LocalMux I__12435 (
            .O(N__51783),
            .I(N__51767));
    CascadeMux I__12434 (
            .O(N__51782),
            .I(N__51763));
    Span4Mux_v I__12433 (
            .O(N__51777),
            .I(N__51759));
    Span4Mux_v I__12432 (
            .O(N__51774),
            .I(N__51756));
    Span4Mux_v I__12431 (
            .O(N__51767),
            .I(N__51753));
    InMux I__12430 (
            .O(N__51766),
            .I(N__51748));
    InMux I__12429 (
            .O(N__51763),
            .I(N__51748));
    CascadeMux I__12428 (
            .O(N__51762),
            .I(N__51742));
    Sp12to4 I__12427 (
            .O(N__51759),
            .I(N__51738));
    Sp12to4 I__12426 (
            .O(N__51756),
            .I(N__51735));
    Span4Mux_h I__12425 (
            .O(N__51753),
            .I(N__51732));
    LocalMux I__12424 (
            .O(N__51748),
            .I(N__51729));
    InMux I__12423 (
            .O(N__51747),
            .I(N__51724));
    InMux I__12422 (
            .O(N__51746),
            .I(N__51724));
    InMux I__12421 (
            .O(N__51745),
            .I(N__51717));
    InMux I__12420 (
            .O(N__51742),
            .I(N__51717));
    InMux I__12419 (
            .O(N__51741),
            .I(N__51717));
    Span12Mux_h I__12418 (
            .O(N__51738),
            .I(N__51714));
    Span12Mux_s10_h I__12417 (
            .O(N__51735),
            .I(N__51703));
    Sp12to4 I__12416 (
            .O(N__51732),
            .I(N__51703));
    Sp12to4 I__12415 (
            .O(N__51729),
            .I(N__51703));
    LocalMux I__12414 (
            .O(N__51724),
            .I(N__51703));
    LocalMux I__12413 (
            .O(N__51717),
            .I(N__51703));
    Span12Mux_v I__12412 (
            .O(N__51714),
            .I(N__51700));
    Span12Mux_v I__12411 (
            .O(N__51703),
            .I(N__51697));
    Odrv12 I__12410 (
            .O(N__51700),
            .I(ICE_SPI_CE0));
    Odrv12 I__12409 (
            .O(N__51697),
            .I(ICE_SPI_CE0));
    InMux I__12408 (
            .O(N__51692),
            .I(N__51683));
    InMux I__12407 (
            .O(N__51691),
            .I(N__51683));
    InMux I__12406 (
            .O(N__51690),
            .I(N__51680));
    InMux I__12405 (
            .O(N__51689),
            .I(N__51677));
    InMux I__12404 (
            .O(N__51688),
            .I(N__51674));
    LocalMux I__12403 (
            .O(N__51683),
            .I(N__51666));
    LocalMux I__12402 (
            .O(N__51680),
            .I(N__51663));
    LocalMux I__12401 (
            .O(N__51677),
            .I(N__51658));
    LocalMux I__12400 (
            .O(N__51674),
            .I(N__51658));
    InMux I__12399 (
            .O(N__51673),
            .I(N__51653));
    InMux I__12398 (
            .O(N__51672),
            .I(N__51653));
    InMux I__12397 (
            .O(N__51671),
            .I(N__51648));
    InMux I__12396 (
            .O(N__51670),
            .I(N__51648));
    CascadeMux I__12395 (
            .O(N__51669),
            .I(N__51643));
    Span4Mux_h I__12394 (
            .O(N__51666),
            .I(N__51639));
    Span4Mux_v I__12393 (
            .O(N__51663),
            .I(N__51632));
    Span4Mux_v I__12392 (
            .O(N__51658),
            .I(N__51632));
    LocalMux I__12391 (
            .O(N__51653),
            .I(N__51632));
    LocalMux I__12390 (
            .O(N__51648),
            .I(N__51629));
    InMux I__12389 (
            .O(N__51647),
            .I(N__51620));
    InMux I__12388 (
            .O(N__51646),
            .I(N__51620));
    InMux I__12387 (
            .O(N__51643),
            .I(N__51620));
    InMux I__12386 (
            .O(N__51642),
            .I(N__51620));
    Odrv4 I__12385 (
            .O(N__51639),
            .I(comm_data_vld));
    Odrv4 I__12384 (
            .O(N__51632),
            .I(comm_data_vld));
    Odrv4 I__12383 (
            .O(N__51629),
            .I(comm_data_vld));
    LocalMux I__12382 (
            .O(N__51620),
            .I(comm_data_vld));
    InMux I__12381 (
            .O(N__51611),
            .I(N__51608));
    LocalMux I__12380 (
            .O(N__51608),
            .I(n21129));
    CascadeMux I__12379 (
            .O(N__51605),
            .I(N__51602));
    InMux I__12378 (
            .O(N__51602),
            .I(N__51599));
    LocalMux I__12377 (
            .O(N__51599),
            .I(N__51596));
    Odrv4 I__12376 (
            .O(N__51596),
            .I(n20740));
    CascadeMux I__12375 (
            .O(N__51593),
            .I(n11363_cascade_));
    CascadeMux I__12374 (
            .O(N__51590),
            .I(N__51586));
    InMux I__12373 (
            .O(N__51589),
            .I(N__51581));
    InMux I__12372 (
            .O(N__51586),
            .I(N__51574));
    InMux I__12371 (
            .O(N__51585),
            .I(N__51574));
    InMux I__12370 (
            .O(N__51584),
            .I(N__51574));
    LocalMux I__12369 (
            .O(N__51581),
            .I(N__51570));
    LocalMux I__12368 (
            .O(N__51574),
            .I(N__51565));
    CascadeMux I__12367 (
            .O(N__51573),
            .I(N__51562));
    Span4Mux_v I__12366 (
            .O(N__51570),
            .I(N__51559));
    CascadeMux I__12365 (
            .O(N__51569),
            .I(N__51556));
    InMux I__12364 (
            .O(N__51568),
            .I(N__51553));
    Span4Mux_h I__12363 (
            .O(N__51565),
            .I(N__51546));
    InMux I__12362 (
            .O(N__51562),
            .I(N__51543));
    Span4Mux_v I__12361 (
            .O(N__51559),
            .I(N__51539));
    InMux I__12360 (
            .O(N__51556),
            .I(N__51536));
    LocalMux I__12359 (
            .O(N__51553),
            .I(N__51533));
    InMux I__12358 (
            .O(N__51552),
            .I(N__51530));
    InMux I__12357 (
            .O(N__51551),
            .I(N__51527));
    InMux I__12356 (
            .O(N__51550),
            .I(N__51522));
    InMux I__12355 (
            .O(N__51549),
            .I(N__51522));
    Span4Mux_h I__12354 (
            .O(N__51546),
            .I(N__51519));
    LocalMux I__12353 (
            .O(N__51543),
            .I(N__51516));
    InMux I__12352 (
            .O(N__51542),
            .I(N__51513));
    Sp12to4 I__12351 (
            .O(N__51539),
            .I(N__51508));
    LocalMux I__12350 (
            .O(N__51536),
            .I(N__51508));
    Span4Mux_h I__12349 (
            .O(N__51533),
            .I(N__51505));
    LocalMux I__12348 (
            .O(N__51530),
            .I(N__51498));
    LocalMux I__12347 (
            .O(N__51527),
            .I(N__51498));
    LocalMux I__12346 (
            .O(N__51522),
            .I(N__51498));
    Span4Mux_v I__12345 (
            .O(N__51519),
            .I(N__51493));
    Span4Mux_h I__12344 (
            .O(N__51516),
            .I(N__51493));
    LocalMux I__12343 (
            .O(N__51513),
            .I(n12242));
    Odrv12 I__12342 (
            .O(N__51508),
            .I(n12242));
    Odrv4 I__12341 (
            .O(N__51505),
            .I(n12242));
    Odrv4 I__12340 (
            .O(N__51498),
            .I(n12242));
    Odrv4 I__12339 (
            .O(N__51493),
            .I(n12242));
    InMux I__12338 (
            .O(N__51482),
            .I(N__51478));
    CascadeMux I__12337 (
            .O(N__51481),
            .I(N__51473));
    LocalMux I__12336 (
            .O(N__51478),
            .I(N__51470));
    InMux I__12335 (
            .O(N__51477),
            .I(N__51465));
    InMux I__12334 (
            .O(N__51476),
            .I(N__51465));
    InMux I__12333 (
            .O(N__51473),
            .I(N__51462));
    Odrv4 I__12332 (
            .O(N__51470),
            .I(n12235));
    LocalMux I__12331 (
            .O(N__51465),
            .I(n12235));
    LocalMux I__12330 (
            .O(N__51462),
            .I(n12235));
    InMux I__12329 (
            .O(N__51455),
            .I(N__51452));
    LocalMux I__12328 (
            .O(N__51452),
            .I(N__51449));
    Span4Mux_h I__12327 (
            .O(N__51449),
            .I(N__51446));
    Odrv4 I__12326 (
            .O(N__51446),
            .I(n11869));
    CEMux I__12325 (
            .O(N__51443),
            .I(N__51439));
    InMux I__12324 (
            .O(N__51442),
            .I(N__51436));
    LocalMux I__12323 (
            .O(N__51439),
            .I(N__51432));
    LocalMux I__12322 (
            .O(N__51436),
            .I(N__51429));
    InMux I__12321 (
            .O(N__51435),
            .I(N__51426));
    Span4Mux_h I__12320 (
            .O(N__51432),
            .I(N__51423));
    Span4Mux_h I__12319 (
            .O(N__51429),
            .I(N__51418));
    LocalMux I__12318 (
            .O(N__51426),
            .I(N__51418));
    Span4Mux_v I__12317 (
            .O(N__51423),
            .I(N__51415));
    Span4Mux_v I__12316 (
            .O(N__51418),
            .I(N__51412));
    Odrv4 I__12315 (
            .O(N__51415),
            .I(n11876));
    Odrv4 I__12314 (
            .O(N__51412),
            .I(n11876));
    CascadeMux I__12313 (
            .O(N__51407),
            .I(N__51402));
    InMux I__12312 (
            .O(N__51406),
            .I(N__51399));
    InMux I__12311 (
            .O(N__51405),
            .I(N__51395));
    InMux I__12310 (
            .O(N__51402),
            .I(N__51390));
    LocalMux I__12309 (
            .O(N__51399),
            .I(N__51387));
    CascadeMux I__12308 (
            .O(N__51398),
            .I(N__51384));
    LocalMux I__12307 (
            .O(N__51395),
            .I(N__51380));
    InMux I__12306 (
            .O(N__51394),
            .I(N__51377));
    InMux I__12305 (
            .O(N__51393),
            .I(N__51374));
    LocalMux I__12304 (
            .O(N__51390),
            .I(N__51371));
    Span4Mux_v I__12303 (
            .O(N__51387),
            .I(N__51368));
    InMux I__12302 (
            .O(N__51384),
            .I(N__51365));
    InMux I__12301 (
            .O(N__51383),
            .I(N__51362));
    Span4Mux_v I__12300 (
            .O(N__51380),
            .I(N__51359));
    LocalMux I__12299 (
            .O(N__51377),
            .I(N__51356));
    LocalMux I__12298 (
            .O(N__51374),
            .I(N__51353));
    Span4Mux_v I__12297 (
            .O(N__51371),
            .I(N__51350));
    Span4Mux_h I__12296 (
            .O(N__51368),
            .I(N__51343));
    LocalMux I__12295 (
            .O(N__51365),
            .I(N__51343));
    LocalMux I__12294 (
            .O(N__51362),
            .I(N__51343));
    Span4Mux_h I__12293 (
            .O(N__51359),
            .I(N__51335));
    Span4Mux_v I__12292 (
            .O(N__51356),
            .I(N__51335));
    Span4Mux_h I__12291 (
            .O(N__51353),
            .I(N__51335));
    Span4Mux_v I__12290 (
            .O(N__51350),
            .I(N__51330));
    Span4Mux_v I__12289 (
            .O(N__51343),
            .I(N__51330));
    InMux I__12288 (
            .O(N__51342),
            .I(N__51327));
    Odrv4 I__12287 (
            .O(N__51335),
            .I(comm_rx_buf_7));
    Odrv4 I__12286 (
            .O(N__51330),
            .I(comm_rx_buf_7));
    LocalMux I__12285 (
            .O(N__51327),
            .I(comm_rx_buf_7));
    InMux I__12284 (
            .O(N__51320),
            .I(N__51314));
    InMux I__12283 (
            .O(N__51319),
            .I(N__51314));
    LocalMux I__12282 (
            .O(N__51314),
            .I(N__51308));
    InMux I__12281 (
            .O(N__51313),
            .I(N__51303));
    InMux I__12280 (
            .O(N__51312),
            .I(N__51303));
    InMux I__12279 (
            .O(N__51311),
            .I(N__51300));
    Span4Mux_h I__12278 (
            .O(N__51308),
            .I(N__51293));
    LocalMux I__12277 (
            .O(N__51303),
            .I(N__51293));
    LocalMux I__12276 (
            .O(N__51300),
            .I(N__51290));
    InMux I__12275 (
            .O(N__51299),
            .I(N__51285));
    InMux I__12274 (
            .O(N__51298),
            .I(N__51285));
    Span4Mux_h I__12273 (
            .O(N__51293),
            .I(N__51281));
    Span4Mux_v I__12272 (
            .O(N__51290),
            .I(N__51276));
    LocalMux I__12271 (
            .O(N__51285),
            .I(N__51276));
    InMux I__12270 (
            .O(N__51284),
            .I(N__51273));
    Odrv4 I__12269 (
            .O(N__51281),
            .I(n12244));
    Odrv4 I__12268 (
            .O(N__51276),
            .I(n12244));
    LocalMux I__12267 (
            .O(N__51273),
            .I(n12244));
    InMux I__12266 (
            .O(N__51266),
            .I(N__51262));
    InMux I__12265 (
            .O(N__51265),
            .I(N__51259));
    LocalMux I__12264 (
            .O(N__51262),
            .I(comm_buf_6_7));
    LocalMux I__12263 (
            .O(N__51259),
            .I(comm_buf_6_7));
    InMux I__12262 (
            .O(N__51254),
            .I(N__51251));
    LocalMux I__12261 (
            .O(N__51251),
            .I(N__51248));
    Span4Mux_v I__12260 (
            .O(N__51248),
            .I(N__51245));
    Span4Mux_v I__12259 (
            .O(N__51245),
            .I(N__51242));
    Sp12to4 I__12258 (
            .O(N__51242),
            .I(N__51239));
    Span12Mux_h I__12257 (
            .O(N__51239),
            .I(N__51236));
    Odrv12 I__12256 (
            .O(N__51236),
            .I(THERMOSTAT));
    InMux I__12255 (
            .O(N__51233),
            .I(N__51230));
    LocalMux I__12254 (
            .O(N__51230),
            .I(N__51227));
    Odrv4 I__12253 (
            .O(N__51227),
            .I(buf_control_7));
    CEMux I__12252 (
            .O(N__51224),
            .I(N__51221));
    LocalMux I__12251 (
            .O(N__51221),
            .I(N__51218));
    Span4Mux_v I__12250 (
            .O(N__51218),
            .I(N__51215));
    Odrv4 I__12249 (
            .O(N__51215),
            .I(n11935));
    SRMux I__12248 (
            .O(N__51212),
            .I(N__51209));
    LocalMux I__12247 (
            .O(N__51209),
            .I(N__51205));
    SRMux I__12246 (
            .O(N__51208),
            .I(N__51202));
    Span4Mux_v I__12245 (
            .O(N__51205),
            .I(N__51197));
    LocalMux I__12244 (
            .O(N__51202),
            .I(N__51197));
    Span4Mux_h I__12243 (
            .O(N__51197),
            .I(N__51194));
    Span4Mux_h I__12242 (
            .O(N__51194),
            .I(N__51191));
    Odrv4 I__12241 (
            .O(N__51191),
            .I(n19904));
    CascadeMux I__12240 (
            .O(N__51188),
            .I(N__51184));
    CascadeMux I__12239 (
            .O(N__51187),
            .I(N__51178));
    InMux I__12238 (
            .O(N__51184),
            .I(N__51175));
    InMux I__12237 (
            .O(N__51183),
            .I(N__51172));
    InMux I__12236 (
            .O(N__51182),
            .I(N__51169));
    InMux I__12235 (
            .O(N__51181),
            .I(N__51165));
    InMux I__12234 (
            .O(N__51178),
            .I(N__51162));
    LocalMux I__12233 (
            .O(N__51175),
            .I(N__51157));
    LocalMux I__12232 (
            .O(N__51172),
            .I(N__51157));
    LocalMux I__12231 (
            .O(N__51169),
            .I(N__51154));
    InMux I__12230 (
            .O(N__51168),
            .I(N__51151));
    LocalMux I__12229 (
            .O(N__51165),
            .I(N__51148));
    LocalMux I__12228 (
            .O(N__51162),
            .I(N__51145));
    Span4Mux_v I__12227 (
            .O(N__51157),
            .I(N__51142));
    Span4Mux_v I__12226 (
            .O(N__51154),
            .I(N__51139));
    LocalMux I__12225 (
            .O(N__51151),
            .I(N__51136));
    Span4Mux_v I__12224 (
            .O(N__51148),
            .I(N__51133));
    Span4Mux_v I__12223 (
            .O(N__51145),
            .I(N__51124));
    Span4Mux_h I__12222 (
            .O(N__51142),
            .I(N__51124));
    Span4Mux_v I__12221 (
            .O(N__51139),
            .I(N__51124));
    Span4Mux_v I__12220 (
            .O(N__51136),
            .I(N__51124));
    Odrv4 I__12219 (
            .O(N__51133),
            .I(comm_buf_1_4));
    Odrv4 I__12218 (
            .O(N__51124),
            .I(comm_buf_1_4));
    InMux I__12217 (
            .O(N__51119),
            .I(N__51115));
    InMux I__12216 (
            .O(N__51118),
            .I(N__51112));
    LocalMux I__12215 (
            .O(N__51115),
            .I(N__51109));
    LocalMux I__12214 (
            .O(N__51112),
            .I(N__51106));
    Span4Mux_h I__12213 (
            .O(N__51109),
            .I(N__51103));
    Span4Mux_h I__12212 (
            .O(N__51106),
            .I(N__51100));
    Odrv4 I__12211 (
            .O(N__51103),
            .I(n14_adj_1548));
    Odrv4 I__12210 (
            .O(N__51100),
            .I(n14_adj_1548));
    InMux I__12209 (
            .O(N__51095),
            .I(N__51091));
    CascadeMux I__12208 (
            .O(N__51094),
            .I(N__51088));
    LocalMux I__12207 (
            .O(N__51091),
            .I(N__51085));
    InMux I__12206 (
            .O(N__51088),
            .I(N__51082));
    Span4Mux_v I__12205 (
            .O(N__51085),
            .I(N__51077));
    LocalMux I__12204 (
            .O(N__51082),
            .I(N__51077));
    Span4Mux_h I__12203 (
            .O(N__51077),
            .I(N__51073));
    CascadeMux I__12202 (
            .O(N__51076),
            .I(N__51070));
    Span4Mux_h I__12201 (
            .O(N__51073),
            .I(N__51067));
    InMux I__12200 (
            .O(N__51070),
            .I(N__51064));
    Odrv4 I__12199 (
            .O(N__51067),
            .I(cmd_rdadctmp_20_adj_1430));
    LocalMux I__12198 (
            .O(N__51064),
            .I(cmd_rdadctmp_20_adj_1430));
    CascadeMux I__12197 (
            .O(N__51059),
            .I(N__51056));
    InMux I__12196 (
            .O(N__51056),
            .I(N__51051));
    InMux I__12195 (
            .O(N__51055),
            .I(N__51048));
    InMux I__12194 (
            .O(N__51054),
            .I(N__51044));
    LocalMux I__12193 (
            .O(N__51051),
            .I(N__51039));
    LocalMux I__12192 (
            .O(N__51048),
            .I(N__51036));
    CascadeMux I__12191 (
            .O(N__51047),
            .I(N__51033));
    LocalMux I__12190 (
            .O(N__51044),
            .I(N__51029));
    InMux I__12189 (
            .O(N__51043),
            .I(N__51026));
    InMux I__12188 (
            .O(N__51042),
            .I(N__51023));
    Span4Mux_v I__12187 (
            .O(N__51039),
            .I(N__51018));
    Span4Mux_v I__12186 (
            .O(N__51036),
            .I(N__51018));
    InMux I__12185 (
            .O(N__51033),
            .I(N__51015));
    InMux I__12184 (
            .O(N__51032),
            .I(N__51012));
    Span4Mux_v I__12183 (
            .O(N__51029),
            .I(N__51009));
    LocalMux I__12182 (
            .O(N__51026),
            .I(N__51006));
    LocalMux I__12181 (
            .O(N__51023),
            .I(N__51003));
    Span4Mux_h I__12180 (
            .O(N__51018),
            .I(N__50996));
    LocalMux I__12179 (
            .O(N__51015),
            .I(N__50996));
    LocalMux I__12178 (
            .O(N__51012),
            .I(N__50996));
    Span4Mux_v I__12177 (
            .O(N__51009),
            .I(N__50989));
    Span4Mux_h I__12176 (
            .O(N__51006),
            .I(N__50989));
    Span4Mux_v I__12175 (
            .O(N__51003),
            .I(N__50984));
    Span4Mux_v I__12174 (
            .O(N__50996),
            .I(N__50984));
    InMux I__12173 (
            .O(N__50995),
            .I(N__50981));
    InMux I__12172 (
            .O(N__50994),
            .I(N__50978));
    Odrv4 I__12171 (
            .O(N__50989),
            .I(comm_rx_buf_5));
    Odrv4 I__12170 (
            .O(N__50984),
            .I(comm_rx_buf_5));
    LocalMux I__12169 (
            .O(N__50981),
            .I(comm_rx_buf_5));
    LocalMux I__12168 (
            .O(N__50978),
            .I(comm_rx_buf_5));
    CascadeMux I__12167 (
            .O(N__50969),
            .I(N__50965));
    InMux I__12166 (
            .O(N__50968),
            .I(N__50960));
    InMux I__12165 (
            .O(N__50965),
            .I(N__50960));
    LocalMux I__12164 (
            .O(N__50960),
            .I(comm_buf_6_5));
    CascadeMux I__12163 (
            .O(N__50957),
            .I(n2369_cascade_));
    CascadeMux I__12162 (
            .O(N__50954),
            .I(n21130_cascade_));
    CEMux I__12161 (
            .O(N__50951),
            .I(N__50948));
    LocalMux I__12160 (
            .O(N__50948),
            .I(N__50945));
    Odrv4 I__12159 (
            .O(N__50945),
            .I(n14_adj_1506));
    InMux I__12158 (
            .O(N__50942),
            .I(N__50939));
    LocalMux I__12157 (
            .O(N__50939),
            .I(N__50936));
    Odrv4 I__12156 (
            .O(N__50936),
            .I(n3));
    CascadeMux I__12155 (
            .O(N__50933),
            .I(N__50927));
    InMux I__12154 (
            .O(N__50932),
            .I(N__50922));
    InMux I__12153 (
            .O(N__50931),
            .I(N__50917));
    InMux I__12152 (
            .O(N__50930),
            .I(N__50917));
    InMux I__12151 (
            .O(N__50927),
            .I(N__50914));
    InMux I__12150 (
            .O(N__50926),
            .I(N__50911));
    InMux I__12149 (
            .O(N__50925),
            .I(N__50908));
    LocalMux I__12148 (
            .O(N__50922),
            .I(N__50903));
    LocalMux I__12147 (
            .O(N__50917),
            .I(N__50898));
    LocalMux I__12146 (
            .O(N__50914),
            .I(N__50898));
    LocalMux I__12145 (
            .O(N__50911),
            .I(N__50895));
    LocalMux I__12144 (
            .O(N__50908),
            .I(N__50892));
    InMux I__12143 (
            .O(N__50907),
            .I(N__50887));
    InMux I__12142 (
            .O(N__50906),
            .I(N__50887));
    Span4Mux_h I__12141 (
            .O(N__50903),
            .I(N__50882));
    Span4Mux_v I__12140 (
            .O(N__50898),
            .I(N__50879));
    Span4Mux_h I__12139 (
            .O(N__50895),
            .I(N__50872));
    Span4Mux_h I__12138 (
            .O(N__50892),
            .I(N__50872));
    LocalMux I__12137 (
            .O(N__50887),
            .I(N__50872));
    InMux I__12136 (
            .O(N__50886),
            .I(N__50867));
    InMux I__12135 (
            .O(N__50885),
            .I(N__50867));
    Odrv4 I__12134 (
            .O(N__50882),
            .I(n20681));
    Odrv4 I__12133 (
            .O(N__50879),
            .I(n20681));
    Odrv4 I__12132 (
            .O(N__50872),
            .I(n20681));
    LocalMux I__12131 (
            .O(N__50867),
            .I(n20681));
    CascadeMux I__12130 (
            .O(N__50858),
            .I(n3_cascade_));
    InMux I__12129 (
            .O(N__50855),
            .I(N__50851));
    InMux I__12128 (
            .O(N__50854),
            .I(N__50847));
    LocalMux I__12127 (
            .O(N__50851),
            .I(N__50844));
    InMux I__12126 (
            .O(N__50850),
            .I(N__50841));
    LocalMux I__12125 (
            .O(N__50847),
            .I(n2369));
    Odrv4 I__12124 (
            .O(N__50844),
            .I(n2369));
    LocalMux I__12123 (
            .O(N__50841),
            .I(n2369));
    InMux I__12122 (
            .O(N__50834),
            .I(N__50831));
    LocalMux I__12121 (
            .O(N__50831),
            .I(n19655));
    InMux I__12120 (
            .O(N__50828),
            .I(N__50825));
    LocalMux I__12119 (
            .O(N__50825),
            .I(n23_adj_1501));
    CascadeMux I__12118 (
            .O(N__50822),
            .I(n21_adj_1600_cascade_));
    InMux I__12117 (
            .O(N__50819),
            .I(N__50816));
    LocalMux I__12116 (
            .O(N__50816),
            .I(n17485));
    CEMux I__12115 (
            .O(N__50813),
            .I(N__50810));
    LocalMux I__12114 (
            .O(N__50810),
            .I(N__50807));
    Odrv12 I__12113 (
            .O(N__50807),
            .I(n18_adj_1633));
    CascadeMux I__12112 (
            .O(N__50804),
            .I(\comm_spi.imosi_cascade_ ));
    InMux I__12111 (
            .O(N__50801),
            .I(N__50798));
    LocalMux I__12110 (
            .O(N__50798),
            .I(\comm_spi.n22667 ));
    InMux I__12109 (
            .O(N__50795),
            .I(N__50792));
    LocalMux I__12108 (
            .O(N__50792),
            .I(N__50789));
    Odrv4 I__12107 (
            .O(N__50789),
            .I(\comm_spi.n14630 ));
    CascadeMux I__12106 (
            .O(N__50786),
            .I(\comm_spi.n22667_cascade_ ));
    InMux I__12105 (
            .O(N__50783),
            .I(N__50779));
    InMux I__12104 (
            .O(N__50782),
            .I(N__50772));
    LocalMux I__12103 (
            .O(N__50779),
            .I(N__50768));
    InMux I__12102 (
            .O(N__50778),
            .I(N__50765));
    InMux I__12101 (
            .O(N__50777),
            .I(N__50762));
    InMux I__12100 (
            .O(N__50776),
            .I(N__50758));
    InMux I__12099 (
            .O(N__50775),
            .I(N__50755));
    LocalMux I__12098 (
            .O(N__50772),
            .I(N__50752));
    InMux I__12097 (
            .O(N__50771),
            .I(N__50749));
    Span4Mux_h I__12096 (
            .O(N__50768),
            .I(N__50742));
    LocalMux I__12095 (
            .O(N__50765),
            .I(N__50742));
    LocalMux I__12094 (
            .O(N__50762),
            .I(N__50742));
    InMux I__12093 (
            .O(N__50761),
            .I(N__50739));
    LocalMux I__12092 (
            .O(N__50758),
            .I(N__50736));
    LocalMux I__12091 (
            .O(N__50755),
            .I(N__50733));
    Span4Mux_v I__12090 (
            .O(N__50752),
            .I(N__50728));
    LocalMux I__12089 (
            .O(N__50749),
            .I(N__50728));
    Span4Mux_v I__12088 (
            .O(N__50742),
            .I(N__50723));
    LocalMux I__12087 (
            .O(N__50739),
            .I(N__50723));
    Span12Mux_h I__12086 (
            .O(N__50736),
            .I(N__50720));
    Span4Mux_v I__12085 (
            .O(N__50733),
            .I(N__50715));
    Span4Mux_v I__12084 (
            .O(N__50728),
            .I(N__50715));
    Span4Mux_h I__12083 (
            .O(N__50723),
            .I(N__50712));
    Odrv12 I__12082 (
            .O(N__50720),
            .I(comm_rx_buf_0));
    Odrv4 I__12081 (
            .O(N__50715),
            .I(comm_rx_buf_0));
    Odrv4 I__12080 (
            .O(N__50712),
            .I(comm_rx_buf_0));
    CascadeMux I__12079 (
            .O(N__50705),
            .I(comm_rx_buf_0_cascade_));
    InMux I__12078 (
            .O(N__50702),
            .I(N__50698));
    InMux I__12077 (
            .O(N__50701),
            .I(N__50695));
    LocalMux I__12076 (
            .O(N__50698),
            .I(N__50692));
    LocalMux I__12075 (
            .O(N__50695),
            .I(comm_buf_6_0));
    Odrv12 I__12074 (
            .O(N__50692),
            .I(comm_buf_6_0));
    InMux I__12073 (
            .O(N__50687),
            .I(N__50671));
    InMux I__12072 (
            .O(N__50686),
            .I(N__50671));
    InMux I__12071 (
            .O(N__50685),
            .I(N__50671));
    InMux I__12070 (
            .O(N__50684),
            .I(N__50659));
    InMux I__12069 (
            .O(N__50683),
            .I(N__50652));
    InMux I__12068 (
            .O(N__50682),
            .I(N__50652));
    InMux I__12067 (
            .O(N__50681),
            .I(N__50652));
    InMux I__12066 (
            .O(N__50680),
            .I(N__50645));
    InMux I__12065 (
            .O(N__50679),
            .I(N__50645));
    InMux I__12064 (
            .O(N__50678),
            .I(N__50645));
    LocalMux I__12063 (
            .O(N__50671),
            .I(N__50642));
    InMux I__12062 (
            .O(N__50670),
            .I(N__50637));
    InMux I__12061 (
            .O(N__50669),
            .I(N__50637));
    CascadeMux I__12060 (
            .O(N__50668),
            .I(N__50633));
    InMux I__12059 (
            .O(N__50667),
            .I(N__50626));
    InMux I__12058 (
            .O(N__50666),
            .I(N__50626));
    InMux I__12057 (
            .O(N__50665),
            .I(N__50619));
    InMux I__12056 (
            .O(N__50664),
            .I(N__50619));
    InMux I__12055 (
            .O(N__50663),
            .I(N__50619));
    InMux I__12054 (
            .O(N__50662),
            .I(N__50616));
    LocalMux I__12053 (
            .O(N__50659),
            .I(N__50613));
    LocalMux I__12052 (
            .O(N__50652),
            .I(N__50604));
    LocalMux I__12051 (
            .O(N__50645),
            .I(N__50604));
    Span4Mux_v I__12050 (
            .O(N__50642),
            .I(N__50604));
    LocalMux I__12049 (
            .O(N__50637),
            .I(N__50604));
    InMux I__12048 (
            .O(N__50636),
            .I(N__50601));
    InMux I__12047 (
            .O(N__50633),
            .I(N__50598));
    InMux I__12046 (
            .O(N__50632),
            .I(N__50593));
    InMux I__12045 (
            .O(N__50631),
            .I(N__50593));
    LocalMux I__12044 (
            .O(N__50626),
            .I(N__50590));
    LocalMux I__12043 (
            .O(N__50619),
            .I(N__50585));
    LocalMux I__12042 (
            .O(N__50616),
            .I(N__50585));
    Span4Mux_v I__12041 (
            .O(N__50613),
            .I(N__50580));
    Span4Mux_h I__12040 (
            .O(N__50604),
            .I(N__50580));
    LocalMux I__12039 (
            .O(N__50601),
            .I(comm_index_2));
    LocalMux I__12038 (
            .O(N__50598),
            .I(comm_index_2));
    LocalMux I__12037 (
            .O(N__50593),
            .I(comm_index_2));
    Odrv4 I__12036 (
            .O(N__50590),
            .I(comm_index_2));
    Odrv4 I__12035 (
            .O(N__50585),
            .I(comm_index_2));
    Odrv4 I__12034 (
            .O(N__50580),
            .I(comm_index_2));
    InMux I__12033 (
            .O(N__50567),
            .I(N__50564));
    LocalMux I__12032 (
            .O(N__50564),
            .I(N__50561));
    Span4Mux_h I__12031 (
            .O(N__50561),
            .I(N__50558));
    Odrv4 I__12030 (
            .O(N__50558),
            .I(comm_buf_2_5));
    CascadeMux I__12029 (
            .O(N__50555),
            .I(N__50549));
    InMux I__12028 (
            .O(N__50554),
            .I(N__50539));
    InMux I__12027 (
            .O(N__50553),
            .I(N__50539));
    InMux I__12026 (
            .O(N__50552),
            .I(N__50529));
    InMux I__12025 (
            .O(N__50549),
            .I(N__50526));
    InMux I__12024 (
            .O(N__50548),
            .I(N__50523));
    InMux I__12023 (
            .O(N__50547),
            .I(N__50518));
    InMux I__12022 (
            .O(N__50546),
            .I(N__50518));
    InMux I__12021 (
            .O(N__50545),
            .I(N__50513));
    InMux I__12020 (
            .O(N__50544),
            .I(N__50513));
    LocalMux I__12019 (
            .O(N__50539),
            .I(N__50510));
    InMux I__12018 (
            .O(N__50538),
            .I(N__50507));
    InMux I__12017 (
            .O(N__50537),
            .I(N__50499));
    InMux I__12016 (
            .O(N__50536),
            .I(N__50499));
    InMux I__12015 (
            .O(N__50535),
            .I(N__50499));
    InMux I__12014 (
            .O(N__50534),
            .I(N__50496));
    InMux I__12013 (
            .O(N__50533),
            .I(N__50488));
    InMux I__12012 (
            .O(N__50532),
            .I(N__50488));
    LocalMux I__12011 (
            .O(N__50529),
            .I(N__50485));
    LocalMux I__12010 (
            .O(N__50526),
            .I(N__50478));
    LocalMux I__12009 (
            .O(N__50523),
            .I(N__50475));
    LocalMux I__12008 (
            .O(N__50518),
            .I(N__50466));
    LocalMux I__12007 (
            .O(N__50513),
            .I(N__50466));
    Span4Mux_v I__12006 (
            .O(N__50510),
            .I(N__50466));
    LocalMux I__12005 (
            .O(N__50507),
            .I(N__50466));
    InMux I__12004 (
            .O(N__50506),
            .I(N__50463));
    LocalMux I__12003 (
            .O(N__50499),
            .I(N__50458));
    LocalMux I__12002 (
            .O(N__50496),
            .I(N__50458));
    InMux I__12001 (
            .O(N__50495),
            .I(N__50451));
    InMux I__12000 (
            .O(N__50494),
            .I(N__50451));
    InMux I__11999 (
            .O(N__50493),
            .I(N__50451));
    LocalMux I__11998 (
            .O(N__50488),
            .I(N__50448));
    Span4Mux_h I__11997 (
            .O(N__50485),
            .I(N__50445));
    InMux I__11996 (
            .O(N__50484),
            .I(N__50436));
    InMux I__11995 (
            .O(N__50483),
            .I(N__50436));
    InMux I__11994 (
            .O(N__50482),
            .I(N__50436));
    InMux I__11993 (
            .O(N__50481),
            .I(N__50436));
    Span4Mux_h I__11992 (
            .O(N__50478),
            .I(N__50429));
    Span4Mux_h I__11991 (
            .O(N__50475),
            .I(N__50429));
    Span4Mux_h I__11990 (
            .O(N__50466),
            .I(N__50429));
    LocalMux I__11989 (
            .O(N__50463),
            .I(comm_index_1));
    Odrv4 I__11988 (
            .O(N__50458),
            .I(comm_index_1));
    LocalMux I__11987 (
            .O(N__50451),
            .I(comm_index_1));
    Odrv12 I__11986 (
            .O(N__50448),
            .I(comm_index_1));
    Odrv4 I__11985 (
            .O(N__50445),
            .I(comm_index_1));
    LocalMux I__11984 (
            .O(N__50436),
            .I(comm_index_1));
    Odrv4 I__11983 (
            .O(N__50429),
            .I(comm_index_1));
    InMux I__11982 (
            .O(N__50414),
            .I(N__50411));
    LocalMux I__11981 (
            .O(N__50411),
            .I(N__50408));
    Odrv12 I__11980 (
            .O(N__50408),
            .I(n22172));
    SRMux I__11979 (
            .O(N__50405),
            .I(N__50402));
    LocalMux I__11978 (
            .O(N__50402),
            .I(N__50399));
    Odrv4 I__11977 (
            .O(N__50399),
            .I(n14671));
    InMux I__11976 (
            .O(N__50396),
            .I(N__50393));
    LocalMux I__11975 (
            .O(N__50393),
            .I(\SIG_DDS.n21331 ));
    CascadeMux I__11974 (
            .O(N__50390),
            .I(N__50387));
    InMux I__11973 (
            .O(N__50387),
            .I(N__50384));
    LocalMux I__11972 (
            .O(N__50384),
            .I(\SIG_DDS.n10 ));
    CEMux I__11971 (
            .O(N__50381),
            .I(N__50377));
    CEMux I__11970 (
            .O(N__50380),
            .I(N__50374));
    LocalMux I__11969 (
            .O(N__50377),
            .I(N__50371));
    LocalMux I__11968 (
            .O(N__50374),
            .I(\SIG_DDS.n9 ));
    Odrv4 I__11967 (
            .O(N__50371),
            .I(\SIG_DDS.n9 ));
    InMux I__11966 (
            .O(N__50366),
            .I(N__50363));
    LocalMux I__11965 (
            .O(N__50363),
            .I(N__50355));
    CascadeMux I__11964 (
            .O(N__50362),
            .I(N__50350));
    InMux I__11963 (
            .O(N__50361),
            .I(N__50346));
    InMux I__11962 (
            .O(N__50360),
            .I(N__50343));
    InMux I__11961 (
            .O(N__50359),
            .I(N__50340));
    InMux I__11960 (
            .O(N__50358),
            .I(N__50337));
    Span12Mux_s8_v I__11959 (
            .O(N__50355),
            .I(N__50334));
    InMux I__11958 (
            .O(N__50354),
            .I(N__50329));
    InMux I__11957 (
            .O(N__50353),
            .I(N__50329));
    InMux I__11956 (
            .O(N__50350),
            .I(N__50324));
    InMux I__11955 (
            .O(N__50349),
            .I(N__50324));
    LocalMux I__11954 (
            .O(N__50346),
            .I(dds_state_0));
    LocalMux I__11953 (
            .O(N__50343),
            .I(dds_state_0));
    LocalMux I__11952 (
            .O(N__50340),
            .I(dds_state_0));
    LocalMux I__11951 (
            .O(N__50337),
            .I(dds_state_0));
    Odrv12 I__11950 (
            .O(N__50334),
            .I(dds_state_0));
    LocalMux I__11949 (
            .O(N__50329),
            .I(dds_state_0));
    LocalMux I__11948 (
            .O(N__50324),
            .I(dds_state_0));
    InMux I__11947 (
            .O(N__50309),
            .I(N__50278));
    InMux I__11946 (
            .O(N__50308),
            .I(N__50278));
    InMux I__11945 (
            .O(N__50307),
            .I(N__50278));
    InMux I__11944 (
            .O(N__50306),
            .I(N__50278));
    InMux I__11943 (
            .O(N__50305),
            .I(N__50278));
    InMux I__11942 (
            .O(N__50304),
            .I(N__50278));
    InMux I__11941 (
            .O(N__50303),
            .I(N__50278));
    InMux I__11940 (
            .O(N__50302),
            .I(N__50278));
    InMux I__11939 (
            .O(N__50301),
            .I(N__50263));
    InMux I__11938 (
            .O(N__50300),
            .I(N__50263));
    InMux I__11937 (
            .O(N__50299),
            .I(N__50263));
    InMux I__11936 (
            .O(N__50298),
            .I(N__50263));
    InMux I__11935 (
            .O(N__50297),
            .I(N__50263));
    InMux I__11934 (
            .O(N__50296),
            .I(N__50263));
    InMux I__11933 (
            .O(N__50295),
            .I(N__50263));
    LocalMux I__11932 (
            .O(N__50278),
            .I(N__50255));
    LocalMux I__11931 (
            .O(N__50263),
            .I(N__50255));
    InMux I__11930 (
            .O(N__50262),
            .I(N__50251));
    InMux I__11929 (
            .O(N__50261),
            .I(N__50243));
    InMux I__11928 (
            .O(N__50260),
            .I(N__50243));
    Span4Mux_v I__11927 (
            .O(N__50255),
            .I(N__50240));
    InMux I__11926 (
            .O(N__50254),
            .I(N__50237));
    LocalMux I__11925 (
            .O(N__50251),
            .I(N__50234));
    InMux I__11924 (
            .O(N__50250),
            .I(N__50230));
    InMux I__11923 (
            .O(N__50249),
            .I(N__50225));
    InMux I__11922 (
            .O(N__50248),
            .I(N__50225));
    LocalMux I__11921 (
            .O(N__50243),
            .I(N__50220));
    Span4Mux_h I__11920 (
            .O(N__50240),
            .I(N__50213));
    LocalMux I__11919 (
            .O(N__50237),
            .I(N__50213));
    Span4Mux_v I__11918 (
            .O(N__50234),
            .I(N__50213));
    InMux I__11917 (
            .O(N__50233),
            .I(N__50210));
    LocalMux I__11916 (
            .O(N__50230),
            .I(N__50205));
    LocalMux I__11915 (
            .O(N__50225),
            .I(N__50205));
    InMux I__11914 (
            .O(N__50224),
            .I(N__50200));
    InMux I__11913 (
            .O(N__50223),
            .I(N__50200));
    Span4Mux_v I__11912 (
            .O(N__50220),
            .I(N__50197));
    Odrv4 I__11911 (
            .O(N__50213),
            .I(dds_state_2));
    LocalMux I__11910 (
            .O(N__50210),
            .I(dds_state_2));
    Odrv12 I__11909 (
            .O(N__50205),
            .I(dds_state_2));
    LocalMux I__11908 (
            .O(N__50200),
            .I(dds_state_2));
    Odrv4 I__11907 (
            .O(N__50197),
            .I(dds_state_2));
    SRMux I__11906 (
            .O(N__50186),
            .I(N__50173));
    InMux I__11905 (
            .O(N__50185),
            .I(N__50158));
    InMux I__11904 (
            .O(N__50184),
            .I(N__50158));
    InMux I__11903 (
            .O(N__50183),
            .I(N__50158));
    InMux I__11902 (
            .O(N__50182),
            .I(N__50158));
    InMux I__11901 (
            .O(N__50181),
            .I(N__50158));
    InMux I__11900 (
            .O(N__50180),
            .I(N__50158));
    InMux I__11899 (
            .O(N__50179),
            .I(N__50158));
    InMux I__11898 (
            .O(N__50178),
            .I(N__50151));
    InMux I__11897 (
            .O(N__50177),
            .I(N__50151));
    CEMux I__11896 (
            .O(N__50176),
            .I(N__50148));
    LocalMux I__11895 (
            .O(N__50173),
            .I(N__50145));
    LocalMux I__11894 (
            .O(N__50158),
            .I(N__50142));
    CascadeMux I__11893 (
            .O(N__50157),
            .I(N__50134));
    InMux I__11892 (
            .O(N__50156),
            .I(N__50127));
    LocalMux I__11891 (
            .O(N__50151),
            .I(N__50124));
    LocalMux I__11890 (
            .O(N__50148),
            .I(N__50121));
    Span4Mux_v I__11889 (
            .O(N__50145),
            .I(N__50116));
    Span4Mux_h I__11888 (
            .O(N__50142),
            .I(N__50116));
    InMux I__11887 (
            .O(N__50141),
            .I(N__50099));
    InMux I__11886 (
            .O(N__50140),
            .I(N__50099));
    InMux I__11885 (
            .O(N__50139),
            .I(N__50099));
    InMux I__11884 (
            .O(N__50138),
            .I(N__50099));
    InMux I__11883 (
            .O(N__50137),
            .I(N__50099));
    InMux I__11882 (
            .O(N__50134),
            .I(N__50099));
    InMux I__11881 (
            .O(N__50133),
            .I(N__50099));
    InMux I__11880 (
            .O(N__50132),
            .I(N__50099));
    InMux I__11879 (
            .O(N__50131),
            .I(N__50095));
    InMux I__11878 (
            .O(N__50130),
            .I(N__50092));
    LocalMux I__11877 (
            .O(N__50127),
            .I(N__50087));
    Span4Mux_h I__11876 (
            .O(N__50124),
            .I(N__50087));
    Span4Mux_h I__11875 (
            .O(N__50121),
            .I(N__50077));
    Span4Mux_h I__11874 (
            .O(N__50116),
            .I(N__50077));
    LocalMux I__11873 (
            .O(N__50099),
            .I(N__50074));
    InMux I__11872 (
            .O(N__50098),
            .I(N__50071));
    LocalMux I__11871 (
            .O(N__50095),
            .I(N__50064));
    LocalMux I__11870 (
            .O(N__50092),
            .I(N__50064));
    Span4Mux_h I__11869 (
            .O(N__50087),
            .I(N__50064));
    InMux I__11868 (
            .O(N__50086),
            .I(N__50057));
    InMux I__11867 (
            .O(N__50085),
            .I(N__50057));
    InMux I__11866 (
            .O(N__50084),
            .I(N__50057));
    InMux I__11865 (
            .O(N__50083),
            .I(N__50052));
    InMux I__11864 (
            .O(N__50082),
            .I(N__50052));
    Odrv4 I__11863 (
            .O(N__50077),
            .I(dds_state_1));
    Odrv12 I__11862 (
            .O(N__50074),
            .I(dds_state_1));
    LocalMux I__11861 (
            .O(N__50071),
            .I(dds_state_1));
    Odrv4 I__11860 (
            .O(N__50064),
            .I(dds_state_1));
    LocalMux I__11859 (
            .O(N__50057),
            .I(dds_state_1));
    LocalMux I__11858 (
            .O(N__50052),
            .I(dds_state_1));
    IoInMux I__11857 (
            .O(N__50039),
            .I(N__50036));
    LocalMux I__11856 (
            .O(N__50036),
            .I(N__50033));
    IoSpan4Mux I__11855 (
            .O(N__50033),
            .I(N__50030));
    IoSpan4Mux I__11854 (
            .O(N__50030),
            .I(N__50027));
    Span4Mux_s3_v I__11853 (
            .O(N__50027),
            .I(N__50023));
    CascadeMux I__11852 (
            .O(N__50026),
            .I(N__50020));
    Span4Mux_v I__11851 (
            .O(N__50023),
            .I(N__50017));
    InMux I__11850 (
            .O(N__50020),
            .I(N__50014));
    Odrv4 I__11849 (
            .O(N__50017),
            .I(DDS_SCK));
    LocalMux I__11848 (
            .O(N__50014),
            .I(DDS_SCK));
    InMux I__11847 (
            .O(N__50009),
            .I(N__50006));
    LocalMux I__11846 (
            .O(N__50006),
            .I(N__50003));
    Span4Mux_v I__11845 (
            .O(N__50003),
            .I(N__49999));
    InMux I__11844 (
            .O(N__50002),
            .I(N__49995));
    Sp12to4 I__11843 (
            .O(N__49999),
            .I(N__49992));
    InMux I__11842 (
            .O(N__49998),
            .I(N__49989));
    LocalMux I__11841 (
            .O(N__49995),
            .I(N__49986));
    Odrv12 I__11840 (
            .O(N__49992),
            .I(wdtick_flag));
    LocalMux I__11839 (
            .O(N__49989),
            .I(wdtick_flag));
    Odrv4 I__11838 (
            .O(N__49986),
            .I(wdtick_flag));
    InMux I__11837 (
            .O(N__49979),
            .I(N__49975));
    InMux I__11836 (
            .O(N__49978),
            .I(N__49972));
    LocalMux I__11835 (
            .O(N__49975),
            .I(N__49968));
    LocalMux I__11834 (
            .O(N__49972),
            .I(N__49965));
    InMux I__11833 (
            .O(N__49971),
            .I(N__49962));
    Span4Mux_v I__11832 (
            .O(N__49968),
            .I(N__49959));
    Odrv4 I__11831 (
            .O(N__49965),
            .I(buf_control_0));
    LocalMux I__11830 (
            .O(N__49962),
            .I(buf_control_0));
    Odrv4 I__11829 (
            .O(N__49959),
            .I(buf_control_0));
    IoInMux I__11828 (
            .O(N__49952),
            .I(N__49949));
    LocalMux I__11827 (
            .O(N__49949),
            .I(N__49946));
    IoSpan4Mux I__11826 (
            .O(N__49946),
            .I(N__49943));
    Span4Mux_s3_v I__11825 (
            .O(N__49943),
            .I(N__49940));
    Span4Mux_v I__11824 (
            .O(N__49940),
            .I(N__49937));
    Odrv4 I__11823 (
            .O(N__49937),
            .I(CONT_SD));
    InMux I__11822 (
            .O(N__49934),
            .I(N__49931));
    LocalMux I__11821 (
            .O(N__49931),
            .I(N__49928));
    Odrv4 I__11820 (
            .O(N__49928),
            .I(n20608));
    CascadeMux I__11819 (
            .O(N__49925),
            .I(N__49911));
    CascadeMux I__11818 (
            .O(N__49924),
            .I(N__49905));
    CascadeMux I__11817 (
            .O(N__49923),
            .I(N__49901));
    InMux I__11816 (
            .O(N__49922),
            .I(N__49890));
    InMux I__11815 (
            .O(N__49921),
            .I(N__49890));
    InMux I__11814 (
            .O(N__49920),
            .I(N__49887));
    InMux I__11813 (
            .O(N__49919),
            .I(N__49882));
    InMux I__11812 (
            .O(N__49918),
            .I(N__49882));
    CascadeMux I__11811 (
            .O(N__49917),
            .I(N__49879));
    CascadeMux I__11810 (
            .O(N__49916),
            .I(N__49876));
    CascadeMux I__11809 (
            .O(N__49915),
            .I(N__49872));
    InMux I__11808 (
            .O(N__49914),
            .I(N__49868));
    InMux I__11807 (
            .O(N__49911),
            .I(N__49861));
    InMux I__11806 (
            .O(N__49910),
            .I(N__49861));
    InMux I__11805 (
            .O(N__49909),
            .I(N__49861));
    InMux I__11804 (
            .O(N__49908),
            .I(N__49856));
    InMux I__11803 (
            .O(N__49905),
            .I(N__49856));
    InMux I__11802 (
            .O(N__49904),
            .I(N__49849));
    InMux I__11801 (
            .O(N__49901),
            .I(N__49849));
    InMux I__11800 (
            .O(N__49900),
            .I(N__49849));
    InMux I__11799 (
            .O(N__49899),
            .I(N__49840));
    InMux I__11798 (
            .O(N__49898),
            .I(N__49840));
    InMux I__11797 (
            .O(N__49897),
            .I(N__49840));
    InMux I__11796 (
            .O(N__49896),
            .I(N__49840));
    CascadeMux I__11795 (
            .O(N__49895),
            .I(N__49835));
    LocalMux I__11794 (
            .O(N__49890),
            .I(N__49820));
    LocalMux I__11793 (
            .O(N__49887),
            .I(N__49815));
    LocalMux I__11792 (
            .O(N__49882),
            .I(N__49815));
    InMux I__11791 (
            .O(N__49879),
            .I(N__49810));
    InMux I__11790 (
            .O(N__49876),
            .I(N__49810));
    InMux I__11789 (
            .O(N__49875),
            .I(N__49803));
    InMux I__11788 (
            .O(N__49872),
            .I(N__49803));
    InMux I__11787 (
            .O(N__49871),
            .I(N__49803));
    LocalMux I__11786 (
            .O(N__49868),
            .I(N__49792));
    LocalMux I__11785 (
            .O(N__49861),
            .I(N__49792));
    LocalMux I__11784 (
            .O(N__49856),
            .I(N__49792));
    LocalMux I__11783 (
            .O(N__49849),
            .I(N__49792));
    LocalMux I__11782 (
            .O(N__49840),
            .I(N__49792));
    InMux I__11781 (
            .O(N__49839),
            .I(N__49785));
    InMux I__11780 (
            .O(N__49838),
            .I(N__49785));
    InMux I__11779 (
            .O(N__49835),
            .I(N__49785));
    InMux I__11778 (
            .O(N__49834),
            .I(N__49782));
    CascadeMux I__11777 (
            .O(N__49833),
            .I(N__49777));
    CascadeMux I__11776 (
            .O(N__49832),
            .I(N__49768));
    InMux I__11775 (
            .O(N__49831),
            .I(N__49762));
    InMux I__11774 (
            .O(N__49830),
            .I(N__49762));
    CascadeMux I__11773 (
            .O(N__49829),
            .I(N__49759));
    InMux I__11772 (
            .O(N__49828),
            .I(N__49755));
    CascadeMux I__11771 (
            .O(N__49827),
            .I(N__49751));
    CascadeMux I__11770 (
            .O(N__49826),
            .I(N__49746));
    CascadeMux I__11769 (
            .O(N__49825),
            .I(N__49743));
    CascadeMux I__11768 (
            .O(N__49824),
            .I(N__49740));
    CascadeMux I__11767 (
            .O(N__49823),
            .I(N__49736));
    Span4Mux_h I__11766 (
            .O(N__49820),
            .I(N__49721));
    Span4Mux_v I__11765 (
            .O(N__49815),
            .I(N__49721));
    LocalMux I__11764 (
            .O(N__49810),
            .I(N__49721));
    LocalMux I__11763 (
            .O(N__49803),
            .I(N__49721));
    Span4Mux_v I__11762 (
            .O(N__49792),
            .I(N__49721));
    LocalMux I__11761 (
            .O(N__49785),
            .I(N__49721));
    LocalMux I__11760 (
            .O(N__49782),
            .I(N__49717));
    InMux I__11759 (
            .O(N__49781),
            .I(N__49714));
    CascadeMux I__11758 (
            .O(N__49780),
            .I(N__49711));
    InMux I__11757 (
            .O(N__49777),
            .I(N__49705));
    InMux I__11756 (
            .O(N__49776),
            .I(N__49702));
    CascadeMux I__11755 (
            .O(N__49775),
            .I(N__49695));
    CascadeMux I__11754 (
            .O(N__49774),
            .I(N__49692));
    CascadeMux I__11753 (
            .O(N__49773),
            .I(N__49688));
    CascadeMux I__11752 (
            .O(N__49772),
            .I(N__49683));
    CascadeMux I__11751 (
            .O(N__49771),
            .I(N__49679));
    InMux I__11750 (
            .O(N__49768),
            .I(N__49674));
    InMux I__11749 (
            .O(N__49767),
            .I(N__49674));
    LocalMux I__11748 (
            .O(N__49762),
            .I(N__49671));
    InMux I__11747 (
            .O(N__49759),
            .I(N__49668));
    CascadeMux I__11746 (
            .O(N__49758),
            .I(N__49665));
    LocalMux I__11745 (
            .O(N__49755),
            .I(N__49660));
    InMux I__11744 (
            .O(N__49754),
            .I(N__49657));
    InMux I__11743 (
            .O(N__49751),
            .I(N__49652));
    InMux I__11742 (
            .O(N__49750),
            .I(N__49652));
    InMux I__11741 (
            .O(N__49749),
            .I(N__49647));
    InMux I__11740 (
            .O(N__49746),
            .I(N__49647));
    InMux I__11739 (
            .O(N__49743),
            .I(N__49642));
    InMux I__11738 (
            .O(N__49740),
            .I(N__49642));
    InMux I__11737 (
            .O(N__49739),
            .I(N__49639));
    InMux I__11736 (
            .O(N__49736),
            .I(N__49631));
    InMux I__11735 (
            .O(N__49735),
            .I(N__49631));
    InMux I__11734 (
            .O(N__49734),
            .I(N__49631));
    Span4Mux_v I__11733 (
            .O(N__49721),
            .I(N__49623));
    InMux I__11732 (
            .O(N__49720),
            .I(N__49620));
    Span4Mux_v I__11731 (
            .O(N__49717),
            .I(N__49617));
    LocalMux I__11730 (
            .O(N__49714),
            .I(N__49614));
    InMux I__11729 (
            .O(N__49711),
            .I(N__49605));
    InMux I__11728 (
            .O(N__49710),
            .I(N__49605));
    InMux I__11727 (
            .O(N__49709),
            .I(N__49605));
    InMux I__11726 (
            .O(N__49708),
            .I(N__49605));
    LocalMux I__11725 (
            .O(N__49705),
            .I(N__49602));
    LocalMux I__11724 (
            .O(N__49702),
            .I(N__49599));
    CascadeMux I__11723 (
            .O(N__49701),
            .I(N__49596));
    CascadeMux I__11722 (
            .O(N__49700),
            .I(N__49587));
    InMux I__11721 (
            .O(N__49699),
            .I(N__49576));
    InMux I__11720 (
            .O(N__49698),
            .I(N__49576));
    InMux I__11719 (
            .O(N__49695),
            .I(N__49576));
    InMux I__11718 (
            .O(N__49692),
            .I(N__49576));
    InMux I__11717 (
            .O(N__49691),
            .I(N__49576));
    InMux I__11716 (
            .O(N__49688),
            .I(N__49569));
    InMux I__11715 (
            .O(N__49687),
            .I(N__49569));
    InMux I__11714 (
            .O(N__49686),
            .I(N__49569));
    InMux I__11713 (
            .O(N__49683),
            .I(N__49562));
    InMux I__11712 (
            .O(N__49682),
            .I(N__49562));
    InMux I__11711 (
            .O(N__49679),
            .I(N__49562));
    LocalMux I__11710 (
            .O(N__49674),
            .I(N__49555));
    Span4Mux_h I__11709 (
            .O(N__49671),
            .I(N__49555));
    LocalMux I__11708 (
            .O(N__49668),
            .I(N__49555));
    InMux I__11707 (
            .O(N__49665),
            .I(N__49548));
    InMux I__11706 (
            .O(N__49664),
            .I(N__49548));
    InMux I__11705 (
            .O(N__49663),
            .I(N__49548));
    Span4Mux_v I__11704 (
            .O(N__49660),
            .I(N__49539));
    LocalMux I__11703 (
            .O(N__49657),
            .I(N__49539));
    LocalMux I__11702 (
            .O(N__49652),
            .I(N__49539));
    LocalMux I__11701 (
            .O(N__49647),
            .I(N__49539));
    LocalMux I__11700 (
            .O(N__49642),
            .I(N__49536));
    LocalMux I__11699 (
            .O(N__49639),
            .I(N__49533));
    InMux I__11698 (
            .O(N__49638),
            .I(N__49530));
    LocalMux I__11697 (
            .O(N__49631),
            .I(N__49527));
    InMux I__11696 (
            .O(N__49630),
            .I(N__49524));
    CascadeMux I__11695 (
            .O(N__49629),
            .I(N__49518));
    InMux I__11694 (
            .O(N__49628),
            .I(N__49515));
    InMux I__11693 (
            .O(N__49627),
            .I(N__49512));
    InMux I__11692 (
            .O(N__49626),
            .I(N__49509));
    Span4Mux_h I__11691 (
            .O(N__49623),
            .I(N__49506));
    LocalMux I__11690 (
            .O(N__49620),
            .I(N__49497));
    Span4Mux_h I__11689 (
            .O(N__49617),
            .I(N__49497));
    Span4Mux_v I__11688 (
            .O(N__49614),
            .I(N__49497));
    LocalMux I__11687 (
            .O(N__49605),
            .I(N__49497));
    Span4Mux_v I__11686 (
            .O(N__49602),
            .I(N__49492));
    Span4Mux_v I__11685 (
            .O(N__49599),
            .I(N__49492));
    InMux I__11684 (
            .O(N__49596),
            .I(N__49489));
    InMux I__11683 (
            .O(N__49595),
            .I(N__49482));
    InMux I__11682 (
            .O(N__49594),
            .I(N__49482));
    InMux I__11681 (
            .O(N__49593),
            .I(N__49482));
    InMux I__11680 (
            .O(N__49592),
            .I(N__49473));
    InMux I__11679 (
            .O(N__49591),
            .I(N__49473));
    InMux I__11678 (
            .O(N__49590),
            .I(N__49473));
    InMux I__11677 (
            .O(N__49587),
            .I(N__49473));
    LocalMux I__11676 (
            .O(N__49576),
            .I(N__49462));
    LocalMux I__11675 (
            .O(N__49569),
            .I(N__49462));
    LocalMux I__11674 (
            .O(N__49562),
            .I(N__49462));
    Span4Mux_v I__11673 (
            .O(N__49555),
            .I(N__49462));
    LocalMux I__11672 (
            .O(N__49548),
            .I(N__49462));
    Span4Mux_v I__11671 (
            .O(N__49539),
            .I(N__49457));
    Span4Mux_v I__11670 (
            .O(N__49536),
            .I(N__49457));
    Span4Mux_h I__11669 (
            .O(N__49533),
            .I(N__49450));
    LocalMux I__11668 (
            .O(N__49530),
            .I(N__49450));
    Span4Mux_h I__11667 (
            .O(N__49527),
            .I(N__49450));
    LocalMux I__11666 (
            .O(N__49524),
            .I(N__49445));
    InMux I__11665 (
            .O(N__49523),
            .I(N__49436));
    InMux I__11664 (
            .O(N__49522),
            .I(N__49436));
    InMux I__11663 (
            .O(N__49521),
            .I(N__49436));
    InMux I__11662 (
            .O(N__49518),
            .I(N__49436));
    LocalMux I__11661 (
            .O(N__49515),
            .I(N__49433));
    LocalMux I__11660 (
            .O(N__49512),
            .I(N__49428));
    LocalMux I__11659 (
            .O(N__49509),
            .I(N__49428));
    Span4Mux_h I__11658 (
            .O(N__49506),
            .I(N__49423));
    Span4Mux_v I__11657 (
            .O(N__49497),
            .I(N__49423));
    Span4Mux_v I__11656 (
            .O(N__49492),
            .I(N__49418));
    LocalMux I__11655 (
            .O(N__49489),
            .I(N__49418));
    LocalMux I__11654 (
            .O(N__49482),
            .I(N__49407));
    LocalMux I__11653 (
            .O(N__49473),
            .I(N__49407));
    Span4Mux_h I__11652 (
            .O(N__49462),
            .I(N__49407));
    Span4Mux_h I__11651 (
            .O(N__49457),
            .I(N__49407));
    Span4Mux_h I__11650 (
            .O(N__49450),
            .I(N__49407));
    InMux I__11649 (
            .O(N__49449),
            .I(N__49404));
    InMux I__11648 (
            .O(N__49448),
            .I(N__49401));
    Sp12to4 I__11647 (
            .O(N__49445),
            .I(N__49396));
    LocalMux I__11646 (
            .O(N__49436),
            .I(N__49396));
    Span4Mux_h I__11645 (
            .O(N__49433),
            .I(N__49389));
    Span4Mux_v I__11644 (
            .O(N__49428),
            .I(N__49389));
    Span4Mux_v I__11643 (
            .O(N__49423),
            .I(N__49389));
    Span4Mux_h I__11642 (
            .O(N__49418),
            .I(N__49384));
    Span4Mux_v I__11641 (
            .O(N__49407),
            .I(N__49384));
    LocalMux I__11640 (
            .O(N__49404),
            .I(n9321));
    LocalMux I__11639 (
            .O(N__49401),
            .I(n9321));
    Odrv12 I__11638 (
            .O(N__49396),
            .I(n9321));
    Odrv4 I__11637 (
            .O(N__49389),
            .I(n9321));
    Odrv4 I__11636 (
            .O(N__49384),
            .I(n9321));
    InMux I__11635 (
            .O(N__49373),
            .I(N__49363));
    InMux I__11634 (
            .O(N__49372),
            .I(N__49360));
    InMux I__11633 (
            .O(N__49371),
            .I(N__49345));
    InMux I__11632 (
            .O(N__49370),
            .I(N__49345));
    InMux I__11631 (
            .O(N__49369),
            .I(N__49345));
    InMux I__11630 (
            .O(N__49368),
            .I(N__49345));
    InMux I__11629 (
            .O(N__49367),
            .I(N__49345));
    InMux I__11628 (
            .O(N__49366),
            .I(N__49339));
    LocalMux I__11627 (
            .O(N__49363),
            .I(N__49336));
    LocalMux I__11626 (
            .O(N__49360),
            .I(N__49333));
    InMux I__11625 (
            .O(N__49359),
            .I(N__49326));
    InMux I__11624 (
            .O(N__49358),
            .I(N__49326));
    InMux I__11623 (
            .O(N__49357),
            .I(N__49326));
    InMux I__11622 (
            .O(N__49356),
            .I(N__49323));
    LocalMux I__11621 (
            .O(N__49345),
            .I(N__49320));
    InMux I__11620 (
            .O(N__49344),
            .I(N__49317));
    InMux I__11619 (
            .O(N__49343),
            .I(N__49312));
    InMux I__11618 (
            .O(N__49342),
            .I(N__49312));
    LocalMux I__11617 (
            .O(N__49339),
            .I(N__49309));
    Span4Mux_v I__11616 (
            .O(N__49336),
            .I(N__49306));
    Span4Mux_v I__11615 (
            .O(N__49333),
            .I(N__49303));
    LocalMux I__11614 (
            .O(N__49326),
            .I(N__49296));
    LocalMux I__11613 (
            .O(N__49323),
            .I(N__49296));
    Span4Mux_h I__11612 (
            .O(N__49320),
            .I(N__49296));
    LocalMux I__11611 (
            .O(N__49317),
            .I(n12441));
    LocalMux I__11610 (
            .O(N__49312),
            .I(n12441));
    Odrv4 I__11609 (
            .O(N__49309),
            .I(n12441));
    Odrv4 I__11608 (
            .O(N__49306),
            .I(n12441));
    Odrv4 I__11607 (
            .O(N__49303),
            .I(n12441));
    Odrv4 I__11606 (
            .O(N__49296),
            .I(n12441));
    InMux I__11605 (
            .O(N__49283),
            .I(N__49279));
    InMux I__11604 (
            .O(N__49282),
            .I(N__49276));
    LocalMux I__11603 (
            .O(N__49279),
            .I(N__49272));
    LocalMux I__11602 (
            .O(N__49276),
            .I(N__49269));
    InMux I__11601 (
            .O(N__49275),
            .I(N__49266));
    Span4Mux_h I__11600 (
            .O(N__49272),
            .I(N__49263));
    Span4Mux_h I__11599 (
            .O(N__49269),
            .I(N__49260));
    LocalMux I__11598 (
            .O(N__49266),
            .I(acadc_skipCount_4));
    Odrv4 I__11597 (
            .O(N__49263),
            .I(acadc_skipCount_4));
    Odrv4 I__11596 (
            .O(N__49260),
            .I(acadc_skipCount_4));
    InMux I__11595 (
            .O(N__49253),
            .I(N__49250));
    LocalMux I__11594 (
            .O(N__49250),
            .I(N__49246));
    CascadeMux I__11593 (
            .O(N__49249),
            .I(N__49243));
    Span4Mux_h I__11592 (
            .O(N__49246),
            .I(N__49240));
    InMux I__11591 (
            .O(N__49243),
            .I(N__49237));
    Span4Mux_v I__11590 (
            .O(N__49240),
            .I(N__49234));
    LocalMux I__11589 (
            .O(N__49237),
            .I(data_idxvec_7));
    Odrv4 I__11588 (
            .O(N__49234),
            .I(data_idxvec_7));
    InMux I__11587 (
            .O(N__49229),
            .I(N__49226));
    LocalMux I__11586 (
            .O(N__49226),
            .I(N__49221));
    InMux I__11585 (
            .O(N__49225),
            .I(N__49218));
    InMux I__11584 (
            .O(N__49224),
            .I(N__49215));
    Span4Mux_h I__11583 (
            .O(N__49221),
            .I(N__49212));
    LocalMux I__11582 (
            .O(N__49218),
            .I(data_cntvec_7));
    LocalMux I__11581 (
            .O(N__49215),
            .I(data_cntvec_7));
    Odrv4 I__11580 (
            .O(N__49212),
            .I(data_cntvec_7));
    InMux I__11579 (
            .O(N__49205),
            .I(N__49202));
    LocalMux I__11578 (
            .O(N__49202),
            .I(N__49199));
    Span4Mux_v I__11577 (
            .O(N__49199),
            .I(N__49196));
    Odrv4 I__11576 (
            .O(N__49196),
            .I(buf_data_iac_15));
    CascadeMux I__11575 (
            .O(N__49193),
            .I(n26_adj_1500_cascade_));
    CascadeMux I__11574 (
            .O(N__49190),
            .I(n20810_cascade_));
    InMux I__11573 (
            .O(N__49187),
            .I(N__49184));
    LocalMux I__11572 (
            .O(N__49184),
            .I(n22058));
    CascadeMux I__11571 (
            .O(N__49181),
            .I(N__49177));
    InMux I__11570 (
            .O(N__49180),
            .I(N__49173));
    InMux I__11569 (
            .O(N__49177),
            .I(N__49170));
    InMux I__11568 (
            .O(N__49176),
            .I(N__49167));
    LocalMux I__11567 (
            .O(N__49173),
            .I(N__49162));
    LocalMux I__11566 (
            .O(N__49170),
            .I(N__49162));
    LocalMux I__11565 (
            .O(N__49167),
            .I(acadc_skipCount_7));
    Odrv12 I__11564 (
            .O(N__49162),
            .I(acadc_skipCount_7));
    CascadeMux I__11563 (
            .O(N__49157),
            .I(N__49154));
    InMux I__11562 (
            .O(N__49154),
            .I(N__49149));
    InMux I__11561 (
            .O(N__49153),
            .I(N__49146));
    InMux I__11560 (
            .O(N__49152),
            .I(N__49143));
    LocalMux I__11559 (
            .O(N__49149),
            .I(N__49140));
    LocalMux I__11558 (
            .O(N__49146),
            .I(req_data_cnt_7));
    LocalMux I__11557 (
            .O(N__49143),
            .I(req_data_cnt_7));
    Odrv4 I__11556 (
            .O(N__49140),
            .I(req_data_cnt_7));
    InMux I__11555 (
            .O(N__49133),
            .I(N__49130));
    LocalMux I__11554 (
            .O(N__49130),
            .I(n20809));
    CascadeMux I__11553 (
            .O(N__49127),
            .I(N__49095));
    InMux I__11552 (
            .O(N__49126),
            .I(N__49092));
    InMux I__11551 (
            .O(N__49125),
            .I(N__49089));
    InMux I__11550 (
            .O(N__49124),
            .I(N__49086));
    InMux I__11549 (
            .O(N__49123),
            .I(N__49079));
    InMux I__11548 (
            .O(N__49122),
            .I(N__49079));
    InMux I__11547 (
            .O(N__49121),
            .I(N__49079));
    InMux I__11546 (
            .O(N__49120),
            .I(N__49069));
    InMux I__11545 (
            .O(N__49119),
            .I(N__49069));
    InMux I__11544 (
            .O(N__49118),
            .I(N__49066));
    InMux I__11543 (
            .O(N__49117),
            .I(N__49063));
    InMux I__11542 (
            .O(N__49116),
            .I(N__49060));
    InMux I__11541 (
            .O(N__49115),
            .I(N__49046));
    InMux I__11540 (
            .O(N__49114),
            .I(N__49039));
    InMux I__11539 (
            .O(N__49113),
            .I(N__49039));
    InMux I__11538 (
            .O(N__49112),
            .I(N__49039));
    InMux I__11537 (
            .O(N__49111),
            .I(N__49030));
    InMux I__11536 (
            .O(N__49110),
            .I(N__49030));
    InMux I__11535 (
            .O(N__49109),
            .I(N__49030));
    InMux I__11534 (
            .O(N__49108),
            .I(N__49030));
    InMux I__11533 (
            .O(N__49107),
            .I(N__49021));
    InMux I__11532 (
            .O(N__49106),
            .I(N__49021));
    InMux I__11531 (
            .O(N__49105),
            .I(N__49021));
    InMux I__11530 (
            .O(N__49104),
            .I(N__49021));
    InMux I__11529 (
            .O(N__49103),
            .I(N__49014));
    InMux I__11528 (
            .O(N__49102),
            .I(N__49014));
    InMux I__11527 (
            .O(N__49101),
            .I(N__49014));
    InMux I__11526 (
            .O(N__49100),
            .I(N__49007));
    InMux I__11525 (
            .O(N__49099),
            .I(N__49004));
    InMux I__11524 (
            .O(N__49098),
            .I(N__49000));
    InMux I__11523 (
            .O(N__49095),
            .I(N__48994));
    LocalMux I__11522 (
            .O(N__49092),
            .I(N__48991));
    LocalMux I__11521 (
            .O(N__49089),
            .I(N__48984));
    LocalMux I__11520 (
            .O(N__49086),
            .I(N__48984));
    LocalMux I__11519 (
            .O(N__49079),
            .I(N__48984));
    InMux I__11518 (
            .O(N__49078),
            .I(N__48977));
    InMux I__11517 (
            .O(N__49077),
            .I(N__48977));
    InMux I__11516 (
            .O(N__49076),
            .I(N__48977));
    InMux I__11515 (
            .O(N__49075),
            .I(N__48974));
    InMux I__11514 (
            .O(N__49074),
            .I(N__48971));
    LocalMux I__11513 (
            .O(N__49069),
            .I(N__48966));
    LocalMux I__11512 (
            .O(N__49066),
            .I(N__48966));
    LocalMux I__11511 (
            .O(N__49063),
            .I(N__48961));
    LocalMux I__11510 (
            .O(N__49060),
            .I(N__48961));
    InMux I__11509 (
            .O(N__49059),
            .I(N__48958));
    InMux I__11508 (
            .O(N__49058),
            .I(N__48955));
    InMux I__11507 (
            .O(N__49057),
            .I(N__48946));
    InMux I__11506 (
            .O(N__49056),
            .I(N__48946));
    InMux I__11505 (
            .O(N__49055),
            .I(N__48941));
    InMux I__11504 (
            .O(N__49054),
            .I(N__48941));
    InMux I__11503 (
            .O(N__49053),
            .I(N__48938));
    InMux I__11502 (
            .O(N__49052),
            .I(N__48935));
    InMux I__11501 (
            .O(N__49051),
            .I(N__48928));
    InMux I__11500 (
            .O(N__49050),
            .I(N__48928));
    InMux I__11499 (
            .O(N__49049),
            .I(N__48928));
    LocalMux I__11498 (
            .O(N__49046),
            .I(N__48919));
    LocalMux I__11497 (
            .O(N__49039),
            .I(N__48919));
    LocalMux I__11496 (
            .O(N__49030),
            .I(N__48919));
    LocalMux I__11495 (
            .O(N__49021),
            .I(N__48919));
    LocalMux I__11494 (
            .O(N__49014),
            .I(N__48916));
    InMux I__11493 (
            .O(N__49013),
            .I(N__48911));
    InMux I__11492 (
            .O(N__49012),
            .I(N__48911));
    InMux I__11491 (
            .O(N__49011),
            .I(N__48906));
    InMux I__11490 (
            .O(N__49010),
            .I(N__48906));
    LocalMux I__11489 (
            .O(N__49007),
            .I(N__48903));
    LocalMux I__11488 (
            .O(N__49004),
            .I(N__48900));
    InMux I__11487 (
            .O(N__49003),
            .I(N__48897));
    LocalMux I__11486 (
            .O(N__49000),
            .I(N__48894));
    InMux I__11485 (
            .O(N__48999),
            .I(N__48887));
    InMux I__11484 (
            .O(N__48998),
            .I(N__48887));
    InMux I__11483 (
            .O(N__48997),
            .I(N__48887));
    LocalMux I__11482 (
            .O(N__48994),
            .I(N__48880));
    Span4Mux_v I__11481 (
            .O(N__48991),
            .I(N__48880));
    Span4Mux_v I__11480 (
            .O(N__48984),
            .I(N__48880));
    LocalMux I__11479 (
            .O(N__48977),
            .I(N__48877));
    LocalMux I__11478 (
            .O(N__48974),
            .I(N__48870));
    LocalMux I__11477 (
            .O(N__48971),
            .I(N__48865));
    Span4Mux_v I__11476 (
            .O(N__48966),
            .I(N__48865));
    Span4Mux_v I__11475 (
            .O(N__48961),
            .I(N__48860));
    LocalMux I__11474 (
            .O(N__48958),
            .I(N__48860));
    LocalMux I__11473 (
            .O(N__48955),
            .I(N__48857));
    InMux I__11472 (
            .O(N__48954),
            .I(N__48853));
    InMux I__11471 (
            .O(N__48953),
            .I(N__48846));
    InMux I__11470 (
            .O(N__48952),
            .I(N__48846));
    InMux I__11469 (
            .O(N__48951),
            .I(N__48846));
    LocalMux I__11468 (
            .O(N__48946),
            .I(N__48841));
    LocalMux I__11467 (
            .O(N__48941),
            .I(N__48841));
    LocalMux I__11466 (
            .O(N__48938),
            .I(N__48838));
    LocalMux I__11465 (
            .O(N__48935),
            .I(N__48835));
    LocalMux I__11464 (
            .O(N__48928),
            .I(N__48826));
    Span4Mux_v I__11463 (
            .O(N__48919),
            .I(N__48826));
    Span4Mux_h I__11462 (
            .O(N__48916),
            .I(N__48826));
    LocalMux I__11461 (
            .O(N__48911),
            .I(N__48826));
    LocalMux I__11460 (
            .O(N__48906),
            .I(N__48817));
    Span4Mux_h I__11459 (
            .O(N__48903),
            .I(N__48817));
    Span4Mux_h I__11458 (
            .O(N__48900),
            .I(N__48817));
    LocalMux I__11457 (
            .O(N__48897),
            .I(N__48817));
    Span4Mux_v I__11456 (
            .O(N__48894),
            .I(N__48810));
    LocalMux I__11455 (
            .O(N__48887),
            .I(N__48810));
    Span4Mux_h I__11454 (
            .O(N__48880),
            .I(N__48807));
    Span12Mux_h I__11453 (
            .O(N__48877),
            .I(N__48804));
    InMux I__11452 (
            .O(N__48876),
            .I(N__48795));
    InMux I__11451 (
            .O(N__48875),
            .I(N__48795));
    InMux I__11450 (
            .O(N__48874),
            .I(N__48795));
    InMux I__11449 (
            .O(N__48873),
            .I(N__48795));
    Span4Mux_v I__11448 (
            .O(N__48870),
            .I(N__48786));
    Span4Mux_v I__11447 (
            .O(N__48865),
            .I(N__48786));
    Span4Mux_v I__11446 (
            .O(N__48860),
            .I(N__48786));
    Span4Mux_v I__11445 (
            .O(N__48857),
            .I(N__48786));
    InMux I__11444 (
            .O(N__48856),
            .I(N__48783));
    LocalMux I__11443 (
            .O(N__48853),
            .I(N__48776));
    LocalMux I__11442 (
            .O(N__48846),
            .I(N__48776));
    Span12Mux_v I__11441 (
            .O(N__48841),
            .I(N__48776));
    Span4Mux_h I__11440 (
            .O(N__48838),
            .I(N__48767));
    Span4Mux_v I__11439 (
            .O(N__48835),
            .I(N__48767));
    Span4Mux_h I__11438 (
            .O(N__48826),
            .I(N__48767));
    Span4Mux_v I__11437 (
            .O(N__48817),
            .I(N__48767));
    InMux I__11436 (
            .O(N__48816),
            .I(N__48762));
    InMux I__11435 (
            .O(N__48815),
            .I(N__48762));
    Odrv4 I__11434 (
            .O(N__48810),
            .I(comm_cmd_2));
    Odrv4 I__11433 (
            .O(N__48807),
            .I(comm_cmd_2));
    Odrv12 I__11432 (
            .O(N__48804),
            .I(comm_cmd_2));
    LocalMux I__11431 (
            .O(N__48795),
            .I(comm_cmd_2));
    Odrv4 I__11430 (
            .O(N__48786),
            .I(comm_cmd_2));
    LocalMux I__11429 (
            .O(N__48783),
            .I(comm_cmd_2));
    Odrv12 I__11428 (
            .O(N__48776),
            .I(comm_cmd_2));
    Odrv4 I__11427 (
            .O(N__48767),
            .I(comm_cmd_2));
    LocalMux I__11426 (
            .O(N__48762),
            .I(comm_cmd_2));
    CascadeMux I__11425 (
            .O(N__48743),
            .I(N__48731));
    InMux I__11424 (
            .O(N__48742),
            .I(N__48724));
    CascadeMux I__11423 (
            .O(N__48741),
            .I(N__48720));
    InMux I__11422 (
            .O(N__48740),
            .I(N__48715));
    InMux I__11421 (
            .O(N__48739),
            .I(N__48709));
    InMux I__11420 (
            .O(N__48738),
            .I(N__48709));
    InMux I__11419 (
            .O(N__48737),
            .I(N__48704));
    InMux I__11418 (
            .O(N__48736),
            .I(N__48704));
    InMux I__11417 (
            .O(N__48735),
            .I(N__48697));
    InMux I__11416 (
            .O(N__48734),
            .I(N__48692));
    InMux I__11415 (
            .O(N__48731),
            .I(N__48692));
    InMux I__11414 (
            .O(N__48730),
            .I(N__48689));
    InMux I__11413 (
            .O(N__48729),
            .I(N__48682));
    CascadeMux I__11412 (
            .O(N__48728),
            .I(N__48678));
    InMux I__11411 (
            .O(N__48727),
            .I(N__48673));
    LocalMux I__11410 (
            .O(N__48724),
            .I(N__48670));
    InMux I__11409 (
            .O(N__48723),
            .I(N__48665));
    InMux I__11408 (
            .O(N__48720),
            .I(N__48662));
    InMux I__11407 (
            .O(N__48719),
            .I(N__48659));
    CascadeMux I__11406 (
            .O(N__48718),
            .I(N__48656));
    LocalMux I__11405 (
            .O(N__48715),
            .I(N__48653));
    InMux I__11404 (
            .O(N__48714),
            .I(N__48650));
    LocalMux I__11403 (
            .O(N__48709),
            .I(N__48645));
    LocalMux I__11402 (
            .O(N__48704),
            .I(N__48645));
    InMux I__11401 (
            .O(N__48703),
            .I(N__48642));
    InMux I__11400 (
            .O(N__48702),
            .I(N__48639));
    InMux I__11399 (
            .O(N__48701),
            .I(N__48636));
    InMux I__11398 (
            .O(N__48700),
            .I(N__48633));
    LocalMux I__11397 (
            .O(N__48697),
            .I(N__48626));
    LocalMux I__11396 (
            .O(N__48692),
            .I(N__48626));
    LocalMux I__11395 (
            .O(N__48689),
            .I(N__48626));
    InMux I__11394 (
            .O(N__48688),
            .I(N__48621));
    InMux I__11393 (
            .O(N__48687),
            .I(N__48621));
    InMux I__11392 (
            .O(N__48686),
            .I(N__48614));
    InMux I__11391 (
            .O(N__48685),
            .I(N__48614));
    LocalMux I__11390 (
            .O(N__48682),
            .I(N__48611));
    InMux I__11389 (
            .O(N__48681),
            .I(N__48608));
    InMux I__11388 (
            .O(N__48678),
            .I(N__48602));
    InMux I__11387 (
            .O(N__48677),
            .I(N__48602));
    InMux I__11386 (
            .O(N__48676),
            .I(N__48599));
    LocalMux I__11385 (
            .O(N__48673),
            .I(N__48594));
    Span4Mux_v I__11384 (
            .O(N__48670),
            .I(N__48591));
    InMux I__11383 (
            .O(N__48669),
            .I(N__48588));
    InMux I__11382 (
            .O(N__48668),
            .I(N__48585));
    LocalMux I__11381 (
            .O(N__48665),
            .I(N__48578));
    LocalMux I__11380 (
            .O(N__48662),
            .I(N__48578));
    LocalMux I__11379 (
            .O(N__48659),
            .I(N__48578));
    InMux I__11378 (
            .O(N__48656),
            .I(N__48575));
    Span4Mux_h I__11377 (
            .O(N__48653),
            .I(N__48569));
    LocalMux I__11376 (
            .O(N__48650),
            .I(N__48569));
    Span4Mux_h I__11375 (
            .O(N__48645),
            .I(N__48564));
    LocalMux I__11374 (
            .O(N__48642),
            .I(N__48564));
    LocalMux I__11373 (
            .O(N__48639),
            .I(N__48553));
    LocalMux I__11372 (
            .O(N__48636),
            .I(N__48553));
    LocalMux I__11371 (
            .O(N__48633),
            .I(N__48553));
    Span4Mux_v I__11370 (
            .O(N__48626),
            .I(N__48553));
    LocalMux I__11369 (
            .O(N__48621),
            .I(N__48553));
    CascadeMux I__11368 (
            .O(N__48620),
            .I(N__48550));
    InMux I__11367 (
            .O(N__48619),
            .I(N__48547));
    LocalMux I__11366 (
            .O(N__48614),
            .I(N__48544));
    Span4Mux_v I__11365 (
            .O(N__48611),
            .I(N__48539));
    LocalMux I__11364 (
            .O(N__48608),
            .I(N__48539));
    InMux I__11363 (
            .O(N__48607),
            .I(N__48533));
    LocalMux I__11362 (
            .O(N__48602),
            .I(N__48528));
    LocalMux I__11361 (
            .O(N__48599),
            .I(N__48528));
    InMux I__11360 (
            .O(N__48598),
            .I(N__48523));
    InMux I__11359 (
            .O(N__48597),
            .I(N__48523));
    Span4Mux_h I__11358 (
            .O(N__48594),
            .I(N__48518));
    Span4Mux_v I__11357 (
            .O(N__48591),
            .I(N__48518));
    LocalMux I__11356 (
            .O(N__48588),
            .I(N__48515));
    LocalMux I__11355 (
            .O(N__48585),
            .I(N__48510));
    Span4Mux_h I__11354 (
            .O(N__48578),
            .I(N__48510));
    LocalMux I__11353 (
            .O(N__48575),
            .I(N__48507));
    InMux I__11352 (
            .O(N__48574),
            .I(N__48504));
    Span4Mux_v I__11351 (
            .O(N__48569),
            .I(N__48496));
    Span4Mux_v I__11350 (
            .O(N__48564),
            .I(N__48496));
    Span4Mux_h I__11349 (
            .O(N__48553),
            .I(N__48496));
    InMux I__11348 (
            .O(N__48550),
            .I(N__48493));
    LocalMux I__11347 (
            .O(N__48547),
            .I(N__48488));
    Span4Mux_v I__11346 (
            .O(N__48544),
            .I(N__48488));
    Span4Mux_h I__11345 (
            .O(N__48539),
            .I(N__48485));
    InMux I__11344 (
            .O(N__48538),
            .I(N__48482));
    InMux I__11343 (
            .O(N__48537),
            .I(N__48477));
    InMux I__11342 (
            .O(N__48536),
            .I(N__48477));
    LocalMux I__11341 (
            .O(N__48533),
            .I(N__48468));
    Span12Mux_v I__11340 (
            .O(N__48528),
            .I(N__48468));
    LocalMux I__11339 (
            .O(N__48523),
            .I(N__48468));
    Sp12to4 I__11338 (
            .O(N__48518),
            .I(N__48468));
    Sp12to4 I__11337 (
            .O(N__48515),
            .I(N__48465));
    Span4Mux_v I__11336 (
            .O(N__48510),
            .I(N__48460));
    Span4Mux_h I__11335 (
            .O(N__48507),
            .I(N__48460));
    LocalMux I__11334 (
            .O(N__48504),
            .I(N__48457));
    InMux I__11333 (
            .O(N__48503),
            .I(N__48454));
    Span4Mux_h I__11332 (
            .O(N__48496),
            .I(N__48451));
    LocalMux I__11331 (
            .O(N__48493),
            .I(N__48440));
    Span4Mux_h I__11330 (
            .O(N__48488),
            .I(N__48440));
    Span4Mux_v I__11329 (
            .O(N__48485),
            .I(N__48440));
    LocalMux I__11328 (
            .O(N__48482),
            .I(N__48440));
    LocalMux I__11327 (
            .O(N__48477),
            .I(N__48440));
    Odrv12 I__11326 (
            .O(N__48468),
            .I(comm_cmd_3));
    Odrv12 I__11325 (
            .O(N__48465),
            .I(comm_cmd_3));
    Odrv4 I__11324 (
            .O(N__48460),
            .I(comm_cmd_3));
    Odrv12 I__11323 (
            .O(N__48457),
            .I(comm_cmd_3));
    LocalMux I__11322 (
            .O(N__48454),
            .I(comm_cmd_3));
    Odrv4 I__11321 (
            .O(N__48451),
            .I(comm_cmd_3));
    Odrv4 I__11320 (
            .O(N__48440),
            .I(comm_cmd_3));
    CascadeMux I__11319 (
            .O(N__48425),
            .I(N__48420));
    CascadeMux I__11318 (
            .O(N__48424),
            .I(N__48411));
    CascadeMux I__11317 (
            .O(N__48423),
            .I(N__48405));
    InMux I__11316 (
            .O(N__48420),
            .I(N__48402));
    InMux I__11315 (
            .O(N__48419),
            .I(N__48399));
    InMux I__11314 (
            .O(N__48418),
            .I(N__48395));
    InMux I__11313 (
            .O(N__48417),
            .I(N__48388));
    InMux I__11312 (
            .O(N__48416),
            .I(N__48388));
    InMux I__11311 (
            .O(N__48415),
            .I(N__48388));
    InMux I__11310 (
            .O(N__48414),
            .I(N__48385));
    InMux I__11309 (
            .O(N__48411),
            .I(N__48381));
    InMux I__11308 (
            .O(N__48410),
            .I(N__48378));
    CascadeMux I__11307 (
            .O(N__48409),
            .I(N__48366));
    InMux I__11306 (
            .O(N__48408),
            .I(N__48354));
    InMux I__11305 (
            .O(N__48405),
            .I(N__48354));
    LocalMux I__11304 (
            .O(N__48402),
            .I(N__48351));
    LocalMux I__11303 (
            .O(N__48399),
            .I(N__48348));
    InMux I__11302 (
            .O(N__48398),
            .I(N__48345));
    LocalMux I__11301 (
            .O(N__48395),
            .I(N__48328));
    LocalMux I__11300 (
            .O(N__48388),
            .I(N__48328));
    LocalMux I__11299 (
            .O(N__48385),
            .I(N__48328));
    InMux I__11298 (
            .O(N__48384),
            .I(N__48325));
    LocalMux I__11297 (
            .O(N__48381),
            .I(N__48322));
    LocalMux I__11296 (
            .O(N__48378),
            .I(N__48319));
    InMux I__11295 (
            .O(N__48377),
            .I(N__48305));
    InMux I__11294 (
            .O(N__48376),
            .I(N__48300));
    InMux I__11293 (
            .O(N__48375),
            .I(N__48300));
    InMux I__11292 (
            .O(N__48374),
            .I(N__48289));
    InMux I__11291 (
            .O(N__48373),
            .I(N__48286));
    InMux I__11290 (
            .O(N__48372),
            .I(N__48278));
    InMux I__11289 (
            .O(N__48371),
            .I(N__48278));
    InMux I__11288 (
            .O(N__48370),
            .I(N__48278));
    InMux I__11287 (
            .O(N__48369),
            .I(N__48273));
    InMux I__11286 (
            .O(N__48366),
            .I(N__48273));
    CascadeMux I__11285 (
            .O(N__48365),
            .I(N__48270));
    CascadeMux I__11284 (
            .O(N__48364),
            .I(N__48267));
    InMux I__11283 (
            .O(N__48363),
            .I(N__48259));
    InMux I__11282 (
            .O(N__48362),
            .I(N__48259));
    InMux I__11281 (
            .O(N__48361),
            .I(N__48259));
    InMux I__11280 (
            .O(N__48360),
            .I(N__48256));
    InMux I__11279 (
            .O(N__48359),
            .I(N__48253));
    LocalMux I__11278 (
            .O(N__48354),
            .I(N__48248));
    Span4Mux_v I__11277 (
            .O(N__48351),
            .I(N__48248));
    Span4Mux_v I__11276 (
            .O(N__48348),
            .I(N__48243));
    LocalMux I__11275 (
            .O(N__48345),
            .I(N__48243));
    InMux I__11274 (
            .O(N__48344),
            .I(N__48236));
    InMux I__11273 (
            .O(N__48343),
            .I(N__48236));
    InMux I__11272 (
            .O(N__48342),
            .I(N__48236));
    InMux I__11271 (
            .O(N__48341),
            .I(N__48233));
    InMux I__11270 (
            .O(N__48340),
            .I(N__48229));
    InMux I__11269 (
            .O(N__48339),
            .I(N__48223));
    InMux I__11268 (
            .O(N__48338),
            .I(N__48223));
    InMux I__11267 (
            .O(N__48337),
            .I(N__48218));
    InMux I__11266 (
            .O(N__48336),
            .I(N__48218));
    InMux I__11265 (
            .O(N__48335),
            .I(N__48212));
    Span4Mux_v I__11264 (
            .O(N__48328),
            .I(N__48203));
    LocalMux I__11263 (
            .O(N__48325),
            .I(N__48203));
    Span4Mux_h I__11262 (
            .O(N__48322),
            .I(N__48203));
    Span4Mux_h I__11261 (
            .O(N__48319),
            .I(N__48203));
    InMux I__11260 (
            .O(N__48318),
            .I(N__48196));
    InMux I__11259 (
            .O(N__48317),
            .I(N__48196));
    InMux I__11258 (
            .O(N__48316),
            .I(N__48196));
    InMux I__11257 (
            .O(N__48315),
            .I(N__48191));
    InMux I__11256 (
            .O(N__48314),
            .I(N__48188));
    InMux I__11255 (
            .O(N__48313),
            .I(N__48185));
    InMux I__11254 (
            .O(N__48312),
            .I(N__48180));
    InMux I__11253 (
            .O(N__48311),
            .I(N__48180));
    InMux I__11252 (
            .O(N__48310),
            .I(N__48177));
    InMux I__11251 (
            .O(N__48309),
            .I(N__48172));
    InMux I__11250 (
            .O(N__48308),
            .I(N__48172));
    LocalMux I__11249 (
            .O(N__48305),
            .I(N__48167));
    LocalMux I__11248 (
            .O(N__48300),
            .I(N__48164));
    InMux I__11247 (
            .O(N__48299),
            .I(N__48161));
    InMux I__11246 (
            .O(N__48298),
            .I(N__48154));
    InMux I__11245 (
            .O(N__48297),
            .I(N__48154));
    InMux I__11244 (
            .O(N__48296),
            .I(N__48154));
    InMux I__11243 (
            .O(N__48295),
            .I(N__48148));
    InMux I__11242 (
            .O(N__48294),
            .I(N__48141));
    InMux I__11241 (
            .O(N__48293),
            .I(N__48141));
    InMux I__11240 (
            .O(N__48292),
            .I(N__48141));
    LocalMux I__11239 (
            .O(N__48289),
            .I(N__48136));
    LocalMux I__11238 (
            .O(N__48286),
            .I(N__48136));
    InMux I__11237 (
            .O(N__48285),
            .I(N__48133));
    LocalMux I__11236 (
            .O(N__48278),
            .I(N__48128));
    LocalMux I__11235 (
            .O(N__48273),
            .I(N__48128));
    InMux I__11234 (
            .O(N__48270),
            .I(N__48123));
    InMux I__11233 (
            .O(N__48267),
            .I(N__48123));
    InMux I__11232 (
            .O(N__48266),
            .I(N__48120));
    LocalMux I__11231 (
            .O(N__48259),
            .I(N__48117));
    LocalMux I__11230 (
            .O(N__48256),
            .I(N__48114));
    LocalMux I__11229 (
            .O(N__48253),
            .I(N__48111));
    Span4Mux_h I__11228 (
            .O(N__48248),
            .I(N__48102));
    Span4Mux_v I__11227 (
            .O(N__48243),
            .I(N__48102));
    LocalMux I__11226 (
            .O(N__48236),
            .I(N__48102));
    LocalMux I__11225 (
            .O(N__48233),
            .I(N__48102));
    InMux I__11224 (
            .O(N__48232),
            .I(N__48099));
    LocalMux I__11223 (
            .O(N__48229),
            .I(N__48095));
    InMux I__11222 (
            .O(N__48228),
            .I(N__48091));
    LocalMux I__11221 (
            .O(N__48223),
            .I(N__48085));
    LocalMux I__11220 (
            .O(N__48218),
            .I(N__48085));
    InMux I__11219 (
            .O(N__48217),
            .I(N__48078));
    InMux I__11218 (
            .O(N__48216),
            .I(N__48078));
    InMux I__11217 (
            .O(N__48215),
            .I(N__48078));
    LocalMux I__11216 (
            .O(N__48212),
            .I(N__48073));
    Span4Mux_h I__11215 (
            .O(N__48203),
            .I(N__48073));
    LocalMux I__11214 (
            .O(N__48196),
            .I(N__48070));
    InMux I__11213 (
            .O(N__48195),
            .I(N__48065));
    InMux I__11212 (
            .O(N__48194),
            .I(N__48065));
    LocalMux I__11211 (
            .O(N__48191),
            .I(N__48054));
    LocalMux I__11210 (
            .O(N__48188),
            .I(N__48054));
    LocalMux I__11209 (
            .O(N__48185),
            .I(N__48054));
    LocalMux I__11208 (
            .O(N__48180),
            .I(N__48054));
    LocalMux I__11207 (
            .O(N__48177),
            .I(N__48054));
    LocalMux I__11206 (
            .O(N__48172),
            .I(N__48051));
    InMux I__11205 (
            .O(N__48171),
            .I(N__48046));
    InMux I__11204 (
            .O(N__48170),
            .I(N__48046));
    Span4Mux_v I__11203 (
            .O(N__48167),
            .I(N__48037));
    Span4Mux_h I__11202 (
            .O(N__48164),
            .I(N__48037));
    LocalMux I__11201 (
            .O(N__48161),
            .I(N__48037));
    LocalMux I__11200 (
            .O(N__48154),
            .I(N__48037));
    InMux I__11199 (
            .O(N__48153),
            .I(N__48030));
    InMux I__11198 (
            .O(N__48152),
            .I(N__48030));
    InMux I__11197 (
            .O(N__48151),
            .I(N__48030));
    LocalMux I__11196 (
            .O(N__48148),
            .I(N__48027));
    LocalMux I__11195 (
            .O(N__48141),
            .I(N__48024));
    Span4Mux_v I__11194 (
            .O(N__48136),
            .I(N__48021));
    LocalMux I__11193 (
            .O(N__48133),
            .I(N__48014));
    Span4Mux_v I__11192 (
            .O(N__48128),
            .I(N__48014));
    LocalMux I__11191 (
            .O(N__48123),
            .I(N__48014));
    LocalMux I__11190 (
            .O(N__48120),
            .I(N__48011));
    Span4Mux_h I__11189 (
            .O(N__48117),
            .I(N__48008));
    Span4Mux_h I__11188 (
            .O(N__48114),
            .I(N__47999));
    Span4Mux_h I__11187 (
            .O(N__48111),
            .I(N__47999));
    Span4Mux_h I__11186 (
            .O(N__48102),
            .I(N__47999));
    LocalMux I__11185 (
            .O(N__48099),
            .I(N__47999));
    InMux I__11184 (
            .O(N__48098),
            .I(N__47994));
    Span4Mux_h I__11183 (
            .O(N__48095),
            .I(N__47991));
    InMux I__11182 (
            .O(N__48094),
            .I(N__47988));
    LocalMux I__11181 (
            .O(N__48091),
            .I(N__47985));
    InMux I__11180 (
            .O(N__48090),
            .I(N__47982));
    Span4Mux_h I__11179 (
            .O(N__48085),
            .I(N__47975));
    LocalMux I__11178 (
            .O(N__48078),
            .I(N__47975));
    Span4Mux_v I__11177 (
            .O(N__48073),
            .I(N__47975));
    Span4Mux_h I__11176 (
            .O(N__48070),
            .I(N__47970));
    LocalMux I__11175 (
            .O(N__48065),
            .I(N__47970));
    Span4Mux_v I__11174 (
            .O(N__48054),
            .I(N__47961));
    Span4Mux_v I__11173 (
            .O(N__48051),
            .I(N__47961));
    LocalMux I__11172 (
            .O(N__48046),
            .I(N__47961));
    Span4Mux_v I__11171 (
            .O(N__48037),
            .I(N__47961));
    LocalMux I__11170 (
            .O(N__48030),
            .I(N__47950));
    Span4Mux_v I__11169 (
            .O(N__48027),
            .I(N__47950));
    Span4Mux_v I__11168 (
            .O(N__48024),
            .I(N__47950));
    Span4Mux_h I__11167 (
            .O(N__48021),
            .I(N__47950));
    Span4Mux_v I__11166 (
            .O(N__48014),
            .I(N__47950));
    Span4Mux_v I__11165 (
            .O(N__48011),
            .I(N__47943));
    Span4Mux_v I__11164 (
            .O(N__48008),
            .I(N__47943));
    Span4Mux_v I__11163 (
            .O(N__47999),
            .I(N__47943));
    InMux I__11162 (
            .O(N__47998),
            .I(N__47938));
    InMux I__11161 (
            .O(N__47997),
            .I(N__47938));
    LocalMux I__11160 (
            .O(N__47994),
            .I(comm_cmd_1));
    Odrv4 I__11159 (
            .O(N__47991),
            .I(comm_cmd_1));
    LocalMux I__11158 (
            .O(N__47988),
            .I(comm_cmd_1));
    Odrv12 I__11157 (
            .O(N__47985),
            .I(comm_cmd_1));
    LocalMux I__11156 (
            .O(N__47982),
            .I(comm_cmd_1));
    Odrv4 I__11155 (
            .O(N__47975),
            .I(comm_cmd_1));
    Odrv4 I__11154 (
            .O(N__47970),
            .I(comm_cmd_1));
    Odrv4 I__11153 (
            .O(N__47961),
            .I(comm_cmd_1));
    Odrv4 I__11152 (
            .O(N__47950),
            .I(comm_cmd_1));
    Odrv4 I__11151 (
            .O(N__47943),
            .I(comm_cmd_1));
    LocalMux I__11150 (
            .O(N__47938),
            .I(comm_cmd_1));
    CascadeMux I__11149 (
            .O(N__47915),
            .I(N__47912));
    InMux I__11148 (
            .O(N__47912),
            .I(N__47908));
    InMux I__11147 (
            .O(N__47911),
            .I(N__47905));
    LocalMux I__11146 (
            .O(N__47908),
            .I(N__47902));
    LocalMux I__11145 (
            .O(N__47905),
            .I(N__47899));
    Span4Mux_v I__11144 (
            .O(N__47902),
            .I(N__47894));
    Span4Mux_h I__11143 (
            .O(N__47899),
            .I(N__47894));
    Span4Mux_v I__11142 (
            .O(N__47894),
            .I(N__47891));
    Odrv4 I__11141 (
            .O(N__47891),
            .I(comm_length_1));
    InMux I__11140 (
            .O(N__47888),
            .I(N__47884));
    InMux I__11139 (
            .O(N__47887),
            .I(N__47881));
    LocalMux I__11138 (
            .O(N__47884),
            .I(comm_length_2));
    LocalMux I__11137 (
            .O(N__47881),
            .I(comm_length_2));
    CascadeMux I__11136 (
            .O(N__47876),
            .I(N__47873));
    InMux I__11135 (
            .O(N__47873),
            .I(N__47870));
    LocalMux I__11134 (
            .O(N__47870),
            .I(comm_length_0));
    InMux I__11133 (
            .O(N__47867),
            .I(N__47863));
    InMux I__11132 (
            .O(N__47866),
            .I(N__47860));
    LocalMux I__11131 (
            .O(N__47863),
            .I(N__47857));
    LocalMux I__11130 (
            .O(N__47860),
            .I(N__47854));
    Span4Mux_v I__11129 (
            .O(N__47857),
            .I(N__47851));
    Span12Mux_v I__11128 (
            .O(N__47854),
            .I(N__47848));
    Odrv4 I__11127 (
            .O(N__47851),
            .I(n4));
    Odrv12 I__11126 (
            .O(N__47848),
            .I(n4));
    InMux I__11125 (
            .O(N__47843),
            .I(N__47838));
    InMux I__11124 (
            .O(N__47842),
            .I(N__47835));
    CascadeMux I__11123 (
            .O(N__47841),
            .I(N__47832));
    LocalMux I__11122 (
            .O(N__47838),
            .I(N__47829));
    LocalMux I__11121 (
            .O(N__47835),
            .I(N__47826));
    InMux I__11120 (
            .O(N__47832),
            .I(N__47823));
    Span4Mux_v I__11119 (
            .O(N__47829),
            .I(N__47818));
    Span4Mux_h I__11118 (
            .O(N__47826),
            .I(N__47818));
    LocalMux I__11117 (
            .O(N__47823),
            .I(N__47815));
    Span4Mux_h I__11116 (
            .O(N__47818),
            .I(N__47812));
    Span4Mux_h I__11115 (
            .O(N__47815),
            .I(N__47809));
    Span4Mux_h I__11114 (
            .O(N__47812),
            .I(N__47806));
    Span4Mux_v I__11113 (
            .O(N__47809),
            .I(N__47803));
    Span4Mux_v I__11112 (
            .O(N__47806),
            .I(N__47800));
    Odrv4 I__11111 (
            .O(N__47803),
            .I(n14_adj_1579));
    Odrv4 I__11110 (
            .O(N__47800),
            .I(n14_adj_1579));
    CascadeMux I__11109 (
            .O(N__47795),
            .I(N__47791));
    InMux I__11108 (
            .O(N__47794),
            .I(N__47788));
    InMux I__11107 (
            .O(N__47791),
            .I(N__47784));
    LocalMux I__11106 (
            .O(N__47788),
            .I(N__47781));
    CascadeMux I__11105 (
            .O(N__47787),
            .I(N__47778));
    LocalMux I__11104 (
            .O(N__47784),
            .I(N__47773));
    Span4Mux_h I__11103 (
            .O(N__47781),
            .I(N__47773));
    InMux I__11102 (
            .O(N__47778),
            .I(N__47770));
    Odrv4 I__11101 (
            .O(N__47773),
            .I(acadc_skipCount_15));
    LocalMux I__11100 (
            .O(N__47770),
            .I(acadc_skipCount_15));
    CascadeMux I__11099 (
            .O(N__47765),
            .I(N__47762));
    InMux I__11098 (
            .O(N__47762),
            .I(N__47759));
    LocalMux I__11097 (
            .O(N__47759),
            .I(N__47756));
    Odrv12 I__11096 (
            .O(N__47756),
            .I(n23_adj_1527));
    InMux I__11095 (
            .O(N__47753),
            .I(N__47749));
    InMux I__11094 (
            .O(N__47752),
            .I(N__47746));
    LocalMux I__11093 (
            .O(N__47749),
            .I(N__47740));
    LocalMux I__11092 (
            .O(N__47746),
            .I(N__47740));
    InMux I__11091 (
            .O(N__47745),
            .I(N__47737));
    Odrv12 I__11090 (
            .O(N__47740),
            .I(data_cntvec_5));
    LocalMux I__11089 (
            .O(N__47737),
            .I(data_cntvec_5));
    InMux I__11088 (
            .O(N__47732),
            .I(N__47727));
    InMux I__11087 (
            .O(N__47731),
            .I(N__47724));
    InMux I__11086 (
            .O(N__47730),
            .I(N__47721));
    LocalMux I__11085 (
            .O(N__47727),
            .I(N__47718));
    LocalMux I__11084 (
            .O(N__47724),
            .I(N__47715));
    LocalMux I__11083 (
            .O(N__47721),
            .I(data_cntvec_3));
    Odrv4 I__11082 (
            .O(N__47718),
            .I(data_cntvec_3));
    Odrv4 I__11081 (
            .O(N__47715),
            .I(data_cntvec_3));
    InMux I__11080 (
            .O(N__47708),
            .I(N__47705));
    LocalMux I__11079 (
            .O(N__47705),
            .I(N__47702));
    Span4Mux_h I__11078 (
            .O(N__47702),
            .I(N__47697));
    InMux I__11077 (
            .O(N__47701),
            .I(N__47692));
    InMux I__11076 (
            .O(N__47700),
            .I(N__47692));
    Odrv4 I__11075 (
            .O(N__47697),
            .I(req_data_cnt_3));
    LocalMux I__11074 (
            .O(N__47692),
            .I(req_data_cnt_3));
    InMux I__11073 (
            .O(N__47687),
            .I(N__47684));
    LocalMux I__11072 (
            .O(N__47684),
            .I(n20_adj_1596));
    CascadeMux I__11071 (
            .O(N__47681),
            .I(N__47677));
    CascadeMux I__11070 (
            .O(N__47680),
            .I(N__47674));
    InMux I__11069 (
            .O(N__47677),
            .I(N__47669));
    InMux I__11068 (
            .O(N__47674),
            .I(N__47666));
    CascadeMux I__11067 (
            .O(N__47673),
            .I(N__47663));
    InMux I__11066 (
            .O(N__47672),
            .I(N__47660));
    LocalMux I__11065 (
            .O(N__47669),
            .I(N__47657));
    LocalMux I__11064 (
            .O(N__47666),
            .I(N__47653));
    InMux I__11063 (
            .O(N__47663),
            .I(N__47650));
    LocalMux I__11062 (
            .O(N__47660),
            .I(N__47647));
    Span4Mux_v I__11061 (
            .O(N__47657),
            .I(N__47644));
    InMux I__11060 (
            .O(N__47656),
            .I(N__47641));
    Span4Mux_v I__11059 (
            .O(N__47653),
            .I(N__47634));
    LocalMux I__11058 (
            .O(N__47650),
            .I(N__47634));
    Span4Mux_h I__11057 (
            .O(N__47647),
            .I(N__47634));
    Span4Mux_v I__11056 (
            .O(N__47644),
            .I(N__47631));
    LocalMux I__11055 (
            .O(N__47641),
            .I(N__47627));
    Span4Mux_h I__11054 (
            .O(N__47634),
            .I(N__47624));
    Span4Mux_h I__11053 (
            .O(N__47631),
            .I(N__47621));
    InMux I__11052 (
            .O(N__47630),
            .I(N__47618));
    Span4Mux_v I__11051 (
            .O(N__47627),
            .I(N__47613));
    Span4Mux_v I__11050 (
            .O(N__47624),
            .I(N__47613));
    Odrv4 I__11049 (
            .O(N__47621),
            .I(comm_buf_1_7));
    LocalMux I__11048 (
            .O(N__47618),
            .I(comm_buf_1_7));
    Odrv4 I__11047 (
            .O(N__47613),
            .I(comm_buf_1_7));
    InMux I__11046 (
            .O(N__47606),
            .I(N__47603));
    LocalMux I__11045 (
            .O(N__47603),
            .I(N__47600));
    Span12Mux_v I__11044 (
            .O(N__47600),
            .I(N__47597));
    Odrv12 I__11043 (
            .O(N__47597),
            .I(n14_adj_1546));
    CascadeMux I__11042 (
            .O(N__47594),
            .I(n14_adj_1546_cascade_));
    CascadeMux I__11041 (
            .O(N__47591),
            .I(N__47588));
    InMux I__11040 (
            .O(N__47588),
            .I(N__47584));
    InMux I__11039 (
            .O(N__47587),
            .I(N__47581));
    LocalMux I__11038 (
            .O(N__47584),
            .I(N__47576));
    LocalMux I__11037 (
            .O(N__47581),
            .I(N__47576));
    Span4Mux_v I__11036 (
            .O(N__47576),
            .I(N__47572));
    InMux I__11035 (
            .O(N__47575),
            .I(N__47569));
    Span4Mux_h I__11034 (
            .O(N__47572),
            .I(N__47566));
    LocalMux I__11033 (
            .O(N__47569),
            .I(N__47563));
    Sp12to4 I__11032 (
            .O(N__47566),
            .I(N__47560));
    Odrv12 I__11031 (
            .O(N__47563),
            .I(n14_adj_1577));
    Odrv12 I__11030 (
            .O(N__47560),
            .I(n14_adj_1577));
    InMux I__11029 (
            .O(N__47555),
            .I(N__47552));
    LocalMux I__11028 (
            .O(N__47552),
            .I(N__47548));
    InMux I__11027 (
            .O(N__47551),
            .I(N__47544));
    Span12Mux_h I__11026 (
            .O(N__47548),
            .I(N__47541));
    InMux I__11025 (
            .O(N__47547),
            .I(N__47538));
    LocalMux I__11024 (
            .O(N__47544),
            .I(req_data_cnt_13));
    Odrv12 I__11023 (
            .O(N__47541),
            .I(req_data_cnt_13));
    LocalMux I__11022 (
            .O(N__47538),
            .I(req_data_cnt_13));
    InMux I__11021 (
            .O(N__47531),
            .I(N__47527));
    InMux I__11020 (
            .O(N__47530),
            .I(N__47523));
    LocalMux I__11019 (
            .O(N__47527),
            .I(N__47520));
    InMux I__11018 (
            .O(N__47526),
            .I(N__47517));
    LocalMux I__11017 (
            .O(N__47523),
            .I(data_cntvec_9));
    Odrv4 I__11016 (
            .O(N__47520),
            .I(data_cntvec_9));
    LocalMux I__11015 (
            .O(N__47517),
            .I(data_cntvec_9));
    InMux I__11014 (
            .O(N__47510),
            .I(N__47507));
    LocalMux I__11013 (
            .O(N__47507),
            .I(N__47503));
    InMux I__11012 (
            .O(N__47506),
            .I(N__47499));
    Span4Mux_h I__11011 (
            .O(N__47503),
            .I(N__47496));
    InMux I__11010 (
            .O(N__47502),
            .I(N__47493));
    LocalMux I__11009 (
            .O(N__47499),
            .I(req_data_cnt_15));
    Odrv4 I__11008 (
            .O(N__47496),
            .I(req_data_cnt_15));
    LocalMux I__11007 (
            .O(N__47493),
            .I(req_data_cnt_15));
    CascadeMux I__11006 (
            .O(N__47486),
            .I(N__47482));
    InMux I__11005 (
            .O(N__47485),
            .I(N__47479));
    InMux I__11004 (
            .O(N__47482),
            .I(N__47476));
    LocalMux I__11003 (
            .O(N__47479),
            .I(N__47471));
    LocalMux I__11002 (
            .O(N__47476),
            .I(N__47471));
    Odrv4 I__11001 (
            .O(N__47471),
            .I(data_cntvec_15));
    InMux I__11000 (
            .O(N__47468),
            .I(N__47465));
    LocalMux I__10999 (
            .O(N__47465),
            .I(n24));
    InMux I__10998 (
            .O(N__47462),
            .I(N__47458));
    InMux I__10997 (
            .O(N__47461),
            .I(N__47455));
    LocalMux I__10996 (
            .O(N__47458),
            .I(N__47452));
    LocalMux I__10995 (
            .O(N__47455),
            .I(N__47449));
    Span4Mux_v I__10994 (
            .O(N__47452),
            .I(N__47446));
    Sp12to4 I__10993 (
            .O(N__47449),
            .I(N__47443));
    Span4Mux_h I__10992 (
            .O(N__47446),
            .I(N__47440));
    Span12Mux_v I__10991 (
            .O(N__47443),
            .I(N__47437));
    Odrv4 I__10990 (
            .O(N__47440),
            .I(n14_adj_1574));
    Odrv12 I__10989 (
            .O(N__47437),
            .I(n14_adj_1574));
    InMux I__10988 (
            .O(N__47432),
            .I(N__47429));
    LocalMux I__10987 (
            .O(N__47429),
            .I(N__47424));
    InMux I__10986 (
            .O(N__47428),
            .I(N__47419));
    InMux I__10985 (
            .O(N__47427),
            .I(N__47419));
    Odrv4 I__10984 (
            .O(N__47424),
            .I(req_data_cnt_9));
    LocalMux I__10983 (
            .O(N__47419),
            .I(req_data_cnt_9));
    InMux I__10982 (
            .O(N__47414),
            .I(N__47406));
    InMux I__10981 (
            .O(N__47413),
            .I(N__47406));
    InMux I__10980 (
            .O(N__47412),
            .I(N__47401));
    InMux I__10979 (
            .O(N__47411),
            .I(N__47401));
    LocalMux I__10978 (
            .O(N__47406),
            .I(N__47398));
    LocalMux I__10977 (
            .O(N__47401),
            .I(N__47392));
    Span4Mux_h I__10976 (
            .O(N__47398),
            .I(N__47389));
    InMux I__10975 (
            .O(N__47397),
            .I(N__47382));
    InMux I__10974 (
            .O(N__47396),
            .I(N__47382));
    InMux I__10973 (
            .O(N__47395),
            .I(N__47382));
    Span4Mux_v I__10972 (
            .O(N__47392),
            .I(N__47372));
    Span4Mux_h I__10971 (
            .O(N__47389),
            .I(N__47367));
    LocalMux I__10970 (
            .O(N__47382),
            .I(N__47367));
    InMux I__10969 (
            .O(N__47381),
            .I(N__47358));
    InMux I__10968 (
            .O(N__47380),
            .I(N__47358));
    InMux I__10967 (
            .O(N__47379),
            .I(N__47358));
    InMux I__10966 (
            .O(N__47378),
            .I(N__47358));
    InMux I__10965 (
            .O(N__47377),
            .I(N__47351));
    InMux I__10964 (
            .O(N__47376),
            .I(N__47351));
    InMux I__10963 (
            .O(N__47375),
            .I(N__47351));
    Span4Mux_h I__10962 (
            .O(N__47372),
            .I(N__47347));
    Span4Mux_v I__10961 (
            .O(N__47367),
            .I(N__47344));
    LocalMux I__10960 (
            .O(N__47358),
            .I(N__47339));
    LocalMux I__10959 (
            .O(N__47351),
            .I(N__47339));
    InMux I__10958 (
            .O(N__47350),
            .I(N__47336));
    Odrv4 I__10957 (
            .O(N__47347),
            .I(n12467));
    Odrv4 I__10956 (
            .O(N__47344),
            .I(n12467));
    Odrv12 I__10955 (
            .O(N__47339),
            .I(n12467));
    LocalMux I__10954 (
            .O(N__47336),
            .I(n12467));
    CascadeMux I__10953 (
            .O(N__47327),
            .I(N__47323));
    InMux I__10952 (
            .O(N__47326),
            .I(N__47319));
    InMux I__10951 (
            .O(N__47323),
            .I(N__47316));
    InMux I__10950 (
            .O(N__47322),
            .I(N__47313));
    LocalMux I__10949 (
            .O(N__47319),
            .I(N__47310));
    LocalMux I__10948 (
            .O(N__47316),
            .I(N__47307));
    LocalMux I__10947 (
            .O(N__47313),
            .I(N__47304));
    Span4Mux_v I__10946 (
            .O(N__47310),
            .I(N__47301));
    Span12Mux_v I__10945 (
            .O(N__47307),
            .I(N__47296));
    Span12Mux_h I__10944 (
            .O(N__47304),
            .I(N__47296));
    Odrv4 I__10943 (
            .O(N__47301),
            .I(n14_adj_1578));
    Odrv12 I__10942 (
            .O(N__47296),
            .I(n14_adj_1578));
    CascadeMux I__10941 (
            .O(N__47291),
            .I(N__47288));
    InMux I__10940 (
            .O(N__47288),
            .I(N__47285));
    LocalMux I__10939 (
            .O(N__47285),
            .I(N__47280));
    CascadeMux I__10938 (
            .O(N__47284),
            .I(N__47277));
    InMux I__10937 (
            .O(N__47283),
            .I(N__47274));
    Span4Mux_v I__10936 (
            .O(N__47280),
            .I(N__47271));
    InMux I__10935 (
            .O(N__47277),
            .I(N__47268));
    LocalMux I__10934 (
            .O(N__47274),
            .I(N__47263));
    Span4Mux_v I__10933 (
            .O(N__47271),
            .I(N__47263));
    LocalMux I__10932 (
            .O(N__47268),
            .I(N__47260));
    Odrv4 I__10931 (
            .O(N__47263),
            .I(req_data_cnt_5));
    Odrv4 I__10930 (
            .O(N__47260),
            .I(req_data_cnt_5));
    CascadeMux I__10929 (
            .O(N__47255),
            .I(n22211_cascade_));
    CascadeMux I__10928 (
            .O(N__47252),
            .I(N__47249));
    InMux I__10927 (
            .O(N__47249),
            .I(N__47243));
    CascadeMux I__10926 (
            .O(N__47248),
            .I(N__47238));
    InMux I__10925 (
            .O(N__47247),
            .I(N__47235));
    InMux I__10924 (
            .O(N__47246),
            .I(N__47231));
    LocalMux I__10923 (
            .O(N__47243),
            .I(N__47228));
    InMux I__10922 (
            .O(N__47242),
            .I(N__47225));
    InMux I__10921 (
            .O(N__47241),
            .I(N__47222));
    InMux I__10920 (
            .O(N__47238),
            .I(N__47218));
    LocalMux I__10919 (
            .O(N__47235),
            .I(N__47215));
    InMux I__10918 (
            .O(N__47234),
            .I(N__47212));
    LocalMux I__10917 (
            .O(N__47231),
            .I(N__47209));
    Span4Mux_v I__10916 (
            .O(N__47228),
            .I(N__47202));
    LocalMux I__10915 (
            .O(N__47225),
            .I(N__47202));
    LocalMux I__10914 (
            .O(N__47222),
            .I(N__47202));
    InMux I__10913 (
            .O(N__47221),
            .I(N__47199));
    LocalMux I__10912 (
            .O(N__47218),
            .I(N__47196));
    Sp12to4 I__10911 (
            .O(N__47215),
            .I(N__47191));
    LocalMux I__10910 (
            .O(N__47212),
            .I(N__47191));
    Span4Mux_v I__10909 (
            .O(N__47209),
            .I(N__47188));
    Span4Mux_v I__10908 (
            .O(N__47202),
            .I(N__47185));
    LocalMux I__10907 (
            .O(N__47199),
            .I(N__47182));
    Span12Mux_h I__10906 (
            .O(N__47196),
            .I(N__47178));
    Span12Mux_v I__10905 (
            .O(N__47191),
            .I(N__47175));
    Span4Mux_v I__10904 (
            .O(N__47188),
            .I(N__47170));
    Span4Mux_v I__10903 (
            .O(N__47185),
            .I(N__47170));
    Span4Mux_h I__10902 (
            .O(N__47182),
            .I(N__47167));
    InMux I__10901 (
            .O(N__47181),
            .I(N__47164));
    Odrv12 I__10900 (
            .O(N__47178),
            .I(comm_rx_buf_2));
    Odrv12 I__10899 (
            .O(N__47175),
            .I(comm_rx_buf_2));
    Odrv4 I__10898 (
            .O(N__47170),
            .I(comm_rx_buf_2));
    Odrv4 I__10897 (
            .O(N__47167),
            .I(comm_rx_buf_2));
    LocalMux I__10896 (
            .O(N__47164),
            .I(comm_rx_buf_2));
    CascadeMux I__10895 (
            .O(N__47153),
            .I(n30_adj_1518_cascade_));
    CascadeMux I__10894 (
            .O(N__47150),
            .I(N__47147));
    InMux I__10893 (
            .O(N__47147),
            .I(N__47144));
    LocalMux I__10892 (
            .O(N__47144),
            .I(N__47140));
    CascadeMux I__10891 (
            .O(N__47143),
            .I(N__47136));
    Span4Mux_v I__10890 (
            .O(N__47140),
            .I(N__47130));
    InMux I__10889 (
            .O(N__47139),
            .I(N__47127));
    InMux I__10888 (
            .O(N__47136),
            .I(N__47124));
    InMux I__10887 (
            .O(N__47135),
            .I(N__47121));
    InMux I__10886 (
            .O(N__47134),
            .I(N__47118));
    InMux I__10885 (
            .O(N__47133),
            .I(N__47115));
    Span4Mux_h I__10884 (
            .O(N__47130),
            .I(N__47110));
    LocalMux I__10883 (
            .O(N__47127),
            .I(N__47110));
    LocalMux I__10882 (
            .O(N__47124),
            .I(N__47105));
    LocalMux I__10881 (
            .O(N__47121),
            .I(N__47105));
    LocalMux I__10880 (
            .O(N__47118),
            .I(N__47102));
    LocalMux I__10879 (
            .O(N__47115),
            .I(N__47099));
    Span4Mux_v I__10878 (
            .O(N__47110),
            .I(N__47096));
    Span12Mux_h I__10877 (
            .O(N__47105),
            .I(N__47093));
    Span4Mux_h I__10876 (
            .O(N__47102),
            .I(N__47090));
    Span4Mux_v I__10875 (
            .O(N__47099),
            .I(N__47087));
    Span4Mux_h I__10874 (
            .O(N__47096),
            .I(N__47084));
    Odrv12 I__10873 (
            .O(N__47093),
            .I(comm_buf_1_2));
    Odrv4 I__10872 (
            .O(N__47090),
            .I(comm_buf_1_2));
    Odrv4 I__10871 (
            .O(N__47087),
            .I(comm_buf_1_2));
    Odrv4 I__10870 (
            .O(N__47084),
            .I(comm_buf_1_2));
    CEMux I__10869 (
            .O(N__47075),
            .I(N__47072));
    LocalMux I__10868 (
            .O(N__47072),
            .I(N__47065));
    CEMux I__10867 (
            .O(N__47071),
            .I(N__47062));
    CEMux I__10866 (
            .O(N__47070),
            .I(N__47058));
    CEMux I__10865 (
            .O(N__47069),
            .I(N__47055));
    CEMux I__10864 (
            .O(N__47068),
            .I(N__47050));
    Span4Mux_h I__10863 (
            .O(N__47065),
            .I(N__47045));
    LocalMux I__10862 (
            .O(N__47062),
            .I(N__47045));
    CEMux I__10861 (
            .O(N__47061),
            .I(N__47042));
    LocalMux I__10860 (
            .O(N__47058),
            .I(N__47039));
    LocalMux I__10859 (
            .O(N__47055),
            .I(N__47036));
    CEMux I__10858 (
            .O(N__47054),
            .I(N__47033));
    CEMux I__10857 (
            .O(N__47053),
            .I(N__47030));
    LocalMux I__10856 (
            .O(N__47050),
            .I(N__47022));
    Span4Mux_h I__10855 (
            .O(N__47045),
            .I(N__47022));
    LocalMux I__10854 (
            .O(N__47042),
            .I(N__47022));
    Span4Mux_h I__10853 (
            .O(N__47039),
            .I(N__47015));
    Span4Mux_h I__10852 (
            .O(N__47036),
            .I(N__47015));
    LocalMux I__10851 (
            .O(N__47033),
            .I(N__47015));
    LocalMux I__10850 (
            .O(N__47030),
            .I(N__47012));
    InMux I__10849 (
            .O(N__47029),
            .I(N__47009));
    Odrv4 I__10848 (
            .O(N__47022),
            .I(n12047));
    Odrv4 I__10847 (
            .O(N__47015),
            .I(n12047));
    Odrv12 I__10846 (
            .O(N__47012),
            .I(n12047));
    LocalMux I__10845 (
            .O(N__47009),
            .I(n12047));
    SRMux I__10844 (
            .O(N__47000),
            .I(N__46997));
    LocalMux I__10843 (
            .O(N__46997),
            .I(N__46990));
    SRMux I__10842 (
            .O(N__46996),
            .I(N__46986));
    SRMux I__10841 (
            .O(N__46995),
            .I(N__46983));
    SRMux I__10840 (
            .O(N__46994),
            .I(N__46980));
    SRMux I__10839 (
            .O(N__46993),
            .I(N__46977));
    Span4Mux_v I__10838 (
            .O(N__46990),
            .I(N__46974));
    SRMux I__10837 (
            .O(N__46989),
            .I(N__46971));
    LocalMux I__10836 (
            .O(N__46986),
            .I(N__46966));
    LocalMux I__10835 (
            .O(N__46983),
            .I(N__46963));
    LocalMux I__10834 (
            .O(N__46980),
            .I(N__46960));
    LocalMux I__10833 (
            .O(N__46977),
            .I(N__46957));
    Span4Mux_h I__10832 (
            .O(N__46974),
            .I(N__46952));
    LocalMux I__10831 (
            .O(N__46971),
            .I(N__46952));
    SRMux I__10830 (
            .O(N__46970),
            .I(N__46949));
    SRMux I__10829 (
            .O(N__46969),
            .I(N__46946));
    Span4Mux_v I__10828 (
            .O(N__46966),
            .I(N__46941));
    Span4Mux_v I__10827 (
            .O(N__46963),
            .I(N__46941));
    Span4Mux_v I__10826 (
            .O(N__46960),
            .I(N__46936));
    Span4Mux_h I__10825 (
            .O(N__46957),
            .I(N__46936));
    Span4Mux_h I__10824 (
            .O(N__46952),
            .I(N__46933));
    LocalMux I__10823 (
            .O(N__46949),
            .I(N__46930));
    LocalMux I__10822 (
            .O(N__46946),
            .I(N__46927));
    Odrv4 I__10821 (
            .O(N__46941),
            .I(n14773));
    Odrv4 I__10820 (
            .O(N__46936),
            .I(n14773));
    Odrv4 I__10819 (
            .O(N__46933),
            .I(n14773));
    Odrv12 I__10818 (
            .O(N__46930),
            .I(n14773));
    Odrv12 I__10817 (
            .O(N__46927),
            .I(n14773));
    InMux I__10816 (
            .O(N__46916),
            .I(N__46913));
    LocalMux I__10815 (
            .O(N__46913),
            .I(N__46910));
    Span4Mux_h I__10814 (
            .O(N__46910),
            .I(N__46907));
    Span4Mux_h I__10813 (
            .O(N__46907),
            .I(N__46904));
    Odrv4 I__10812 (
            .O(N__46904),
            .I(n19_adj_1516));
    CascadeMux I__10811 (
            .O(N__46901),
            .I(N__46898));
    InMux I__10810 (
            .O(N__46898),
            .I(N__46895));
    LocalMux I__10809 (
            .O(N__46895),
            .I(N__46892));
    Span12Mux_h I__10808 (
            .O(N__46892),
            .I(N__46888));
    InMux I__10807 (
            .O(N__46891),
            .I(N__46885));
    Odrv12 I__10806 (
            .O(N__46888),
            .I(buf_readRTD_2));
    LocalMux I__10805 (
            .O(N__46885),
            .I(buf_readRTD_2));
    InMux I__10804 (
            .O(N__46880),
            .I(N__46877));
    LocalMux I__10803 (
            .O(N__46877),
            .I(n21956));
    InMux I__10802 (
            .O(N__46874),
            .I(N__46871));
    LocalMux I__10801 (
            .O(N__46871),
            .I(N__46867));
    CascadeMux I__10800 (
            .O(N__46870),
            .I(N__46864));
    Span4Mux_h I__10799 (
            .O(N__46867),
            .I(N__46861));
    InMux I__10798 (
            .O(N__46864),
            .I(N__46858));
    Span4Mux_h I__10797 (
            .O(N__46861),
            .I(N__46855));
    LocalMux I__10796 (
            .O(N__46858),
            .I(data_idxvec_2));
    Odrv4 I__10795 (
            .O(N__46855),
            .I(data_idxvec_2));
    InMux I__10794 (
            .O(N__46850),
            .I(N__46846));
    InMux I__10793 (
            .O(N__46849),
            .I(N__46842));
    LocalMux I__10792 (
            .O(N__46846),
            .I(N__46839));
    InMux I__10791 (
            .O(N__46845),
            .I(N__46836));
    LocalMux I__10790 (
            .O(N__46842),
            .I(N__46833));
    Span4Mux_h I__10789 (
            .O(N__46839),
            .I(N__46830));
    LocalMux I__10788 (
            .O(N__46836),
            .I(data_cntvec_2));
    Odrv4 I__10787 (
            .O(N__46833),
            .I(data_cntvec_2));
    Odrv4 I__10786 (
            .O(N__46830),
            .I(data_cntvec_2));
    InMux I__10785 (
            .O(N__46823),
            .I(N__46820));
    LocalMux I__10784 (
            .O(N__46820),
            .I(n26_adj_1517));
    InMux I__10783 (
            .O(N__46817),
            .I(N__46813));
    InMux I__10782 (
            .O(N__46816),
            .I(N__46810));
    LocalMux I__10781 (
            .O(N__46813),
            .I(N__46807));
    LocalMux I__10780 (
            .O(N__46810),
            .I(N__46804));
    Span4Mux_h I__10779 (
            .O(N__46807),
            .I(N__46799));
    Span4Mux_v I__10778 (
            .O(N__46804),
            .I(N__46799));
    Odrv4 I__10777 (
            .O(N__46799),
            .I(n14_adj_1550));
    InMux I__10776 (
            .O(N__46796),
            .I(N__46792));
    InMux I__10775 (
            .O(N__46795),
            .I(N__46789));
    LocalMux I__10774 (
            .O(N__46792),
            .I(N__46786));
    LocalMux I__10773 (
            .O(N__46789),
            .I(N__46783));
    Span4Mux_h I__10772 (
            .O(N__46786),
            .I(N__46780));
    Span4Mux_h I__10771 (
            .O(N__46783),
            .I(N__46777));
    Odrv4 I__10770 (
            .O(N__46780),
            .I(n14_adj_1544));
    Odrv4 I__10769 (
            .O(N__46777),
            .I(n14_adj_1544));
    InMux I__10768 (
            .O(N__46772),
            .I(N__46769));
    LocalMux I__10767 (
            .O(N__46769),
            .I(N__46764));
    InMux I__10766 (
            .O(N__46768),
            .I(N__46761));
    InMux I__10765 (
            .O(N__46767),
            .I(N__46758));
    Span4Mux_h I__10764 (
            .O(N__46764),
            .I(N__46755));
    LocalMux I__10763 (
            .O(N__46761),
            .I(N__46752));
    LocalMux I__10762 (
            .O(N__46758),
            .I(data_cntvec_1));
    Odrv4 I__10761 (
            .O(N__46755),
            .I(data_cntvec_1));
    Odrv4 I__10760 (
            .O(N__46752),
            .I(data_cntvec_1));
    InMux I__10759 (
            .O(N__46745),
            .I(N__46741));
    InMux I__10758 (
            .O(N__46744),
            .I(N__46737));
    LocalMux I__10757 (
            .O(N__46741),
            .I(N__46734));
    InMux I__10756 (
            .O(N__46740),
            .I(N__46731));
    LocalMux I__10755 (
            .O(N__46737),
            .I(data_cntvec_4));
    Odrv4 I__10754 (
            .O(N__46734),
            .I(data_cntvec_4));
    LocalMux I__10753 (
            .O(N__46731),
            .I(data_cntvec_4));
    InMux I__10752 (
            .O(N__46724),
            .I(N__46720));
    CascadeMux I__10751 (
            .O(N__46723),
            .I(N__46717));
    LocalMux I__10750 (
            .O(N__46720),
            .I(N__46713));
    InMux I__10749 (
            .O(N__46717),
            .I(N__46710));
    InMux I__10748 (
            .O(N__46716),
            .I(N__46707));
    Span4Mux_h I__10747 (
            .O(N__46713),
            .I(N__46704));
    LocalMux I__10746 (
            .O(N__46710),
            .I(N__46701));
    LocalMux I__10745 (
            .O(N__46707),
            .I(req_data_cnt_4));
    Odrv4 I__10744 (
            .O(N__46704),
            .I(req_data_cnt_4));
    Odrv4 I__10743 (
            .O(N__46701),
            .I(req_data_cnt_4));
    InMux I__10742 (
            .O(N__46694),
            .I(N__46691));
    LocalMux I__10741 (
            .O(N__46691),
            .I(N__46686));
    InMux I__10740 (
            .O(N__46690),
            .I(N__46681));
    InMux I__10739 (
            .O(N__46689),
            .I(N__46681));
    Odrv4 I__10738 (
            .O(N__46686),
            .I(req_data_cnt_1));
    LocalMux I__10737 (
            .O(N__46681),
            .I(req_data_cnt_1));
    InMux I__10736 (
            .O(N__46676),
            .I(N__46673));
    LocalMux I__10735 (
            .O(N__46673),
            .I(n18));
    InMux I__10734 (
            .O(N__46670),
            .I(N__46667));
    LocalMux I__10733 (
            .O(N__46667),
            .I(N__46663));
    CascadeMux I__10732 (
            .O(N__46666),
            .I(N__46660));
    Span12Mux_v I__10731 (
            .O(N__46663),
            .I(N__46657));
    InMux I__10730 (
            .O(N__46660),
            .I(N__46654));
    Odrv12 I__10729 (
            .O(N__46657),
            .I(buf_adcdata_vdc_13));
    LocalMux I__10728 (
            .O(N__46654),
            .I(buf_adcdata_vdc_13));
    InMux I__10727 (
            .O(N__46649),
            .I(N__46646));
    LocalMux I__10726 (
            .O(N__46646),
            .I(N__46643));
    Span4Mux_v I__10725 (
            .O(N__46643),
            .I(N__46639));
    InMux I__10724 (
            .O(N__46642),
            .I(N__46636));
    Span4Mux_h I__10723 (
            .O(N__46639),
            .I(N__46630));
    LocalMux I__10722 (
            .O(N__46636),
            .I(N__46630));
    InMux I__10721 (
            .O(N__46635),
            .I(N__46627));
    Span4Mux_h I__10720 (
            .O(N__46630),
            .I(N__46624));
    LocalMux I__10719 (
            .O(N__46627),
            .I(buf_adcdata_vac_13));
    Odrv4 I__10718 (
            .O(N__46624),
            .I(buf_adcdata_vac_13));
    InMux I__10717 (
            .O(N__46619),
            .I(N__46616));
    LocalMux I__10716 (
            .O(N__46616),
            .I(n19_adj_1497));
    InMux I__10715 (
            .O(N__46613),
            .I(N__46610));
    LocalMux I__10714 (
            .O(N__46610),
            .I(N__46606));
    InMux I__10713 (
            .O(N__46609),
            .I(N__46603));
    Span4Mux_v I__10712 (
            .O(N__46606),
            .I(N__46600));
    LocalMux I__10711 (
            .O(N__46603),
            .I(N__46597));
    Sp12to4 I__10710 (
            .O(N__46600),
            .I(N__46594));
    Span4Mux_h I__10709 (
            .O(N__46597),
            .I(N__46591));
    Odrv12 I__10708 (
            .O(N__46594),
            .I(n9));
    Odrv4 I__10707 (
            .O(N__46591),
            .I(n9));
    InMux I__10706 (
            .O(N__46586),
            .I(N__46582));
    InMux I__10705 (
            .O(N__46585),
            .I(N__46578));
    LocalMux I__10704 (
            .O(N__46582),
            .I(N__46575));
    InMux I__10703 (
            .O(N__46581),
            .I(N__46572));
    LocalMux I__10702 (
            .O(N__46578),
            .I(N__46566));
    Span4Mux_v I__10701 (
            .O(N__46575),
            .I(N__46566));
    LocalMux I__10700 (
            .O(N__46572),
            .I(N__46563));
    InMux I__10699 (
            .O(N__46571),
            .I(N__46560));
    Span4Mux_h I__10698 (
            .O(N__46566),
            .I(N__46555));
    Span4Mux_v I__10697 (
            .O(N__46563),
            .I(N__46555));
    LocalMux I__10696 (
            .O(N__46560),
            .I(n20663));
    Odrv4 I__10695 (
            .O(N__46555),
            .I(n20663));
    CascadeMux I__10694 (
            .O(N__46550),
            .I(n12467_cascade_));
    InMux I__10693 (
            .O(N__46547),
            .I(N__46544));
    LocalMux I__10692 (
            .O(N__46544),
            .I(N__46540));
    InMux I__10691 (
            .O(N__46543),
            .I(N__46537));
    Span4Mux_h I__10690 (
            .O(N__46540),
            .I(N__46532));
    LocalMux I__10689 (
            .O(N__46537),
            .I(N__46532));
    Span4Mux_h I__10688 (
            .O(N__46532),
            .I(N__46529));
    Span4Mux_h I__10687 (
            .O(N__46529),
            .I(N__46526));
    Odrv4 I__10686 (
            .O(N__46526),
            .I(n14_adj_1533));
    InMux I__10685 (
            .O(N__46523),
            .I(N__46518));
    InMux I__10684 (
            .O(N__46522),
            .I(N__46515));
    InMux I__10683 (
            .O(N__46521),
            .I(N__46512));
    LocalMux I__10682 (
            .O(N__46518),
            .I(N__46509));
    LocalMux I__10681 (
            .O(N__46515),
            .I(N__46506));
    LocalMux I__10680 (
            .O(N__46512),
            .I(N__46499));
    Span4Mux_v I__10679 (
            .O(N__46509),
            .I(N__46499));
    Span4Mux_v I__10678 (
            .O(N__46506),
            .I(N__46499));
    Odrv4 I__10677 (
            .O(N__46499),
            .I(data_cntvec_6));
    InMux I__10676 (
            .O(N__46496),
            .I(N__46493));
    LocalMux I__10675 (
            .O(N__46493),
            .I(N__46488));
    InMux I__10674 (
            .O(N__46492),
            .I(N__46485));
    InMux I__10673 (
            .O(N__46491),
            .I(N__46482));
    Span4Mux_h I__10672 (
            .O(N__46488),
            .I(N__46479));
    LocalMux I__10671 (
            .O(N__46485),
            .I(N__46476));
    LocalMux I__10670 (
            .O(N__46482),
            .I(data_cntvec_0));
    Odrv4 I__10669 (
            .O(N__46479),
            .I(data_cntvec_0));
    Odrv4 I__10668 (
            .O(N__46476),
            .I(data_cntvec_0));
    CascadeMux I__10667 (
            .O(N__46469),
            .I(N__46466));
    InMux I__10666 (
            .O(N__46466),
            .I(N__46462));
    CascadeMux I__10665 (
            .O(N__46465),
            .I(N__46458));
    LocalMux I__10664 (
            .O(N__46462),
            .I(N__46455));
    InMux I__10663 (
            .O(N__46461),
            .I(N__46450));
    InMux I__10662 (
            .O(N__46458),
            .I(N__46450));
    Odrv4 I__10661 (
            .O(N__46455),
            .I(req_data_cnt_0));
    LocalMux I__10660 (
            .O(N__46450),
            .I(req_data_cnt_0));
    InMux I__10659 (
            .O(N__46445),
            .I(N__46442));
    LocalMux I__10658 (
            .O(N__46442),
            .I(N__46439));
    Odrv4 I__10657 (
            .O(N__46439),
            .I(n17));
    InMux I__10656 (
            .O(N__46436),
            .I(N__46433));
    LocalMux I__10655 (
            .O(N__46433),
            .I(N__46430));
    Span4Mux_h I__10654 (
            .O(N__46430),
            .I(N__46427));
    Span4Mux_h I__10653 (
            .O(N__46427),
            .I(N__46424));
    Odrv4 I__10652 (
            .O(N__46424),
            .I(n16_adj_1515));
    CascadeMux I__10651 (
            .O(N__46421),
            .I(N__46417));
    CascadeMux I__10650 (
            .O(N__46420),
            .I(N__46414));
    InMux I__10649 (
            .O(N__46417),
            .I(N__46411));
    InMux I__10648 (
            .O(N__46414),
            .I(N__46407));
    LocalMux I__10647 (
            .O(N__46411),
            .I(N__46402));
    CascadeMux I__10646 (
            .O(N__46410),
            .I(N__46399));
    LocalMux I__10645 (
            .O(N__46407),
            .I(N__46396));
    InMux I__10644 (
            .O(N__46406),
            .I(N__46393));
    InMux I__10643 (
            .O(N__46405),
            .I(N__46390));
    Span4Mux_h I__10642 (
            .O(N__46402),
            .I(N__46387));
    InMux I__10641 (
            .O(N__46399),
            .I(N__46384));
    Span4Mux_v I__10640 (
            .O(N__46396),
            .I(N__46379));
    LocalMux I__10639 (
            .O(N__46393),
            .I(N__46379));
    LocalMux I__10638 (
            .O(N__46390),
            .I(N__46376));
    Span4Mux_h I__10637 (
            .O(N__46387),
            .I(N__46371));
    LocalMux I__10636 (
            .O(N__46384),
            .I(N__46371));
    Span4Mux_v I__10635 (
            .O(N__46379),
            .I(N__46368));
    Span4Mux_v I__10634 (
            .O(N__46376),
            .I(N__46362));
    Span4Mux_v I__10633 (
            .O(N__46371),
            .I(N__46362));
    Span4Mux_h I__10632 (
            .O(N__46368),
            .I(N__46359));
    InMux I__10631 (
            .O(N__46367),
            .I(N__46356));
    Span4Mux_h I__10630 (
            .O(N__46362),
            .I(N__46352));
    Span4Mux_h I__10629 (
            .O(N__46359),
            .I(N__46347));
    LocalMux I__10628 (
            .O(N__46356),
            .I(N__46347));
    InMux I__10627 (
            .O(N__46355),
            .I(N__46344));
    Span4Mux_v I__10626 (
            .O(N__46352),
            .I(N__46341));
    Span4Mux_v I__10625 (
            .O(N__46347),
            .I(N__46336));
    LocalMux I__10624 (
            .O(N__46344),
            .I(N__46336));
    Odrv4 I__10623 (
            .O(N__46341),
            .I(comm_buf_0_5));
    Odrv4 I__10622 (
            .O(N__46336),
            .I(comm_buf_0_5));
    InMux I__10621 (
            .O(N__46331),
            .I(N__46328));
    LocalMux I__10620 (
            .O(N__46328),
            .I(N__46325));
    Span4Mux_h I__10619 (
            .O(N__46325),
            .I(N__46320));
    InMux I__10618 (
            .O(N__46324),
            .I(N__46315));
    InMux I__10617 (
            .O(N__46323),
            .I(N__46315));
    Odrv4 I__10616 (
            .O(N__46320),
            .I(req_data_cnt_6));
    LocalMux I__10615 (
            .O(N__46315),
            .I(req_data_cnt_6));
    InMux I__10614 (
            .O(N__46310),
            .I(N__46305));
    InMux I__10613 (
            .O(N__46309),
            .I(N__46302));
    InMux I__10612 (
            .O(N__46308),
            .I(N__46299));
    LocalMux I__10611 (
            .O(N__46305),
            .I(req_data_cnt_2));
    LocalMux I__10610 (
            .O(N__46302),
            .I(req_data_cnt_2));
    LocalMux I__10609 (
            .O(N__46299),
            .I(req_data_cnt_2));
    CascadeMux I__10608 (
            .O(N__46292),
            .I(n22208_cascade_));
    InMux I__10607 (
            .O(N__46289),
            .I(N__46285));
    CascadeMux I__10606 (
            .O(N__46288),
            .I(N__46282));
    LocalMux I__10605 (
            .O(N__46285),
            .I(N__46279));
    InMux I__10604 (
            .O(N__46282),
            .I(N__46275));
    Span4Mux_v I__10603 (
            .O(N__46279),
            .I(N__46272));
    InMux I__10602 (
            .O(N__46278),
            .I(N__46269));
    LocalMux I__10601 (
            .O(N__46275),
            .I(acadc_skipCount_2));
    Odrv4 I__10600 (
            .O(N__46272),
            .I(acadc_skipCount_2));
    LocalMux I__10599 (
            .O(N__46269),
            .I(acadc_skipCount_2));
    InMux I__10598 (
            .O(N__46262),
            .I(N__46259));
    LocalMux I__10597 (
            .O(N__46259),
            .I(N__46256));
    Odrv4 I__10596 (
            .O(N__46256),
            .I(n21959));
    InMux I__10595 (
            .O(N__46253),
            .I(N__46250));
    LocalMux I__10594 (
            .O(N__46250),
            .I(N__46247));
    Span4Mux_v I__10593 (
            .O(N__46247),
            .I(N__46244));
    Odrv4 I__10592 (
            .O(N__46244),
            .I(comm_buf_3_7));
    InMux I__10591 (
            .O(N__46241),
            .I(N__46238));
    LocalMux I__10590 (
            .O(N__46238),
            .I(N__46235));
    Span4Mux_v I__10589 (
            .O(N__46235),
            .I(N__46232));
    Span4Mux_h I__10588 (
            .O(N__46232),
            .I(N__46229));
    Odrv4 I__10587 (
            .O(N__46229),
            .I(comm_buf_2_7));
    CascadeMux I__10586 (
            .O(N__46226),
            .I(n2_adj_1581_cascade_));
    CEMux I__10585 (
            .O(N__46223),
            .I(N__46220));
    LocalMux I__10584 (
            .O(N__46220),
            .I(N__46215));
    InMux I__10583 (
            .O(N__46219),
            .I(N__46209));
    CEMux I__10582 (
            .O(N__46218),
            .I(N__46206));
    Span4Mux_v I__10581 (
            .O(N__46215),
            .I(N__46202));
    CEMux I__10580 (
            .O(N__46214),
            .I(N__46199));
    CEMux I__10579 (
            .O(N__46213),
            .I(N__46195));
    CEMux I__10578 (
            .O(N__46212),
            .I(N__46192));
    LocalMux I__10577 (
            .O(N__46209),
            .I(N__46189));
    LocalMux I__10576 (
            .O(N__46206),
            .I(N__46186));
    CEMux I__10575 (
            .O(N__46205),
            .I(N__46183));
    Span4Mux_h I__10574 (
            .O(N__46202),
            .I(N__46178));
    LocalMux I__10573 (
            .O(N__46199),
            .I(N__46178));
    CEMux I__10572 (
            .O(N__46198),
            .I(N__46175));
    LocalMux I__10571 (
            .O(N__46195),
            .I(N__46172));
    LocalMux I__10570 (
            .O(N__46192),
            .I(N__46169));
    Span4Mux_h I__10569 (
            .O(N__46189),
            .I(N__46166));
    Span4Mux_h I__10568 (
            .O(N__46186),
            .I(N__46161));
    LocalMux I__10567 (
            .O(N__46183),
            .I(N__46161));
    Span4Mux_v I__10566 (
            .O(N__46178),
            .I(N__46156));
    LocalMux I__10565 (
            .O(N__46175),
            .I(N__46156));
    Span4Mux_v I__10564 (
            .O(N__46172),
            .I(N__46149));
    Span4Mux_h I__10563 (
            .O(N__46169),
            .I(N__46149));
    Span4Mux_v I__10562 (
            .O(N__46166),
            .I(N__46149));
    Odrv4 I__10561 (
            .O(N__46161),
            .I(n11503));
    Odrv4 I__10560 (
            .O(N__46156),
            .I(n11503));
    Odrv4 I__10559 (
            .O(N__46149),
            .I(n11503));
    SRMux I__10558 (
            .O(N__46142),
            .I(N__46137));
    SRMux I__10557 (
            .O(N__46141),
            .I(N__46134));
    SRMux I__10556 (
            .O(N__46140),
            .I(N__46129));
    LocalMux I__10555 (
            .O(N__46137),
            .I(N__46126));
    LocalMux I__10554 (
            .O(N__46134),
            .I(N__46123));
    SRMux I__10553 (
            .O(N__46133),
            .I(N__46120));
    SRMux I__10552 (
            .O(N__46132),
            .I(N__46117));
    LocalMux I__10551 (
            .O(N__46129),
            .I(N__46112));
    Span4Mux_v I__10550 (
            .O(N__46126),
            .I(N__46103));
    Span4Mux_h I__10549 (
            .O(N__46123),
            .I(N__46103));
    LocalMux I__10548 (
            .O(N__46120),
            .I(N__46103));
    LocalMux I__10547 (
            .O(N__46117),
            .I(N__46103));
    SRMux I__10546 (
            .O(N__46116),
            .I(N__46100));
    SRMux I__10545 (
            .O(N__46115),
            .I(N__46097));
    Span4Mux_v I__10544 (
            .O(N__46112),
            .I(N__46094));
    Span4Mux_v I__10543 (
            .O(N__46103),
            .I(N__46091));
    LocalMux I__10542 (
            .O(N__46100),
            .I(N__46088));
    LocalMux I__10541 (
            .O(N__46097),
            .I(N__46085));
    Span4Mux_h I__10540 (
            .O(N__46094),
            .I(N__46080));
    Span4Mux_h I__10539 (
            .O(N__46091),
            .I(N__46080));
    Span4Mux_h I__10538 (
            .O(N__46088),
            .I(N__46077));
    Span4Mux_v I__10537 (
            .O(N__46085),
            .I(N__46074));
    Odrv4 I__10536 (
            .O(N__46080),
            .I(n14815));
    Odrv4 I__10535 (
            .O(N__46077),
            .I(n14815));
    Odrv4 I__10534 (
            .O(N__46074),
            .I(n14815));
    CascadeMux I__10533 (
            .O(N__46067),
            .I(N__46063));
    CascadeMux I__10532 (
            .O(N__46066),
            .I(N__46060));
    InMux I__10531 (
            .O(N__46063),
            .I(N__46055));
    InMux I__10530 (
            .O(N__46060),
            .I(N__46052));
    InMux I__10529 (
            .O(N__46059),
            .I(N__46049));
    CascadeMux I__10528 (
            .O(N__46058),
            .I(N__46045));
    LocalMux I__10527 (
            .O(N__46055),
            .I(N__46042));
    LocalMux I__10526 (
            .O(N__46052),
            .I(N__46038));
    LocalMux I__10525 (
            .O(N__46049),
            .I(N__46035));
    InMux I__10524 (
            .O(N__46048),
            .I(N__46032));
    InMux I__10523 (
            .O(N__46045),
            .I(N__46029));
    Span4Mux_v I__10522 (
            .O(N__46042),
            .I(N__46025));
    InMux I__10521 (
            .O(N__46041),
            .I(N__46022));
    Span4Mux_h I__10520 (
            .O(N__46038),
            .I(N__46017));
    Span4Mux_h I__10519 (
            .O(N__46035),
            .I(N__46017));
    LocalMux I__10518 (
            .O(N__46032),
            .I(N__46014));
    LocalMux I__10517 (
            .O(N__46029),
            .I(N__46011));
    CascadeMux I__10516 (
            .O(N__46028),
            .I(N__46008));
    Span4Mux_h I__10515 (
            .O(N__46025),
            .I(N__46005));
    LocalMux I__10514 (
            .O(N__46022),
            .I(N__46002));
    Span4Mux_h I__10513 (
            .O(N__46017),
            .I(N__45997));
    Span4Mux_v I__10512 (
            .O(N__46014),
            .I(N__45997));
    Span4Mux_v I__10511 (
            .O(N__46011),
            .I(N__45994));
    InMux I__10510 (
            .O(N__46008),
            .I(N__45991));
    Span4Mux_h I__10509 (
            .O(N__46005),
            .I(N__45986));
    Span4Mux_h I__10508 (
            .O(N__46002),
            .I(N__45986));
    Sp12to4 I__10507 (
            .O(N__45997),
            .I(N__45983));
    Sp12to4 I__10506 (
            .O(N__45994),
            .I(N__45978));
    LocalMux I__10505 (
            .O(N__45991),
            .I(N__45978));
    Span4Mux_v I__10504 (
            .O(N__45986),
            .I(N__45975));
    Span12Mux_h I__10503 (
            .O(N__45983),
            .I(N__45970));
    Span12Mux_h I__10502 (
            .O(N__45978),
            .I(N__45970));
    Odrv4 I__10501 (
            .O(N__45975),
            .I(comm_buf_0_7));
    Odrv12 I__10500 (
            .O(N__45970),
            .I(comm_buf_0_7));
    InMux I__10499 (
            .O(N__45965),
            .I(N__45962));
    LocalMux I__10498 (
            .O(N__45962),
            .I(n1_adj_1580));
    InMux I__10497 (
            .O(N__45959),
            .I(N__45956));
    LocalMux I__10496 (
            .O(N__45956),
            .I(N__45953));
    Span4Mux_v I__10495 (
            .O(N__45953),
            .I(N__45950));
    Span4Mux_h I__10494 (
            .O(N__45950),
            .I(N__45947));
    Odrv4 I__10493 (
            .O(N__45947),
            .I(comm_buf_5_7));
    InMux I__10492 (
            .O(N__45944),
            .I(N__45941));
    LocalMux I__10491 (
            .O(N__45941),
            .I(N__45938));
    Span4Mux_h I__10490 (
            .O(N__45938),
            .I(N__45935));
    Odrv4 I__10489 (
            .O(N__45935),
            .I(comm_buf_4_7));
    InMux I__10488 (
            .O(N__45932),
            .I(N__45929));
    LocalMux I__10487 (
            .O(N__45929),
            .I(n20966));
    CascadeMux I__10486 (
            .O(N__45926),
            .I(n4_adj_1582_cascade_));
    InMux I__10485 (
            .O(N__45923),
            .I(N__45920));
    LocalMux I__10484 (
            .O(N__45920),
            .I(n21968));
    CascadeMux I__10483 (
            .O(N__45917),
            .I(N__45913));
    InMux I__10482 (
            .O(N__45916),
            .I(N__45908));
    InMux I__10481 (
            .O(N__45913),
            .I(N__45905));
    InMux I__10480 (
            .O(N__45912),
            .I(N__45902));
    InMux I__10479 (
            .O(N__45911),
            .I(N__45899));
    LocalMux I__10478 (
            .O(N__45908),
            .I(N__45896));
    LocalMux I__10477 (
            .O(N__45905),
            .I(N__45893));
    LocalMux I__10476 (
            .O(N__45902),
            .I(N__45890));
    LocalMux I__10475 (
            .O(N__45899),
            .I(N__45887));
    Span4Mux_v I__10474 (
            .O(N__45896),
            .I(N__45883));
    Span4Mux_v I__10473 (
            .O(N__45893),
            .I(N__45880));
    Span4Mux_v I__10472 (
            .O(N__45890),
            .I(N__45877));
    Span4Mux_h I__10471 (
            .O(N__45887),
            .I(N__45874));
    InMux I__10470 (
            .O(N__45886),
            .I(N__45871));
    Sp12to4 I__10469 (
            .O(N__45883),
            .I(N__45868));
    Span4Mux_v I__10468 (
            .O(N__45880),
            .I(N__45863));
    Span4Mux_v I__10467 (
            .O(N__45877),
            .I(N__45863));
    Odrv4 I__10466 (
            .O(N__45874),
            .I(comm_buf_1_5));
    LocalMux I__10465 (
            .O(N__45871),
            .I(comm_buf_1_5));
    Odrv12 I__10464 (
            .O(N__45868),
            .I(comm_buf_1_5));
    Odrv4 I__10463 (
            .O(N__45863),
            .I(comm_buf_1_5));
    InMux I__10462 (
            .O(N__45854),
            .I(N__45851));
    LocalMux I__10461 (
            .O(N__45851),
            .I(N__45848));
    Span4Mux_h I__10460 (
            .O(N__45848),
            .I(N__45845));
    Span4Mux_v I__10459 (
            .O(N__45845),
            .I(N__45842));
    Odrv4 I__10458 (
            .O(N__45842),
            .I(buf_data_iac_9));
    InMux I__10457 (
            .O(N__45839),
            .I(N__45836));
    LocalMux I__10456 (
            .O(N__45836),
            .I(N__45833));
    Odrv4 I__10455 (
            .O(N__45833),
            .I(n21270));
    CascadeMux I__10454 (
            .O(N__45830),
            .I(n22241_cascade_));
    InMux I__10453 (
            .O(N__45827),
            .I(N__45824));
    LocalMux I__10452 (
            .O(N__45824),
            .I(n8_adj_1576));
    InMux I__10451 (
            .O(N__45821),
            .I(N__45815));
    InMux I__10450 (
            .O(N__45820),
            .I(N__45815));
    LocalMux I__10449 (
            .O(N__45815),
            .I(n1272));
    InMux I__10448 (
            .O(N__45812),
            .I(N__45809));
    LocalMux I__10447 (
            .O(N__45809),
            .I(n20697));
    InMux I__10446 (
            .O(N__45806),
            .I(N__45803));
    LocalMux I__10445 (
            .O(N__45803),
            .I(n4_adj_1614));
    InMux I__10444 (
            .O(N__45800),
            .I(N__45794));
    InMux I__10443 (
            .O(N__45799),
            .I(N__45794));
    LocalMux I__10442 (
            .O(N__45794),
            .I(N__45791));
    Odrv12 I__10441 (
            .O(N__45791),
            .I(n20668));
    CEMux I__10440 (
            .O(N__45788),
            .I(N__45785));
    LocalMux I__10439 (
            .O(N__45785),
            .I(N__45782));
    Span4Mux_h I__10438 (
            .O(N__45782),
            .I(N__45779));
    Span4Mux_v I__10437 (
            .O(N__45779),
            .I(N__45776));
    Span4Mux_h I__10436 (
            .O(N__45776),
            .I(N__45773));
    Odrv4 I__10435 (
            .O(N__45773),
            .I(n11866));
    SRMux I__10434 (
            .O(N__45770),
            .I(N__45767));
    LocalMux I__10433 (
            .O(N__45767),
            .I(n14753));
    InMux I__10432 (
            .O(N__45764),
            .I(N__45761));
    LocalMux I__10431 (
            .O(N__45761),
            .I(N__45758));
    Span4Mux_h I__10430 (
            .O(N__45758),
            .I(N__45755));
    Odrv4 I__10429 (
            .O(N__45755),
            .I(n8_adj_1530));
    CascadeMux I__10428 (
            .O(N__45752),
            .I(n4_adj_1598_cascade_));
    CEMux I__10427 (
            .O(N__45749),
            .I(N__45746));
    LocalMux I__10426 (
            .O(N__45746),
            .I(n20573));
    InMux I__10425 (
            .O(N__45743),
            .I(N__45739));
    InMux I__10424 (
            .O(N__45742),
            .I(N__45736));
    LocalMux I__10423 (
            .O(N__45739),
            .I(N__45733));
    LocalMux I__10422 (
            .O(N__45736),
            .I(N__45730));
    Span4Mux_h I__10421 (
            .O(N__45733),
            .I(N__45727));
    Span12Mux_h I__10420 (
            .O(N__45730),
            .I(N__45724));
    Odrv4 I__10419 (
            .O(N__45727),
            .I(comm_state_3_N_420_3));
    Odrv12 I__10418 (
            .O(N__45724),
            .I(comm_state_3_N_420_3));
    CascadeMux I__10417 (
            .O(N__45719),
            .I(n1272_cascade_));
    InMux I__10416 (
            .O(N__45716),
            .I(N__45713));
    LocalMux I__10415 (
            .O(N__45713),
            .I(N__45710));
    Span4Mux_v I__10414 (
            .O(N__45710),
            .I(N__45707));
    Odrv4 I__10413 (
            .O(N__45707),
            .I(comm_buf_4_5));
    InMux I__10412 (
            .O(N__45704),
            .I(N__45701));
    LocalMux I__10411 (
            .O(N__45701),
            .I(n22175));
    InMux I__10410 (
            .O(N__45698),
            .I(N__45695));
    LocalMux I__10409 (
            .O(N__45695),
            .I(n20551));
    InMux I__10408 (
            .O(N__45692),
            .I(N__45689));
    LocalMux I__10407 (
            .O(N__45689),
            .I(N__45686));
    Odrv4 I__10406 (
            .O(N__45686),
            .I(n11420));
    CascadeMux I__10405 (
            .O(N__45683),
            .I(n20551_cascade_));
    InMux I__10404 (
            .O(N__45680),
            .I(N__45677));
    LocalMux I__10403 (
            .O(N__45677),
            .I(N__45674));
    Odrv4 I__10402 (
            .O(N__45674),
            .I(n20717));
    CEMux I__10401 (
            .O(N__45671),
            .I(N__45668));
    LocalMux I__10400 (
            .O(N__45668),
            .I(N__45665));
    Span4Mux_h I__10399 (
            .O(N__45665),
            .I(N__45662));
    Odrv4 I__10398 (
            .O(N__45662),
            .I(n20575));
    InMux I__10397 (
            .O(N__45659),
            .I(N__45656));
    LocalMux I__10396 (
            .O(N__45656),
            .I(N__45653));
    Span4Mux_h I__10395 (
            .O(N__45653),
            .I(N__45650));
    Span4Mux_h I__10394 (
            .O(N__45650),
            .I(N__45647));
    Odrv4 I__10393 (
            .O(N__45647),
            .I(n20962));
    InMux I__10392 (
            .O(N__45644),
            .I(N__45640));
    InMux I__10391 (
            .O(N__45643),
            .I(N__45637));
    LocalMux I__10390 (
            .O(N__45640),
            .I(N__45633));
    LocalMux I__10389 (
            .O(N__45637),
            .I(N__45630));
    CascadeMux I__10388 (
            .O(N__45636),
            .I(N__45627));
    Span4Mux_h I__10387 (
            .O(N__45633),
            .I(N__45622));
    Span4Mux_h I__10386 (
            .O(N__45630),
            .I(N__45622));
    InMux I__10385 (
            .O(N__45627),
            .I(N__45619));
    Odrv4 I__10384 (
            .O(N__45622),
            .I(n14545));
    LocalMux I__10383 (
            .O(N__45619),
            .I(n14545));
    InMux I__10382 (
            .O(N__45614),
            .I(N__45611));
    LocalMux I__10381 (
            .O(N__45611),
            .I(n22238));
    CascadeMux I__10380 (
            .O(N__45608),
            .I(n2_adj_1575_cascade_));
    InMux I__10379 (
            .O(N__45605),
            .I(N__45602));
    LocalMux I__10378 (
            .O(N__45602),
            .I(N__45599));
    Span4Mux_v I__10377 (
            .O(N__45599),
            .I(N__45596));
    Odrv4 I__10376 (
            .O(N__45596),
            .I(comm_buf_2_1));
    InMux I__10375 (
            .O(N__45593),
            .I(N__45590));
    LocalMux I__10374 (
            .O(N__45590),
            .I(N__45587));
    Span4Mux_h I__10373 (
            .O(N__45587),
            .I(N__45584));
    Odrv4 I__10372 (
            .O(N__45584),
            .I(comm_buf_3_1));
    CascadeMux I__10371 (
            .O(N__45581),
            .I(N__45578));
    InMux I__10370 (
            .O(N__45578),
            .I(N__45573));
    CascadeMux I__10369 (
            .O(N__45577),
            .I(N__45570));
    CascadeMux I__10368 (
            .O(N__45576),
            .I(N__45567));
    LocalMux I__10367 (
            .O(N__45573),
            .I(N__45563));
    InMux I__10366 (
            .O(N__45570),
            .I(N__45560));
    InMux I__10365 (
            .O(N__45567),
            .I(N__45557));
    InMux I__10364 (
            .O(N__45566),
            .I(N__45553));
    Span4Mux_v I__10363 (
            .O(N__45563),
            .I(N__45546));
    LocalMux I__10362 (
            .O(N__45560),
            .I(N__45546));
    LocalMux I__10361 (
            .O(N__45557),
            .I(N__45546));
    InMux I__10360 (
            .O(N__45556),
            .I(N__45541));
    LocalMux I__10359 (
            .O(N__45553),
            .I(N__45538));
    Span4Mux_v I__10358 (
            .O(N__45546),
            .I(N__45533));
    InMux I__10357 (
            .O(N__45545),
            .I(N__45530));
    InMux I__10356 (
            .O(N__45544),
            .I(N__45527));
    LocalMux I__10355 (
            .O(N__45541),
            .I(N__45522));
    Span4Mux_v I__10354 (
            .O(N__45538),
            .I(N__45522));
    InMux I__10353 (
            .O(N__45537),
            .I(N__45518));
    InMux I__10352 (
            .O(N__45536),
            .I(N__45515));
    Span4Mux_v I__10351 (
            .O(N__45533),
            .I(N__45510));
    LocalMux I__10350 (
            .O(N__45530),
            .I(N__45510));
    LocalMux I__10349 (
            .O(N__45527),
            .I(N__45505));
    Span4Mux_h I__10348 (
            .O(N__45522),
            .I(N__45505));
    InMux I__10347 (
            .O(N__45521),
            .I(N__45502));
    LocalMux I__10346 (
            .O(N__45518),
            .I(N__45499));
    LocalMux I__10345 (
            .O(N__45515),
            .I(N__45496));
    Span4Mux_v I__10344 (
            .O(N__45510),
            .I(N__45493));
    Sp12to4 I__10343 (
            .O(N__45505),
            .I(N__45488));
    LocalMux I__10342 (
            .O(N__45502),
            .I(N__45488));
    Span4Mux_h I__10341 (
            .O(N__45499),
            .I(N__45485));
    Span12Mux_v I__10340 (
            .O(N__45496),
            .I(N__45482));
    Sp12to4 I__10339 (
            .O(N__45493),
            .I(N__45477));
    Span12Mux_v I__10338 (
            .O(N__45488),
            .I(N__45477));
    Odrv4 I__10337 (
            .O(N__45485),
            .I(comm_buf_0_1));
    Odrv12 I__10336 (
            .O(N__45482),
            .I(comm_buf_0_1));
    Odrv12 I__10335 (
            .O(N__45477),
            .I(comm_buf_0_1));
    CascadeMux I__10334 (
            .O(N__45470),
            .I(n22052_cascade_));
    CascadeMux I__10333 (
            .O(N__45467),
            .I(N__45464));
    InMux I__10332 (
            .O(N__45464),
            .I(N__45461));
    LocalMux I__10331 (
            .O(N__45461),
            .I(N__45458));
    Span4Mux_v I__10330 (
            .O(N__45458),
            .I(N__45450));
    InMux I__10329 (
            .O(N__45457),
            .I(N__45441));
    InMux I__10328 (
            .O(N__45456),
            .I(N__45441));
    InMux I__10327 (
            .O(N__45455),
            .I(N__45441));
    InMux I__10326 (
            .O(N__45454),
            .I(N__45441));
    InMux I__10325 (
            .O(N__45453),
            .I(N__45438));
    Span4Mux_h I__10324 (
            .O(N__45450),
            .I(N__45435));
    LocalMux I__10323 (
            .O(N__45441),
            .I(N__45432));
    LocalMux I__10322 (
            .O(N__45438),
            .I(N__45429));
    Span4Mux_h I__10321 (
            .O(N__45435),
            .I(N__45424));
    Span4Mux_h I__10320 (
            .O(N__45432),
            .I(N__45424));
    Span4Mux_v I__10319 (
            .O(N__45429),
            .I(N__45421));
    Span4Mux_v I__10318 (
            .O(N__45424),
            .I(N__45418));
    Odrv4 I__10317 (
            .O(N__45421),
            .I(comm_buf_1_1));
    Odrv4 I__10316 (
            .O(N__45418),
            .I(comm_buf_1_1));
    InMux I__10315 (
            .O(N__45413),
            .I(N__45410));
    LocalMux I__10314 (
            .O(N__45410),
            .I(n20807));
    CascadeMux I__10313 (
            .O(N__45407),
            .I(n22055_cascade_));
    InMux I__10312 (
            .O(N__45404),
            .I(N__45401));
    LocalMux I__10311 (
            .O(N__45401),
            .I(N__45398));
    Span4Mux_h I__10310 (
            .O(N__45398),
            .I(N__45395));
    Odrv4 I__10309 (
            .O(N__45395),
            .I(comm_buf_5_5));
    InMux I__10308 (
            .O(N__45392),
            .I(N__45389));
    LocalMux I__10307 (
            .O(N__45389),
            .I(N__45386));
    Odrv12 I__10306 (
            .O(N__45386),
            .I(comm_buf_3_5));
    CascadeMux I__10305 (
            .O(N__45383),
            .I(n17404_cascade_));
    CascadeMux I__10304 (
            .O(N__45380),
            .I(n20951_cascade_));
    InMux I__10303 (
            .O(N__45377),
            .I(N__45373));
    CascadeMux I__10302 (
            .O(N__45376),
            .I(N__45369));
    LocalMux I__10301 (
            .O(N__45373),
            .I(N__45366));
    InMux I__10300 (
            .O(N__45372),
            .I(N__45359));
    InMux I__10299 (
            .O(N__45369),
            .I(N__45356));
    Span4Mux_v I__10298 (
            .O(N__45366),
            .I(N__45353));
    InMux I__10297 (
            .O(N__45365),
            .I(N__45350));
    InMux I__10296 (
            .O(N__45364),
            .I(N__45347));
    InMux I__10295 (
            .O(N__45363),
            .I(N__45344));
    InMux I__10294 (
            .O(N__45362),
            .I(N__45341));
    LocalMux I__10293 (
            .O(N__45359),
            .I(N__45338));
    LocalMux I__10292 (
            .O(N__45356),
            .I(N__45335));
    Span4Mux_v I__10291 (
            .O(N__45353),
            .I(N__45330));
    LocalMux I__10290 (
            .O(N__45350),
            .I(N__45330));
    LocalMux I__10289 (
            .O(N__45347),
            .I(N__45323));
    LocalMux I__10288 (
            .O(N__45344),
            .I(N__45323));
    LocalMux I__10287 (
            .O(N__45341),
            .I(N__45323));
    Span4Mux_v I__10286 (
            .O(N__45338),
            .I(N__45318));
    Span4Mux_v I__10285 (
            .O(N__45335),
            .I(N__45315));
    Span4Mux_h I__10284 (
            .O(N__45330),
            .I(N__45312));
    Span4Mux_v I__10283 (
            .O(N__45323),
            .I(N__45309));
    InMux I__10282 (
            .O(N__45322),
            .I(N__45306));
    InMux I__10281 (
            .O(N__45321),
            .I(N__45303));
    Odrv4 I__10280 (
            .O(N__45318),
            .I(comm_rx_buf_1));
    Odrv4 I__10279 (
            .O(N__45315),
            .I(comm_rx_buf_1));
    Odrv4 I__10278 (
            .O(N__45312),
            .I(comm_rx_buf_1));
    Odrv4 I__10277 (
            .O(N__45309),
            .I(comm_rx_buf_1));
    LocalMux I__10276 (
            .O(N__45306),
            .I(comm_rx_buf_1));
    LocalMux I__10275 (
            .O(N__45303),
            .I(comm_rx_buf_1));
    InMux I__10274 (
            .O(N__45290),
            .I(N__45286));
    InMux I__10273 (
            .O(N__45289),
            .I(N__45283));
    LocalMux I__10272 (
            .O(N__45286),
            .I(comm_buf_6_1));
    LocalMux I__10271 (
            .O(N__45283),
            .I(comm_buf_6_1));
    IoInMux I__10270 (
            .O(N__45278),
            .I(N__45275));
    LocalMux I__10269 (
            .O(N__45275),
            .I(N__45272));
    Span4Mux_s3_v I__10268 (
            .O(N__45272),
            .I(N__45269));
    Span4Mux_v I__10267 (
            .O(N__45269),
            .I(N__45266));
    Sp12to4 I__10266 (
            .O(N__45266),
            .I(N__45263));
    Odrv12 I__10265 (
            .O(N__45263),
            .I(DDS_CS));
    CEMux I__10264 (
            .O(N__45260),
            .I(N__45257));
    LocalMux I__10263 (
            .O(N__45257),
            .I(N__45254));
    Span4Mux_v I__10262 (
            .O(N__45254),
            .I(N__45251));
    Span4Mux_h I__10261 (
            .O(N__45251),
            .I(N__45248));
    Odrv4 I__10260 (
            .O(N__45248),
            .I(\SIG_DDS.n9_adj_1394 ));
    InMux I__10259 (
            .O(N__45245),
            .I(N__45242));
    LocalMux I__10258 (
            .O(N__45242),
            .I(N__45239));
    Span4Mux_h I__10257 (
            .O(N__45239),
            .I(N__45236));
    Odrv4 I__10256 (
            .O(N__45236),
            .I(buf_data_iac_20));
    InMux I__10255 (
            .O(N__45233),
            .I(N__45230));
    LocalMux I__10254 (
            .O(N__45230),
            .I(N__45227));
    Span4Mux_h I__10253 (
            .O(N__45227),
            .I(N__45224));
    Odrv4 I__10252 (
            .O(N__45224),
            .I(n20984));
    InMux I__10251 (
            .O(N__45221),
            .I(N__45218));
    LocalMux I__10250 (
            .O(N__45218),
            .I(n17738));
    CascadeMux I__10249 (
            .O(N__45215),
            .I(N__45212));
    InMux I__10248 (
            .O(N__45212),
            .I(N__45209));
    LocalMux I__10247 (
            .O(N__45209),
            .I(n14146));
    CascadeMux I__10246 (
            .O(N__45206),
            .I(N__45202));
    CascadeMux I__10245 (
            .O(N__45205),
            .I(N__45198));
    InMux I__10244 (
            .O(N__45202),
            .I(N__45195));
    InMux I__10243 (
            .O(N__45201),
            .I(N__45188));
    InMux I__10242 (
            .O(N__45198),
            .I(N__45188));
    LocalMux I__10241 (
            .O(N__45195),
            .I(N__45184));
    InMux I__10240 (
            .O(N__45194),
            .I(N__45181));
    InMux I__10239 (
            .O(N__45193),
            .I(N__45178));
    LocalMux I__10238 (
            .O(N__45188),
            .I(N__45175));
    InMux I__10237 (
            .O(N__45187),
            .I(N__45172));
    Span4Mux_v I__10236 (
            .O(N__45184),
            .I(N__45167));
    LocalMux I__10235 (
            .O(N__45181),
            .I(N__45167));
    LocalMux I__10234 (
            .O(N__45178),
            .I(N__45162));
    Span4Mux_h I__10233 (
            .O(N__45175),
            .I(N__45162));
    LocalMux I__10232 (
            .O(N__45172),
            .I(N__45159));
    Span4Mux_v I__10231 (
            .O(N__45167),
            .I(N__45156));
    Span4Mux_v I__10230 (
            .O(N__45162),
            .I(N__45153));
    Span4Mux_h I__10229 (
            .O(N__45159),
            .I(N__45150));
    Sp12to4 I__10228 (
            .O(N__45156),
            .I(N__45147));
    Span4Mux_h I__10227 (
            .O(N__45153),
            .I(N__45144));
    Odrv4 I__10226 (
            .O(N__45150),
            .I(comm_state_3_N_436_2));
    Odrv12 I__10225 (
            .O(N__45147),
            .I(comm_state_3_N_436_2));
    Odrv4 I__10224 (
            .O(N__45144),
            .I(comm_state_3_N_436_2));
    CascadeMux I__10223 (
            .O(N__45137),
            .I(n15_cascade_));
    InMux I__10222 (
            .O(N__45134),
            .I(N__45131));
    LocalMux I__10221 (
            .O(N__45131),
            .I(n12_adj_1649));
    InMux I__10220 (
            .O(N__45128),
            .I(N__45125));
    LocalMux I__10219 (
            .O(N__45125),
            .I(N__45122));
    Span4Mux_h I__10218 (
            .O(N__45122),
            .I(N__45119));
    Odrv4 I__10217 (
            .O(N__45119),
            .I(comm_buf_4_1));
    InMux I__10216 (
            .O(N__45116),
            .I(N__45113));
    LocalMux I__10215 (
            .O(N__45113),
            .I(N__45110));
    Span4Mux_v I__10214 (
            .O(N__45110),
            .I(N__45107));
    Span4Mux_h I__10213 (
            .O(N__45107),
            .I(N__45104));
    Odrv4 I__10212 (
            .O(N__45104),
            .I(comm_buf_5_1));
    CascadeMux I__10211 (
            .O(N__45101),
            .I(n4_adj_1595_cascade_));
    InMux I__10210 (
            .O(N__45098),
            .I(N__45094));
    InMux I__10209 (
            .O(N__45097),
            .I(N__45091));
    LocalMux I__10208 (
            .O(N__45094),
            .I(N__45087));
    LocalMux I__10207 (
            .O(N__45091),
            .I(N__45075));
    ClkMux I__10206 (
            .O(N__45090),
            .I(N__45035));
    Glb2LocalMux I__10205 (
            .O(N__45087),
            .I(N__45035));
    ClkMux I__10204 (
            .O(N__45086),
            .I(N__45035));
    ClkMux I__10203 (
            .O(N__45085),
            .I(N__45035));
    ClkMux I__10202 (
            .O(N__45084),
            .I(N__45035));
    ClkMux I__10201 (
            .O(N__45083),
            .I(N__45035));
    ClkMux I__10200 (
            .O(N__45082),
            .I(N__45035));
    ClkMux I__10199 (
            .O(N__45081),
            .I(N__45035));
    ClkMux I__10198 (
            .O(N__45080),
            .I(N__45035));
    ClkMux I__10197 (
            .O(N__45079),
            .I(N__45035));
    ClkMux I__10196 (
            .O(N__45078),
            .I(N__45035));
    Glb2LocalMux I__10195 (
            .O(N__45075),
            .I(N__45035));
    ClkMux I__10194 (
            .O(N__45074),
            .I(N__45035));
    ClkMux I__10193 (
            .O(N__45073),
            .I(N__45035));
    ClkMux I__10192 (
            .O(N__45072),
            .I(N__45035));
    ClkMux I__10191 (
            .O(N__45071),
            .I(N__45035));
    ClkMux I__10190 (
            .O(N__45070),
            .I(N__45035));
    GlobalMux I__10189 (
            .O(N__45035),
            .I(clk_16MHz));
    InMux I__10188 (
            .O(N__45032),
            .I(N__45029));
    LocalMux I__10187 (
            .O(N__45029),
            .I(N__45025));
    InMux I__10186 (
            .O(N__45028),
            .I(N__45022));
    Odrv4 I__10185 (
            .O(N__45025),
            .I(dds0_mclk));
    LocalMux I__10184 (
            .O(N__45022),
            .I(dds0_mclk));
    InMux I__10183 (
            .O(N__45017),
            .I(N__45013));
    InMux I__10182 (
            .O(N__45016),
            .I(N__45009));
    LocalMux I__10181 (
            .O(N__45013),
            .I(N__45006));
    CascadeMux I__10180 (
            .O(N__45012),
            .I(N__45003));
    LocalMux I__10179 (
            .O(N__45009),
            .I(N__45000));
    Span4Mux_h I__10178 (
            .O(N__45006),
            .I(N__44997));
    InMux I__10177 (
            .O(N__45003),
            .I(N__44994));
    Span12Mux_h I__10176 (
            .O(N__45000),
            .I(N__44989));
    Sp12to4 I__10175 (
            .O(N__44997),
            .I(N__44989));
    LocalMux I__10174 (
            .O(N__44994),
            .I(buf_control_6));
    Odrv12 I__10173 (
            .O(N__44989),
            .I(buf_control_6));
    IoInMux I__10172 (
            .O(N__44984),
            .I(N__44981));
    LocalMux I__10171 (
            .O(N__44981),
            .I(N__44978));
    Span4Mux_s0_v I__10170 (
            .O(N__44978),
            .I(N__44975));
    Span4Mux_v I__10169 (
            .O(N__44975),
            .I(N__44972));
    Sp12to4 I__10168 (
            .O(N__44972),
            .I(N__44969));
    Span12Mux_h I__10167 (
            .O(N__44969),
            .I(N__44966));
    Odrv12 I__10166 (
            .O(N__44966),
            .I(DDS_MCLK));
    InMux I__10165 (
            .O(N__44963),
            .I(N__44960));
    LocalMux I__10164 (
            .O(N__44960),
            .I(N__44956));
    InMux I__10163 (
            .O(N__44959),
            .I(N__44953));
    Span4Mux_h I__10162 (
            .O(N__44956),
            .I(N__44950));
    LocalMux I__10161 (
            .O(N__44953),
            .I(N__44946));
    Span4Mux_h I__10160 (
            .O(N__44950),
            .I(N__44943));
    InMux I__10159 (
            .O(N__44949),
            .I(N__44940));
    Span12Mux_h I__10158 (
            .O(N__44946),
            .I(N__44937));
    Span4Mux_v I__10157 (
            .O(N__44943),
            .I(N__44934));
    LocalMux I__10156 (
            .O(N__44940),
            .I(buf_adcdata_iac_15));
    Odrv12 I__10155 (
            .O(N__44937),
            .I(buf_adcdata_iac_15));
    Odrv4 I__10154 (
            .O(N__44934),
            .I(buf_adcdata_iac_15));
    InMux I__10153 (
            .O(N__44927),
            .I(N__44924));
    LocalMux I__10152 (
            .O(N__44924),
            .I(n16_adj_1503));
    CascadeMux I__10151 (
            .O(N__44921),
            .I(N__44918));
    InMux I__10150 (
            .O(N__44918),
            .I(N__44915));
    LocalMux I__10149 (
            .O(N__44915),
            .I(N__44912));
    Span4Mux_h I__10148 (
            .O(N__44912),
            .I(N__44909));
    Odrv4 I__10147 (
            .O(N__44909),
            .I(n20797));
    InMux I__10146 (
            .O(N__44906),
            .I(N__44902));
    InMux I__10145 (
            .O(N__44905),
            .I(N__44899));
    LocalMux I__10144 (
            .O(N__44902),
            .I(N__44894));
    LocalMux I__10143 (
            .O(N__44899),
            .I(N__44891));
    InMux I__10142 (
            .O(N__44898),
            .I(N__44886));
    InMux I__10141 (
            .O(N__44897),
            .I(N__44886));
    Odrv12 I__10140 (
            .O(N__44894),
            .I(eis_stop));
    Odrv4 I__10139 (
            .O(N__44891),
            .I(eis_stop));
    LocalMux I__10138 (
            .O(N__44886),
            .I(eis_stop));
    InMux I__10137 (
            .O(N__44879),
            .I(N__44876));
    LocalMux I__10136 (
            .O(N__44876),
            .I(N__44873));
    Odrv4 I__10135 (
            .O(N__44873),
            .I(n22034));
    CascadeMux I__10134 (
            .O(N__44870),
            .I(N__44866));
    CascadeMux I__10133 (
            .O(N__44869),
            .I(N__44863));
    InMux I__10132 (
            .O(N__44866),
            .I(N__44854));
    InMux I__10131 (
            .O(N__44863),
            .I(N__44854));
    InMux I__10130 (
            .O(N__44862),
            .I(N__44854));
    InMux I__10129 (
            .O(N__44861),
            .I(N__44851));
    LocalMux I__10128 (
            .O(N__44854),
            .I(\SIG_DDS.bit_cnt_1 ));
    LocalMux I__10127 (
            .O(N__44851),
            .I(\SIG_DDS.bit_cnt_1 ));
    CascadeMux I__10126 (
            .O(N__44846),
            .I(N__44841));
    InMux I__10125 (
            .O(N__44845),
            .I(N__44836));
    InMux I__10124 (
            .O(N__44844),
            .I(N__44836));
    InMux I__10123 (
            .O(N__44841),
            .I(N__44833));
    LocalMux I__10122 (
            .O(N__44836),
            .I(\SIG_DDS.bit_cnt_2 ));
    LocalMux I__10121 (
            .O(N__44833),
            .I(\SIG_DDS.bit_cnt_2 ));
    InMux I__10120 (
            .O(N__44828),
            .I(N__44824));
    InMux I__10119 (
            .O(N__44827),
            .I(N__44821));
    LocalMux I__10118 (
            .O(N__44824),
            .I(\SIG_DDS.bit_cnt_3 ));
    LocalMux I__10117 (
            .O(N__44821),
            .I(\SIG_DDS.bit_cnt_3 ));
    InMux I__10116 (
            .O(N__44816),
            .I(N__44812));
    CascadeMux I__10115 (
            .O(N__44815),
            .I(N__44808));
    LocalMux I__10114 (
            .O(N__44812),
            .I(N__44805));
    CascadeMux I__10113 (
            .O(N__44811),
            .I(N__44802));
    InMux I__10112 (
            .O(N__44808),
            .I(N__44799));
    Span4Mux_v I__10111 (
            .O(N__44805),
            .I(N__44796));
    InMux I__10110 (
            .O(N__44802),
            .I(N__44793));
    LocalMux I__10109 (
            .O(N__44799),
            .I(N__44790));
    Span4Mux_h I__10108 (
            .O(N__44796),
            .I(N__44784));
    LocalMux I__10107 (
            .O(N__44793),
            .I(N__44784));
    Span4Mux_h I__10106 (
            .O(N__44790),
            .I(N__44781));
    InMux I__10105 (
            .O(N__44789),
            .I(N__44778));
    Span4Mux_h I__10104 (
            .O(N__44784),
            .I(N__44775));
    Span4Mux_h I__10103 (
            .O(N__44781),
            .I(N__44772));
    LocalMux I__10102 (
            .O(N__44778),
            .I(trig_dds0));
    Odrv4 I__10101 (
            .O(N__44775),
            .I(trig_dds0));
    Odrv4 I__10100 (
            .O(N__44772),
            .I(trig_dds0));
    SRMux I__10099 (
            .O(N__44765),
            .I(N__44761));
    InMux I__10098 (
            .O(N__44764),
            .I(N__44758));
    LocalMux I__10097 (
            .O(N__44761),
            .I(n14900));
    LocalMux I__10096 (
            .O(N__44758),
            .I(n14900));
    InMux I__10095 (
            .O(N__44753),
            .I(N__44742));
    InMux I__10094 (
            .O(N__44752),
            .I(N__44742));
    InMux I__10093 (
            .O(N__44751),
            .I(N__44742));
    InMux I__10092 (
            .O(N__44750),
            .I(N__44737));
    InMux I__10091 (
            .O(N__44749),
            .I(N__44737));
    LocalMux I__10090 (
            .O(N__44742),
            .I(bit_cnt_0));
    LocalMux I__10089 (
            .O(N__44737),
            .I(bit_cnt_0));
    InMux I__10088 (
            .O(N__44732),
            .I(N__44729));
    LocalMux I__10087 (
            .O(N__44729),
            .I(N__44725));
    CascadeMux I__10086 (
            .O(N__44728),
            .I(N__44722));
    Span4Mux_v I__10085 (
            .O(N__44725),
            .I(N__44719));
    InMux I__10084 (
            .O(N__44722),
            .I(N__44716));
    Span4Mux_h I__10083 (
            .O(N__44719),
            .I(N__44713));
    LocalMux I__10082 (
            .O(N__44716),
            .I(N__44710));
    Odrv4 I__10081 (
            .O(N__44713),
            .I(tmp_buf_15));
    Odrv4 I__10080 (
            .O(N__44710),
            .I(tmp_buf_15));
    IoInMux I__10079 (
            .O(N__44705),
            .I(N__44702));
    LocalMux I__10078 (
            .O(N__44702),
            .I(N__44699));
    Span4Mux_s1_v I__10077 (
            .O(N__44699),
            .I(N__44696));
    Sp12to4 I__10076 (
            .O(N__44696),
            .I(N__44693));
    Span12Mux_h I__10075 (
            .O(N__44693),
            .I(N__44689));
    InMux I__10074 (
            .O(N__44692),
            .I(N__44686));
    Odrv12 I__10073 (
            .O(N__44689),
            .I(DDS_MOSI));
    LocalMux I__10072 (
            .O(N__44686),
            .I(DDS_MOSI));
    InMux I__10071 (
            .O(N__44681),
            .I(N__44678));
    LocalMux I__10070 (
            .O(N__44678),
            .I(N__44675));
    Span4Mux_h I__10069 (
            .O(N__44675),
            .I(N__44672));
    Span4Mux_h I__10068 (
            .O(N__44672),
            .I(N__44669));
    Odrv4 I__10067 (
            .O(N__44669),
            .I(n22226));
    InMux I__10066 (
            .O(N__44666),
            .I(N__44663));
    LocalMux I__10065 (
            .O(N__44663),
            .I(n22229));
    IoInMux I__10064 (
            .O(N__44660),
            .I(N__44657));
    LocalMux I__10063 (
            .O(N__44657),
            .I(N__44654));
    Span4Mux_s0_v I__10062 (
            .O(N__44654),
            .I(N__44650));
    CascadeMux I__10061 (
            .O(N__44653),
            .I(N__44647));
    Span4Mux_v I__10060 (
            .O(N__44650),
            .I(N__44644));
    InMux I__10059 (
            .O(N__44647),
            .I(N__44640));
    Sp12to4 I__10058 (
            .O(N__44644),
            .I(N__44637));
    CascadeMux I__10057 (
            .O(N__44643),
            .I(N__44634));
    LocalMux I__10056 (
            .O(N__44640),
            .I(N__44631));
    Span12Mux_h I__10055 (
            .O(N__44637),
            .I(N__44628));
    InMux I__10054 (
            .O(N__44634),
            .I(N__44625));
    Span4Mux_h I__10053 (
            .O(N__44631),
            .I(N__44622));
    Odrv12 I__10052 (
            .O(N__44628),
            .I(DDS_RNG_0));
    LocalMux I__10051 (
            .O(N__44625),
            .I(DDS_RNG_0));
    Odrv4 I__10050 (
            .O(N__44622),
            .I(DDS_RNG_0));
    InMux I__10049 (
            .O(N__44615),
            .I(N__44612));
    LocalMux I__10048 (
            .O(N__44612),
            .I(N__44609));
    Span4Mux_h I__10047 (
            .O(N__44609),
            .I(N__44604));
    InMux I__10046 (
            .O(N__44608),
            .I(N__44599));
    InMux I__10045 (
            .O(N__44607),
            .I(N__44599));
    Odrv4 I__10044 (
            .O(N__44604),
            .I(acadc_skipCount_9));
    LocalMux I__10043 (
            .O(N__44599),
            .I(acadc_skipCount_9));
    InMux I__10042 (
            .O(N__44594),
            .I(N__44591));
    LocalMux I__10041 (
            .O(N__44591),
            .I(n22037));
    InMux I__10040 (
            .O(N__44588),
            .I(N__44583));
    InMux I__10039 (
            .O(N__44587),
            .I(N__44580));
    InMux I__10038 (
            .O(N__44586),
            .I(N__44577));
    LocalMux I__10037 (
            .O(N__44583),
            .I(N__44572));
    LocalMux I__10036 (
            .O(N__44580),
            .I(N__44572));
    LocalMux I__10035 (
            .O(N__44577),
            .I(buf_dds1_7));
    Odrv12 I__10034 (
            .O(N__44572),
            .I(buf_dds1_7));
    InMux I__10033 (
            .O(N__44567),
            .I(N__44564));
    LocalMux I__10032 (
            .O(N__44564),
            .I(N__44559));
    InMux I__10031 (
            .O(N__44563),
            .I(N__44556));
    InMux I__10030 (
            .O(N__44562),
            .I(N__44553));
    Span4Mux_v I__10029 (
            .O(N__44559),
            .I(N__44550));
    LocalMux I__10028 (
            .O(N__44556),
            .I(N__44547));
    LocalMux I__10027 (
            .O(N__44553),
            .I(buf_dds0_7));
    Odrv4 I__10026 (
            .O(N__44550),
            .I(buf_dds0_7));
    Odrv12 I__10025 (
            .O(N__44547),
            .I(buf_dds0_7));
    CascadeMux I__10024 (
            .O(N__44540),
            .I(N__44537));
    InMux I__10023 (
            .O(N__44537),
            .I(N__44533));
    CascadeMux I__10022 (
            .O(N__44536),
            .I(N__44530));
    LocalMux I__10021 (
            .O(N__44533),
            .I(N__44526));
    InMux I__10020 (
            .O(N__44530),
            .I(N__44523));
    InMux I__10019 (
            .O(N__44529),
            .I(N__44520));
    Span4Mux_h I__10018 (
            .O(N__44526),
            .I(N__44517));
    LocalMux I__10017 (
            .O(N__44523),
            .I(N__44514));
    LocalMux I__10016 (
            .O(N__44520),
            .I(req_data_cnt_11));
    Odrv4 I__10015 (
            .O(N__44517),
            .I(req_data_cnt_11));
    Odrv4 I__10014 (
            .O(N__44514),
            .I(req_data_cnt_11));
    InMux I__10013 (
            .O(N__44507),
            .I(N__44504));
    LocalMux I__10012 (
            .O(N__44504),
            .I(n23_adj_1540));
    InMux I__10011 (
            .O(N__44501),
            .I(N__44498));
    LocalMux I__10010 (
            .O(N__44498),
            .I(N__44495));
    Sp12to4 I__10009 (
            .O(N__44495),
            .I(N__44492));
    Odrv12 I__10008 (
            .O(N__44492),
            .I(n20836));
    CascadeMux I__10007 (
            .O(N__44489),
            .I(N__44485));
    InMux I__10006 (
            .O(N__44488),
            .I(N__44482));
    InMux I__10005 (
            .O(N__44485),
            .I(N__44479));
    LocalMux I__10004 (
            .O(N__44482),
            .I(N__44474));
    LocalMux I__10003 (
            .O(N__44479),
            .I(N__44471));
    InMux I__10002 (
            .O(N__44478),
            .I(N__44468));
    InMux I__10001 (
            .O(N__44477),
            .I(N__44464));
    Span4Mux_v I__10000 (
            .O(N__44474),
            .I(N__44457));
    Span4Mux_v I__9999 (
            .O(N__44471),
            .I(N__44457));
    LocalMux I__9998 (
            .O(N__44468),
            .I(N__44457));
    InMux I__9997 (
            .O(N__44467),
            .I(N__44454));
    LocalMux I__9996 (
            .O(N__44464),
            .I(N__44451));
    Span4Mux_h I__9995 (
            .O(N__44457),
            .I(N__44448));
    LocalMux I__9994 (
            .O(N__44454),
            .I(n14_adj_1545));
    Odrv4 I__9993 (
            .O(N__44451),
            .I(n14_adj_1545));
    Odrv4 I__9992 (
            .O(N__44448),
            .I(n14_adj_1545));
    InMux I__9991 (
            .O(N__44441),
            .I(N__44435));
    CascadeMux I__9990 (
            .O(N__44440),
            .I(N__44431));
    InMux I__9989 (
            .O(N__44439),
            .I(N__44426));
    InMux I__9988 (
            .O(N__44438),
            .I(N__44423));
    LocalMux I__9987 (
            .O(N__44435),
            .I(N__44420));
    InMux I__9986 (
            .O(N__44434),
            .I(N__44415));
    InMux I__9985 (
            .O(N__44431),
            .I(N__44415));
    InMux I__9984 (
            .O(N__44430),
            .I(N__44410));
    InMux I__9983 (
            .O(N__44429),
            .I(N__44410));
    LocalMux I__9982 (
            .O(N__44426),
            .I(N__44405));
    LocalMux I__9981 (
            .O(N__44423),
            .I(N__44405));
    Span4Mux_h I__9980 (
            .O(N__44420),
            .I(N__44402));
    LocalMux I__9979 (
            .O(N__44415),
            .I(N__44399));
    LocalMux I__9978 (
            .O(N__44410),
            .I(N__44396));
    Span4Mux_h I__9977 (
            .O(N__44405),
            .I(N__44393));
    Span4Mux_h I__9976 (
            .O(N__44402),
            .I(N__44390));
    Span4Mux_h I__9975 (
            .O(N__44399),
            .I(N__44387));
    Span4Mux_v I__9974 (
            .O(N__44396),
            .I(N__44382));
    Span4Mux_v I__9973 (
            .O(N__44393),
            .I(N__44382));
    Odrv4 I__9972 (
            .O(N__44390),
            .I(n11931));
    Odrv4 I__9971 (
            .O(N__44387),
            .I(n11931));
    Odrv4 I__9970 (
            .O(N__44382),
            .I(n11931));
    CascadeMux I__9969 (
            .O(N__44375),
            .I(n21073_cascade_));
    CascadeMux I__9968 (
            .O(N__44372),
            .I(n21072_cascade_));
    InMux I__9967 (
            .O(N__44369),
            .I(N__44366));
    LocalMux I__9966 (
            .O(N__44366),
            .I(n23));
    InMux I__9965 (
            .O(N__44363),
            .I(N__44360));
    LocalMux I__9964 (
            .O(N__44360),
            .I(n21_adj_1521));
    CascadeMux I__9963 (
            .O(N__44357),
            .I(n22_adj_1568_cascade_));
    InMux I__9962 (
            .O(N__44354),
            .I(N__44351));
    LocalMux I__9961 (
            .O(N__44351),
            .I(n30_adj_1641));
    InMux I__9960 (
            .O(N__44348),
            .I(N__44344));
    CascadeMux I__9959 (
            .O(N__44347),
            .I(N__44341));
    LocalMux I__9958 (
            .O(N__44344),
            .I(N__44338));
    InMux I__9957 (
            .O(N__44341),
            .I(N__44335));
    Span4Mux_h I__9956 (
            .O(N__44338),
            .I(N__44332));
    LocalMux I__9955 (
            .O(N__44335),
            .I(data_idxvec_9));
    Odrv4 I__9954 (
            .O(N__44332),
            .I(data_idxvec_9));
    InMux I__9953 (
            .O(N__44327),
            .I(N__44324));
    LocalMux I__9952 (
            .O(N__44324),
            .I(N__44321));
    Span4Mux_h I__9951 (
            .O(N__44321),
            .I(N__44318));
    Span4Mux_h I__9950 (
            .O(N__44318),
            .I(N__44315));
    Odrv4 I__9949 (
            .O(N__44315),
            .I(buf_data_iac_17));
    CascadeMux I__9948 (
            .O(N__44312),
            .I(n20812_cascade_));
    CascadeMux I__9947 (
            .O(N__44309),
            .I(N__44304));
    InMux I__9946 (
            .O(N__44308),
            .I(N__44298));
    InMux I__9945 (
            .O(N__44307),
            .I(N__44295));
    InMux I__9944 (
            .O(N__44304),
            .I(N__44292));
    CascadeMux I__9943 (
            .O(N__44303),
            .I(N__44288));
    CascadeMux I__9942 (
            .O(N__44302),
            .I(N__44285));
    CascadeMux I__9941 (
            .O(N__44301),
            .I(N__44282));
    LocalMux I__9940 (
            .O(N__44298),
            .I(N__44278));
    LocalMux I__9939 (
            .O(N__44295),
            .I(N__44275));
    LocalMux I__9938 (
            .O(N__44292),
            .I(N__44272));
    InMux I__9937 (
            .O(N__44291),
            .I(N__44269));
    InMux I__9936 (
            .O(N__44288),
            .I(N__44266));
    InMux I__9935 (
            .O(N__44285),
            .I(N__44263));
    InMux I__9934 (
            .O(N__44282),
            .I(N__44260));
    InMux I__9933 (
            .O(N__44281),
            .I(N__44256));
    Span4Mux_h I__9932 (
            .O(N__44278),
            .I(N__44253));
    Span4Mux_h I__9931 (
            .O(N__44275),
            .I(N__44248));
    Span4Mux_v I__9930 (
            .O(N__44272),
            .I(N__44248));
    LocalMux I__9929 (
            .O(N__44269),
            .I(N__44245));
    LocalMux I__9928 (
            .O(N__44266),
            .I(N__44242));
    LocalMux I__9927 (
            .O(N__44263),
            .I(N__44239));
    LocalMux I__9926 (
            .O(N__44260),
            .I(N__44236));
    InMux I__9925 (
            .O(N__44259),
            .I(N__44233));
    LocalMux I__9924 (
            .O(N__44256),
            .I(N__44228));
    Span4Mux_v I__9923 (
            .O(N__44253),
            .I(N__44228));
    Span4Mux_v I__9922 (
            .O(N__44248),
            .I(N__44223));
    Span4Mux_h I__9921 (
            .O(N__44245),
            .I(N__44223));
    Span4Mux_v I__9920 (
            .O(N__44242),
            .I(N__44220));
    Span4Mux_h I__9919 (
            .O(N__44239),
            .I(N__44215));
    Span4Mux_v I__9918 (
            .O(N__44236),
            .I(N__44215));
    LocalMux I__9917 (
            .O(N__44233),
            .I(N__44208));
    Span4Mux_h I__9916 (
            .O(N__44228),
            .I(N__44208));
    Span4Mux_h I__9915 (
            .O(N__44223),
            .I(N__44208));
    Odrv4 I__9914 (
            .O(N__44220),
            .I(comm_buf_0_3));
    Odrv4 I__9913 (
            .O(N__44215),
            .I(comm_buf_0_3));
    Odrv4 I__9912 (
            .O(N__44208),
            .I(comm_buf_0_3));
    IoInMux I__9911 (
            .O(N__44201),
            .I(N__44198));
    LocalMux I__9910 (
            .O(N__44198),
            .I(N__44194));
    InMux I__9909 (
            .O(N__44197),
            .I(N__44190));
    Span12Mux_s3_v I__9908 (
            .O(N__44194),
            .I(N__44187));
    InMux I__9907 (
            .O(N__44193),
            .I(N__44184));
    LocalMux I__9906 (
            .O(N__44190),
            .I(N__44181));
    Odrv12 I__9905 (
            .O(N__44187),
            .I(SELIRNG1));
    LocalMux I__9904 (
            .O(N__44184),
            .I(SELIRNG1));
    Odrv4 I__9903 (
            .O(N__44181),
            .I(SELIRNG1));
    CascadeMux I__9902 (
            .O(N__44174),
            .I(N__44170));
    InMux I__9901 (
            .O(N__44173),
            .I(N__44165));
    InMux I__9900 (
            .O(N__44170),
            .I(N__44162));
    CascadeMux I__9899 (
            .O(N__44169),
            .I(N__44159));
    CascadeMux I__9898 (
            .O(N__44168),
            .I(N__44156));
    LocalMux I__9897 (
            .O(N__44165),
            .I(N__44152));
    LocalMux I__9896 (
            .O(N__44162),
            .I(N__44149));
    InMux I__9895 (
            .O(N__44159),
            .I(N__44146));
    InMux I__9894 (
            .O(N__44156),
            .I(N__44143));
    InMux I__9893 (
            .O(N__44155),
            .I(N__44140));
    Span4Mux_h I__9892 (
            .O(N__44152),
            .I(N__44136));
    Span4Mux_v I__9891 (
            .O(N__44149),
            .I(N__44133));
    LocalMux I__9890 (
            .O(N__44146),
            .I(N__44128));
    LocalMux I__9889 (
            .O(N__44143),
            .I(N__44128));
    LocalMux I__9888 (
            .O(N__44140),
            .I(N__44124));
    InMux I__9887 (
            .O(N__44139),
            .I(N__44121));
    Span4Mux_h I__9886 (
            .O(N__44136),
            .I(N__44113));
    Span4Mux_h I__9885 (
            .O(N__44133),
            .I(N__44113));
    Span4Mux_h I__9884 (
            .O(N__44128),
            .I(N__44113));
    InMux I__9883 (
            .O(N__44127),
            .I(N__44110));
    Span4Mux_h I__9882 (
            .O(N__44124),
            .I(N__44105));
    LocalMux I__9881 (
            .O(N__44121),
            .I(N__44105));
    InMux I__9880 (
            .O(N__44120),
            .I(N__44102));
    Span4Mux_v I__9879 (
            .O(N__44113),
            .I(N__44099));
    LocalMux I__9878 (
            .O(N__44110),
            .I(N__44094));
    Span4Mux_v I__9877 (
            .O(N__44105),
            .I(N__44094));
    LocalMux I__9876 (
            .O(N__44102),
            .I(N__44091));
    Span4Mux_v I__9875 (
            .O(N__44099),
            .I(N__44088));
    Span4Mux_v I__9874 (
            .O(N__44094),
            .I(N__44085));
    Odrv4 I__9873 (
            .O(N__44091),
            .I(comm_buf_0_4));
    Odrv4 I__9872 (
            .O(N__44088),
            .I(comm_buf_0_4));
    Odrv4 I__9871 (
            .O(N__44085),
            .I(comm_buf_0_4));
    InMux I__9870 (
            .O(N__44078),
            .I(N__44074));
    InMux I__9869 (
            .O(N__44077),
            .I(N__44071));
    LocalMux I__9868 (
            .O(N__44074),
            .I(N__44068));
    LocalMux I__9867 (
            .O(N__44071),
            .I(N__44065));
    Span4Mux_v I__9866 (
            .O(N__44068),
            .I(N__44062));
    Span12Mux_h I__9865 (
            .O(N__44065),
            .I(N__44059));
    Odrv4 I__9864 (
            .O(N__44062),
            .I(n14_adj_1571));
    Odrv12 I__9863 (
            .O(N__44059),
            .I(n14_adj_1571));
    InMux I__9862 (
            .O(N__44054),
            .I(N__44051));
    LocalMux I__9861 (
            .O(N__44051),
            .I(N__44047));
    InMux I__9860 (
            .O(N__44050),
            .I(N__44044));
    Span4Mux_h I__9859 (
            .O(N__44047),
            .I(N__44041));
    LocalMux I__9858 (
            .O(N__44044),
            .I(N__44038));
    Span4Mux_h I__9857 (
            .O(N__44041),
            .I(N__44035));
    Span4Mux_v I__9856 (
            .O(N__44038),
            .I(N__44032));
    Span4Mux_v I__9855 (
            .O(N__44035),
            .I(N__44029));
    Odrv4 I__9854 (
            .O(N__44032),
            .I(n14_adj_1549));
    Odrv4 I__9853 (
            .O(N__44029),
            .I(n14_adj_1549));
    InMux I__9852 (
            .O(N__44024),
            .I(N__44021));
    LocalMux I__9851 (
            .O(N__44021),
            .I(n20814));
    InMux I__9850 (
            .O(N__44018),
            .I(N__44015));
    LocalMux I__9849 (
            .O(N__44015),
            .I(N__44012));
    Span4Mux_h I__9848 (
            .O(N__44012),
            .I(N__44009));
    Odrv4 I__9847 (
            .O(N__44009),
            .I(n22025));
    CascadeMux I__9846 (
            .O(N__44006),
            .I(n22232_cascade_));
    InMux I__9845 (
            .O(N__44003),
            .I(N__44000));
    LocalMux I__9844 (
            .O(N__44000),
            .I(N__43997));
    Span12Mux_v I__9843 (
            .O(N__43997),
            .I(N__43994));
    Odrv12 I__9842 (
            .O(N__43994),
            .I(n22235));
    InMux I__9841 (
            .O(N__43991),
            .I(N__43988));
    LocalMux I__9840 (
            .O(N__43988),
            .I(N__43985));
    Span4Mux_v I__9839 (
            .O(N__43985),
            .I(N__43982));
    Sp12to4 I__9838 (
            .O(N__43982),
            .I(N__43979));
    Span12Mux_h I__9837 (
            .O(N__43979),
            .I(N__43975));
    InMux I__9836 (
            .O(N__43978),
            .I(N__43972));
    Odrv12 I__9835 (
            .O(N__43975),
            .I(buf_adcdata_vdc_17));
    LocalMux I__9834 (
            .O(N__43972),
            .I(buf_adcdata_vdc_17));
    InMux I__9833 (
            .O(N__43967),
            .I(N__43964));
    LocalMux I__9832 (
            .O(N__43964),
            .I(N__43961));
    Span4Mux_h I__9831 (
            .O(N__43961),
            .I(N__43957));
    CascadeMux I__9830 (
            .O(N__43960),
            .I(N__43954));
    Span4Mux_v I__9829 (
            .O(N__43957),
            .I(N__43951));
    InMux I__9828 (
            .O(N__43954),
            .I(N__43948));
    Sp12to4 I__9827 (
            .O(N__43951),
            .I(N__43942));
    LocalMux I__9826 (
            .O(N__43948),
            .I(N__43942));
    InMux I__9825 (
            .O(N__43947),
            .I(N__43939));
    Span12Mux_h I__9824 (
            .O(N__43942),
            .I(N__43936));
    LocalMux I__9823 (
            .O(N__43939),
            .I(buf_adcdata_vac_17));
    Odrv12 I__9822 (
            .O(N__43936),
            .I(buf_adcdata_vac_17));
    CascadeMux I__9821 (
            .O(N__43931),
            .I(n19_adj_1597_cascade_));
    CascadeMux I__9820 (
            .O(N__43928),
            .I(n29_adj_1635_cascade_));
    InMux I__9819 (
            .O(N__43925),
            .I(N__43921));
    CascadeMux I__9818 (
            .O(N__43924),
            .I(N__43917));
    LocalMux I__9817 (
            .O(N__43921),
            .I(N__43914));
    InMux I__9816 (
            .O(N__43920),
            .I(N__43909));
    InMux I__9815 (
            .O(N__43917),
            .I(N__43909));
    Span4Mux_v I__9814 (
            .O(N__43914),
            .I(N__43904));
    LocalMux I__9813 (
            .O(N__43909),
            .I(N__43904));
    Odrv4 I__9812 (
            .O(N__43904),
            .I(n16_adj_1623));
    InMux I__9811 (
            .O(N__43901),
            .I(N__43896));
    InMux I__9810 (
            .O(N__43900),
            .I(N__43891));
    InMux I__9809 (
            .O(N__43899),
            .I(N__43891));
    LocalMux I__9808 (
            .O(N__43896),
            .I(req_data_cnt_8));
    LocalMux I__9807 (
            .O(N__43891),
            .I(req_data_cnt_8));
    InMux I__9806 (
            .O(N__43886),
            .I(N__43883));
    LocalMux I__9805 (
            .O(N__43883),
            .I(N__43880));
    Span4Mux_h I__9804 (
            .O(N__43880),
            .I(N__43875));
    InMux I__9803 (
            .O(N__43879),
            .I(N__43872));
    InMux I__9802 (
            .O(N__43878),
            .I(N__43869));
    Odrv4 I__9801 (
            .O(N__43875),
            .I(n10534));
    LocalMux I__9800 (
            .O(N__43872),
            .I(n10534));
    LocalMux I__9799 (
            .O(N__43869),
            .I(n10534));
    InMux I__9798 (
            .O(N__43862),
            .I(N__43859));
    LocalMux I__9797 (
            .O(N__43859),
            .I(N__43856));
    Span4Mux_h I__9796 (
            .O(N__43856),
            .I(N__43853));
    Odrv4 I__9795 (
            .O(N__43853),
            .I(n20798));
    InMux I__9794 (
            .O(N__43850),
            .I(N__43847));
    LocalMux I__9793 (
            .O(N__43847),
            .I(N__43844));
    Span4Mux_h I__9792 (
            .O(N__43844),
            .I(N__43841));
    Odrv4 I__9791 (
            .O(N__43841),
            .I(n22061));
    SRMux I__9790 (
            .O(N__43838),
            .I(N__43834));
    InMux I__9789 (
            .O(N__43837),
            .I(N__43831));
    LocalMux I__9788 (
            .O(N__43834),
            .I(N__43828));
    LocalMux I__9787 (
            .O(N__43831),
            .I(N__43825));
    Odrv12 I__9786 (
            .O(N__43828),
            .I(n14730));
    Odrv4 I__9785 (
            .O(N__43825),
            .I(n14730));
    ClkMux I__9784 (
            .O(N__43820),
            .I(N__43817));
    LocalMux I__9783 (
            .O(N__43817),
            .I(N__43810));
    ClkMux I__9782 (
            .O(N__43816),
            .I(N__43807));
    ClkMux I__9781 (
            .O(N__43815),
            .I(N__43801));
    ClkMux I__9780 (
            .O(N__43814),
            .I(N__43798));
    ClkMux I__9779 (
            .O(N__43813),
            .I(N__43795));
    Span4Mux_v I__9778 (
            .O(N__43810),
            .I(N__43790));
    LocalMux I__9777 (
            .O(N__43807),
            .I(N__43790));
    ClkMux I__9776 (
            .O(N__43806),
            .I(N__43787));
    ClkMux I__9775 (
            .O(N__43805),
            .I(N__43784));
    ClkMux I__9774 (
            .O(N__43804),
            .I(N__43781));
    LocalMux I__9773 (
            .O(N__43801),
            .I(N__43776));
    LocalMux I__9772 (
            .O(N__43798),
            .I(N__43773));
    LocalMux I__9771 (
            .O(N__43795),
            .I(N__43762));
    Span4Mux_h I__9770 (
            .O(N__43790),
            .I(N__43762));
    LocalMux I__9769 (
            .O(N__43787),
            .I(N__43762));
    LocalMux I__9768 (
            .O(N__43784),
            .I(N__43762));
    LocalMux I__9767 (
            .O(N__43781),
            .I(N__43762));
    ClkMux I__9766 (
            .O(N__43780),
            .I(N__43755));
    ClkMux I__9765 (
            .O(N__43779),
            .I(N__43752));
    Span4Mux_v I__9764 (
            .O(N__43776),
            .I(N__43749));
    Span4Mux_v I__9763 (
            .O(N__43773),
            .I(N__43744));
    Span4Mux_v I__9762 (
            .O(N__43762),
            .I(N__43744));
    ClkMux I__9761 (
            .O(N__43761),
            .I(N__43741));
    ClkMux I__9760 (
            .O(N__43760),
            .I(N__43737));
    ClkMux I__9759 (
            .O(N__43759),
            .I(N__43732));
    ClkMux I__9758 (
            .O(N__43758),
            .I(N__43729));
    LocalMux I__9757 (
            .O(N__43755),
            .I(N__43726));
    LocalMux I__9756 (
            .O(N__43752),
            .I(N__43723));
    Span4Mux_h I__9755 (
            .O(N__43749),
            .I(N__43718));
    Span4Mux_h I__9754 (
            .O(N__43744),
            .I(N__43718));
    LocalMux I__9753 (
            .O(N__43741),
            .I(N__43715));
    ClkMux I__9752 (
            .O(N__43740),
            .I(N__43712));
    LocalMux I__9751 (
            .O(N__43737),
            .I(N__43709));
    ClkMux I__9750 (
            .O(N__43736),
            .I(N__43706));
    ClkMux I__9749 (
            .O(N__43735),
            .I(N__43703));
    LocalMux I__9748 (
            .O(N__43732),
            .I(N__43698));
    LocalMux I__9747 (
            .O(N__43729),
            .I(N__43698));
    Span4Mux_h I__9746 (
            .O(N__43726),
            .I(N__43693));
    Span4Mux_h I__9745 (
            .O(N__43723),
            .I(N__43693));
    Span4Mux_h I__9744 (
            .O(N__43718),
            .I(N__43688));
    Span4Mux_h I__9743 (
            .O(N__43715),
            .I(N__43688));
    LocalMux I__9742 (
            .O(N__43712),
            .I(N__43685));
    Span4Mux_h I__9741 (
            .O(N__43709),
            .I(N__43680));
    LocalMux I__9740 (
            .O(N__43706),
            .I(N__43680));
    LocalMux I__9739 (
            .O(N__43703),
            .I(N__43677));
    Span4Mux_v I__9738 (
            .O(N__43698),
            .I(N__43674));
    Span4Mux_h I__9737 (
            .O(N__43693),
            .I(N__43671));
    Sp12to4 I__9736 (
            .O(N__43688),
            .I(N__43668));
    Span4Mux_h I__9735 (
            .O(N__43685),
            .I(N__43663));
    Span4Mux_h I__9734 (
            .O(N__43680),
            .I(N__43663));
    Span4Mux_h I__9733 (
            .O(N__43677),
            .I(N__43660));
    Span4Mux_h I__9732 (
            .O(N__43674),
            .I(N__43657));
    Span4Mux_v I__9731 (
            .O(N__43671),
            .I(N__43653));
    Span12Mux_h I__9730 (
            .O(N__43668),
            .I(N__43650));
    Span4Mux_h I__9729 (
            .O(N__43663),
            .I(N__43647));
    Span4Mux_v I__9728 (
            .O(N__43660),
            .I(N__43644));
    Span4Mux_h I__9727 (
            .O(N__43657),
            .I(N__43641));
    InMux I__9726 (
            .O(N__43656),
            .I(N__43638));
    Odrv4 I__9725 (
            .O(N__43653),
            .I(clk_RTD));
    Odrv12 I__9724 (
            .O(N__43650),
            .I(clk_RTD));
    Odrv4 I__9723 (
            .O(N__43647),
            .I(clk_RTD));
    Odrv4 I__9722 (
            .O(N__43644),
            .I(clk_RTD));
    Odrv4 I__9721 (
            .O(N__43641),
            .I(clk_RTD));
    LocalMux I__9720 (
            .O(N__43638),
            .I(clk_RTD));
    CascadeMux I__9719 (
            .O(N__43625),
            .I(n22064_cascade_));
    InMux I__9718 (
            .O(N__43622),
            .I(N__43619));
    LocalMux I__9717 (
            .O(N__43619),
            .I(N__43616));
    Span4Mux_h I__9716 (
            .O(N__43616),
            .I(N__43613));
    Span4Mux_h I__9715 (
            .O(N__43613),
            .I(N__43610));
    Odrv4 I__9714 (
            .O(N__43610),
            .I(n16_adj_1519));
    InMux I__9713 (
            .O(N__43607),
            .I(N__43604));
    LocalMux I__9712 (
            .O(N__43604),
            .I(n22067));
    InMux I__9711 (
            .O(N__43601),
            .I(N__43597));
    CascadeMux I__9710 (
            .O(N__43600),
            .I(N__43594));
    LocalMux I__9709 (
            .O(N__43597),
            .I(N__43591));
    InMux I__9708 (
            .O(N__43594),
            .I(N__43588));
    Odrv12 I__9707 (
            .O(N__43591),
            .I(buf_readRTD_5));
    LocalMux I__9706 (
            .O(N__43588),
            .I(buf_readRTD_5));
    InMux I__9705 (
            .O(N__43583),
            .I(N__43580));
    LocalMux I__9704 (
            .O(N__43580),
            .I(N__43575));
    InMux I__9703 (
            .O(N__43579),
            .I(N__43572));
    CascadeMux I__9702 (
            .O(N__43578),
            .I(N__43569));
    Span4Mux_h I__9701 (
            .O(N__43575),
            .I(N__43566));
    LocalMux I__9700 (
            .O(N__43572),
            .I(N__43563));
    InMux I__9699 (
            .O(N__43569),
            .I(N__43560));
    Span4Mux_h I__9698 (
            .O(N__43566),
            .I(N__43557));
    Span12Mux_h I__9697 (
            .O(N__43563),
            .I(N__43554));
    LocalMux I__9696 (
            .O(N__43560),
            .I(buf_adcdata_iac_13));
    Odrv4 I__9695 (
            .O(N__43557),
            .I(buf_adcdata_iac_13));
    Odrv12 I__9694 (
            .O(N__43554),
            .I(buf_adcdata_iac_13));
    CascadeMux I__9693 (
            .O(N__43547),
            .I(n22142_cascade_));
    InMux I__9692 (
            .O(N__43544),
            .I(N__43541));
    LocalMux I__9691 (
            .O(N__43541),
            .I(N__43538));
    Span4Mux_h I__9690 (
            .O(N__43538),
            .I(N__43535));
    Span4Mux_v I__9689 (
            .O(N__43535),
            .I(N__43532));
    Odrv4 I__9688 (
            .O(N__43532),
            .I(n16_adj_1496));
    InMux I__9687 (
            .O(N__43529),
            .I(N__43525));
    CascadeMux I__9686 (
            .O(N__43528),
            .I(N__43521));
    LocalMux I__9685 (
            .O(N__43525),
            .I(N__43518));
    InMux I__9684 (
            .O(N__43524),
            .I(N__43515));
    InMux I__9683 (
            .O(N__43521),
            .I(N__43512));
    Span4Mux_h I__9682 (
            .O(N__43518),
            .I(N__43507));
    LocalMux I__9681 (
            .O(N__43515),
            .I(N__43507));
    LocalMux I__9680 (
            .O(N__43512),
            .I(acadc_skipCount_5));
    Odrv4 I__9679 (
            .O(N__43507),
            .I(acadc_skipCount_5));
    InMux I__9678 (
            .O(N__43502),
            .I(N__43499));
    LocalMux I__9677 (
            .O(N__43499),
            .I(n22145));
    CascadeMux I__9676 (
            .O(N__43496),
            .I(n22133_cascade_));
    CascadeMux I__9675 (
            .O(N__43493),
            .I(n30_adj_1499_cascade_));
    InMux I__9674 (
            .O(N__43490),
            .I(N__43486));
    CascadeMux I__9673 (
            .O(N__43489),
            .I(N__43483));
    LocalMux I__9672 (
            .O(N__43486),
            .I(N__43480));
    InMux I__9671 (
            .O(N__43483),
            .I(N__43477));
    Span4Mux_v I__9670 (
            .O(N__43480),
            .I(N__43474));
    LocalMux I__9669 (
            .O(N__43477),
            .I(data_idxvec_5));
    Odrv4 I__9668 (
            .O(N__43474),
            .I(data_idxvec_5));
    CascadeMux I__9667 (
            .O(N__43469),
            .I(n26_adj_1498_cascade_));
    InMux I__9666 (
            .O(N__43466),
            .I(N__43463));
    LocalMux I__9665 (
            .O(N__43463),
            .I(n22130));
    InMux I__9664 (
            .O(N__43460),
            .I(N__43455));
    InMux I__9663 (
            .O(N__43459),
            .I(N__43452));
    InMux I__9662 (
            .O(N__43458),
            .I(N__43449));
    LocalMux I__9661 (
            .O(N__43455),
            .I(N__43446));
    LocalMux I__9660 (
            .O(N__43452),
            .I(data_cntvec_8));
    LocalMux I__9659 (
            .O(N__43449),
            .I(data_cntvec_8));
    Odrv4 I__9658 (
            .O(N__43446),
            .I(data_cntvec_8));
    CascadeMux I__9657 (
            .O(N__43439),
            .I(N__43435));
    InMux I__9656 (
            .O(N__43438),
            .I(N__43432));
    InMux I__9655 (
            .O(N__43435),
            .I(N__43429));
    LocalMux I__9654 (
            .O(N__43432),
            .I(data_cntvec_13));
    LocalMux I__9653 (
            .O(N__43429),
            .I(data_cntvec_13));
    CascadeMux I__9652 (
            .O(N__43424),
            .I(n14545_cascade_));
    CascadeMux I__9651 (
            .O(N__43421),
            .I(N__43417));
    InMux I__9650 (
            .O(N__43420),
            .I(N__43414));
    InMux I__9649 (
            .O(N__43417),
            .I(N__43411));
    LocalMux I__9648 (
            .O(N__43414),
            .I(N__43408));
    LocalMux I__9647 (
            .O(N__43411),
            .I(data_idxvec_1));
    Odrv12 I__9646 (
            .O(N__43408),
            .I(data_idxvec_1));
    CascadeMux I__9645 (
            .O(N__43403),
            .I(n26_adj_1522_cascade_));
    InMux I__9644 (
            .O(N__43400),
            .I(N__43397));
    LocalMux I__9643 (
            .O(N__43397),
            .I(N__43392));
    InMux I__9642 (
            .O(N__43396),
            .I(N__43389));
    InMux I__9641 (
            .O(N__43395),
            .I(N__43386));
    Span4Mux_h I__9640 (
            .O(N__43392),
            .I(N__43381));
    LocalMux I__9639 (
            .O(N__43389),
            .I(N__43381));
    LocalMux I__9638 (
            .O(N__43386),
            .I(acadc_skipCount_1));
    Odrv4 I__9637 (
            .O(N__43381),
            .I(acadc_skipCount_1));
    CascadeMux I__9636 (
            .O(N__43376),
            .I(n22190_cascade_));
    CascadeMux I__9635 (
            .O(N__43373),
            .I(n22193_cascade_));
    CascadeMux I__9634 (
            .O(N__43370),
            .I(n30_adj_1523_cascade_));
    InMux I__9633 (
            .O(N__43367),
            .I(N__43364));
    LocalMux I__9632 (
            .O(N__43364),
            .I(N__43361));
    Span4Mux_v I__9631 (
            .O(N__43361),
            .I(N__43358));
    Span4Mux_h I__9630 (
            .O(N__43358),
            .I(N__43355));
    Odrv4 I__9629 (
            .O(N__43355),
            .I(n19_adj_1520));
    CascadeMux I__9628 (
            .O(N__43352),
            .I(N__43349));
    InMux I__9627 (
            .O(N__43349),
            .I(N__43346));
    LocalMux I__9626 (
            .O(N__43346),
            .I(N__43343));
    Span4Mux_h I__9625 (
            .O(N__43343),
            .I(N__43340));
    Sp12to4 I__9624 (
            .O(N__43340),
            .I(N__43336));
    InMux I__9623 (
            .O(N__43339),
            .I(N__43333));
    Odrv12 I__9622 (
            .O(N__43336),
            .I(buf_readRTD_1));
    LocalMux I__9621 (
            .O(N__43333),
            .I(buf_readRTD_1));
    InMux I__9620 (
            .O(N__43328),
            .I(N__43325));
    LocalMux I__9619 (
            .O(N__43325),
            .I(N__43322));
    Span4Mux_h I__9618 (
            .O(N__43322),
            .I(N__43319));
    Odrv4 I__9617 (
            .O(N__43319),
            .I(comm_buf_5_2));
    InMux I__9616 (
            .O(N__43316),
            .I(N__43313));
    LocalMux I__9615 (
            .O(N__43313),
            .I(N__43310));
    Odrv4 I__9614 (
            .O(N__43310),
            .I(comm_buf_4_2));
    InMux I__9613 (
            .O(N__43307),
            .I(N__43304));
    LocalMux I__9612 (
            .O(N__43304),
            .I(N__43300));
    InMux I__9611 (
            .O(N__43303),
            .I(N__43297));
    Span4Mux_v I__9610 (
            .O(N__43300),
            .I(N__43294));
    LocalMux I__9609 (
            .O(N__43297),
            .I(N__43291));
    Span4Mux_h I__9608 (
            .O(N__43294),
            .I(N__43288));
    Odrv4 I__9607 (
            .O(N__43291),
            .I(comm_buf_6_2));
    Odrv4 I__9606 (
            .O(N__43288),
            .I(comm_buf_6_2));
    CascadeMux I__9605 (
            .O(N__43283),
            .I(n4_adj_1593_cascade_));
    InMux I__9604 (
            .O(N__43280),
            .I(N__43277));
    LocalMux I__9603 (
            .O(N__43277),
            .I(n22049));
    CascadeMux I__9602 (
            .O(N__43274),
            .I(n20801_cascade_));
    CascadeMux I__9601 (
            .O(N__43271),
            .I(N__43268));
    InMux I__9600 (
            .O(N__43268),
            .I(N__43265));
    LocalMux I__9599 (
            .O(N__43265),
            .I(N__43261));
    InMux I__9598 (
            .O(N__43264),
            .I(N__43258));
    Odrv4 I__9597 (
            .O(N__43261),
            .I(n20596));
    LocalMux I__9596 (
            .O(N__43258),
            .I(n20596));
    InMux I__9595 (
            .O(N__43253),
            .I(N__43250));
    LocalMux I__9594 (
            .O(N__43250),
            .I(N__43247));
    Span4Mux_v I__9593 (
            .O(N__43247),
            .I(N__43244));
    Odrv4 I__9592 (
            .O(N__43244),
            .I(n21094));
    CascadeMux I__9591 (
            .O(N__43241),
            .I(n21092_cascade_));
    InMux I__9590 (
            .O(N__43238),
            .I(N__43235));
    LocalMux I__9589 (
            .O(N__43235),
            .I(n20_adj_1610));
    InMux I__9588 (
            .O(N__43232),
            .I(N__43229));
    LocalMux I__9587 (
            .O(N__43229),
            .I(N__43226));
    Span4Mux_v I__9586 (
            .O(N__43226),
            .I(N__43223));
    Odrv4 I__9585 (
            .O(N__43223),
            .I(n20883));
    CascadeMux I__9584 (
            .O(N__43220),
            .I(n20695_cascade_));
    InMux I__9583 (
            .O(N__43217),
            .I(N__43214));
    LocalMux I__9582 (
            .O(N__43214),
            .I(N__43211));
    Span4Mux_v I__9581 (
            .O(N__43211),
            .I(N__43208));
    Odrv4 I__9580 (
            .O(N__43208),
            .I(n20881));
    InMux I__9579 (
            .O(N__43205),
            .I(N__43202));
    LocalMux I__9578 (
            .O(N__43202),
            .I(N__43198));
    InMux I__9577 (
            .O(N__43201),
            .I(N__43195));
    Span12Mux_v I__9576 (
            .O(N__43198),
            .I(N__43192));
    LocalMux I__9575 (
            .O(N__43195),
            .I(comm_buf_6_6));
    Odrv12 I__9574 (
            .O(N__43192),
            .I(comm_buf_6_6));
    CascadeMux I__9573 (
            .O(N__43187),
            .I(n21329_cascade_));
    CascadeMux I__9572 (
            .O(N__43184),
            .I(n21986_cascade_));
    InMux I__9571 (
            .O(N__43181),
            .I(N__43178));
    LocalMux I__9570 (
            .O(N__43178),
            .I(n2_adj_1584));
    CascadeMux I__9569 (
            .O(N__43175),
            .I(N__43172));
    InMux I__9568 (
            .O(N__43172),
            .I(N__43169));
    LocalMux I__9567 (
            .O(N__43169),
            .I(N__43165));
    InMux I__9566 (
            .O(N__43168),
            .I(N__43162));
    Span4Mux_v I__9565 (
            .O(N__43165),
            .I(N__43156));
    LocalMux I__9564 (
            .O(N__43162),
            .I(N__43156));
    InMux I__9563 (
            .O(N__43161),
            .I(N__43150));
    Span4Mux_v I__9562 (
            .O(N__43156),
            .I(N__43146));
    InMux I__9561 (
            .O(N__43155),
            .I(N__43143));
    InMux I__9560 (
            .O(N__43154),
            .I(N__43140));
    InMux I__9559 (
            .O(N__43153),
            .I(N__43137));
    LocalMux I__9558 (
            .O(N__43150),
            .I(N__43133));
    InMux I__9557 (
            .O(N__43149),
            .I(N__43130));
    Sp12to4 I__9556 (
            .O(N__43146),
            .I(N__43125));
    LocalMux I__9555 (
            .O(N__43143),
            .I(N__43125));
    LocalMux I__9554 (
            .O(N__43140),
            .I(N__43122));
    LocalMux I__9553 (
            .O(N__43137),
            .I(N__43119));
    InMux I__9552 (
            .O(N__43136),
            .I(N__43116));
    Span4Mux_v I__9551 (
            .O(N__43133),
            .I(N__43111));
    LocalMux I__9550 (
            .O(N__43130),
            .I(N__43111));
    Span12Mux_h I__9549 (
            .O(N__43125),
            .I(N__43108));
    Span4Mux_v I__9548 (
            .O(N__43122),
            .I(N__43103));
    Span4Mux_h I__9547 (
            .O(N__43119),
            .I(N__43103));
    LocalMux I__9546 (
            .O(N__43116),
            .I(N__43100));
    Span4Mux_v I__9545 (
            .O(N__43111),
            .I(N__43097));
    Span12Mux_v I__9544 (
            .O(N__43108),
            .I(N__43094));
    Span4Mux_v I__9543 (
            .O(N__43103),
            .I(N__43089));
    Span4Mux_h I__9542 (
            .O(N__43100),
            .I(N__43089));
    Span4Mux_h I__9541 (
            .O(N__43097),
            .I(N__43086));
    Odrv12 I__9540 (
            .O(N__43094),
            .I(comm_buf_0_6));
    Odrv4 I__9539 (
            .O(N__43089),
            .I(comm_buf_0_6));
    Odrv4 I__9538 (
            .O(N__43086),
            .I(comm_buf_0_6));
    InMux I__9537 (
            .O(N__43079),
            .I(N__43076));
    LocalMux I__9536 (
            .O(N__43076),
            .I(N__43073));
    Odrv4 I__9535 (
            .O(N__43073),
            .I(n1_adj_1583));
    CascadeMux I__9534 (
            .O(N__43070),
            .I(N__43067));
    InMux I__9533 (
            .O(N__43067),
            .I(N__43064));
    LocalMux I__9532 (
            .O(N__43064),
            .I(N__43060));
    InMux I__9531 (
            .O(N__43063),
            .I(N__43056));
    Span4Mux_v I__9530 (
            .O(N__43060),
            .I(N__43053));
    InMux I__9529 (
            .O(N__43059),
            .I(N__43050));
    LocalMux I__9528 (
            .O(N__43056),
            .I(n20621));
    Odrv4 I__9527 (
            .O(N__43053),
            .I(n20621));
    LocalMux I__9526 (
            .O(N__43050),
            .I(n20621));
    CascadeMux I__9525 (
            .O(N__43043),
            .I(n7_cascade_));
    InMux I__9524 (
            .O(N__43040),
            .I(N__43037));
    LocalMux I__9523 (
            .O(N__43037),
            .I(N__43034));
    Span4Mux_v I__9522 (
            .O(N__43034),
            .I(N__43031));
    Span4Mux_h I__9521 (
            .O(N__43031),
            .I(N__43028));
    Odrv4 I__9520 (
            .O(N__43028),
            .I(comm_buf_2_2));
    CascadeMux I__9519 (
            .O(N__43025),
            .I(N__43022));
    InMux I__9518 (
            .O(N__43022),
            .I(N__43019));
    LocalMux I__9517 (
            .O(N__43019),
            .I(N__43016));
    Span4Mux_h I__9516 (
            .O(N__43016),
            .I(N__43013));
    Odrv4 I__9515 (
            .O(N__43013),
            .I(comm_buf_3_2));
    CascadeMux I__9514 (
            .O(N__43010),
            .I(N__43006));
    InMux I__9513 (
            .O(N__43009),
            .I(N__43000));
    InMux I__9512 (
            .O(N__43006),
            .I(N__42997));
    CascadeMux I__9511 (
            .O(N__43005),
            .I(N__42994));
    CascadeMux I__9510 (
            .O(N__43004),
            .I(N__42991));
    CascadeMux I__9509 (
            .O(N__43003),
            .I(N__42988));
    LocalMux I__9508 (
            .O(N__43000),
            .I(N__42982));
    LocalMux I__9507 (
            .O(N__42997),
            .I(N__42982));
    InMux I__9506 (
            .O(N__42994),
            .I(N__42979));
    InMux I__9505 (
            .O(N__42991),
            .I(N__42976));
    InMux I__9504 (
            .O(N__42988),
            .I(N__42973));
    InMux I__9503 (
            .O(N__42987),
            .I(N__42967));
    Span4Mux_v I__9502 (
            .O(N__42982),
            .I(N__42962));
    LocalMux I__9501 (
            .O(N__42979),
            .I(N__42962));
    LocalMux I__9500 (
            .O(N__42976),
            .I(N__42959));
    LocalMux I__9499 (
            .O(N__42973),
            .I(N__42956));
    InMux I__9498 (
            .O(N__42972),
            .I(N__42953));
    InMux I__9497 (
            .O(N__42971),
            .I(N__42950));
    InMux I__9496 (
            .O(N__42970),
            .I(N__42947));
    LocalMux I__9495 (
            .O(N__42967),
            .I(N__42944));
    Span4Mux_v I__9494 (
            .O(N__42962),
            .I(N__42941));
    Span4Mux_h I__9493 (
            .O(N__42959),
            .I(N__42936));
    Span4Mux_v I__9492 (
            .O(N__42956),
            .I(N__42936));
    LocalMux I__9491 (
            .O(N__42953),
            .I(N__42933));
    LocalMux I__9490 (
            .O(N__42950),
            .I(N__42930));
    LocalMux I__9489 (
            .O(N__42947),
            .I(N__42923));
    Span4Mux_v I__9488 (
            .O(N__42944),
            .I(N__42923));
    Span4Mux_h I__9487 (
            .O(N__42941),
            .I(N__42923));
    Span4Mux_v I__9486 (
            .O(N__42936),
            .I(N__42920));
    Span4Mux_h I__9485 (
            .O(N__42933),
            .I(N__42917));
    Span4Mux_h I__9484 (
            .O(N__42930),
            .I(N__42914));
    Sp12to4 I__9483 (
            .O(N__42923),
            .I(N__42911));
    Span4Mux_h I__9482 (
            .O(N__42920),
            .I(N__42906));
    Span4Mux_h I__9481 (
            .O(N__42917),
            .I(N__42906));
    Span4Mux_h I__9480 (
            .O(N__42914),
            .I(N__42903));
    Odrv12 I__9479 (
            .O(N__42911),
            .I(comm_buf_0_2));
    Odrv4 I__9478 (
            .O(N__42906),
            .I(comm_buf_0_2));
    Odrv4 I__9477 (
            .O(N__42903),
            .I(comm_buf_0_2));
    CascadeMux I__9476 (
            .O(N__42896),
            .I(n22046_cascade_));
    InMux I__9475 (
            .O(N__42893),
            .I(N__42890));
    LocalMux I__9474 (
            .O(N__42890),
            .I(N__42887));
    Span4Mux_h I__9473 (
            .O(N__42887),
            .I(N__42884));
    Span4Mux_v I__9472 (
            .O(N__42884),
            .I(N__42881));
    Odrv4 I__9471 (
            .O(N__42881),
            .I(n30_adj_1529));
    InMux I__9470 (
            .O(N__42878),
            .I(N__42875));
    LocalMux I__9469 (
            .O(N__42875),
            .I(N__42872));
    Span4Mux_h I__9468 (
            .O(N__42872),
            .I(N__42869));
    Span4Mux_v I__9467 (
            .O(N__42869),
            .I(N__42866));
    Span4Mux_v I__9466 (
            .O(N__42866),
            .I(N__42863));
    Span4Mux_h I__9465 (
            .O(N__42863),
            .I(N__42860));
    Odrv4 I__9464 (
            .O(N__42860),
            .I(n22109));
    SRMux I__9463 (
            .O(N__42857),
            .I(N__42853));
    SRMux I__9462 (
            .O(N__42856),
            .I(N__42848));
    LocalMux I__9461 (
            .O(N__42853),
            .I(N__42844));
    SRMux I__9460 (
            .O(N__42852),
            .I(N__42841));
    SRMux I__9459 (
            .O(N__42851),
            .I(N__42838));
    LocalMux I__9458 (
            .O(N__42848),
            .I(N__42835));
    SRMux I__9457 (
            .O(N__42847),
            .I(N__42832));
    Span4Mux_v I__9456 (
            .O(N__42844),
            .I(N__42826));
    LocalMux I__9455 (
            .O(N__42841),
            .I(N__42826));
    LocalMux I__9454 (
            .O(N__42838),
            .I(N__42823));
    Span4Mux_h I__9453 (
            .O(N__42835),
            .I(N__42820));
    LocalMux I__9452 (
            .O(N__42832),
            .I(N__42817));
    SRMux I__9451 (
            .O(N__42831),
            .I(N__42814));
    Span4Mux_h I__9450 (
            .O(N__42826),
            .I(N__42811));
    Span4Mux_h I__9449 (
            .O(N__42823),
            .I(N__42808));
    Span4Mux_v I__9448 (
            .O(N__42820),
            .I(N__42803));
    Span4Mux_v I__9447 (
            .O(N__42817),
            .I(N__42803));
    LocalMux I__9446 (
            .O(N__42814),
            .I(N__42800));
    Odrv4 I__9445 (
            .O(N__42811),
            .I(n14766));
    Odrv4 I__9444 (
            .O(N__42808),
            .I(n14766));
    Odrv4 I__9443 (
            .O(N__42803),
            .I(n14766));
    Odrv12 I__9442 (
            .O(N__42800),
            .I(n14766));
    CascadeMux I__9441 (
            .O(N__42791),
            .I(n21199_cascade_));
    CascadeMux I__9440 (
            .O(N__42788),
            .I(n20681_cascade_));
    InMux I__9439 (
            .O(N__42785),
            .I(N__42779));
    InMux I__9438 (
            .O(N__42784),
            .I(N__42773));
    InMux I__9437 (
            .O(N__42783),
            .I(N__42773));
    InMux I__9436 (
            .O(N__42782),
            .I(N__42770));
    LocalMux I__9435 (
            .O(N__42779),
            .I(N__42767));
    InMux I__9434 (
            .O(N__42778),
            .I(N__42764));
    LocalMux I__9433 (
            .O(N__42773),
            .I(N__42761));
    LocalMux I__9432 (
            .O(N__42770),
            .I(N__42758));
    Span4Mux_v I__9431 (
            .O(N__42767),
            .I(N__42755));
    LocalMux I__9430 (
            .O(N__42764),
            .I(N__42752));
    Span4Mux_h I__9429 (
            .O(N__42761),
            .I(N__42749));
    Span4Mux_h I__9428 (
            .O(N__42758),
            .I(N__42746));
    Span4Mux_h I__9427 (
            .O(N__42755),
            .I(N__42741));
    Span4Mux_h I__9426 (
            .O(N__42752),
            .I(N__42741));
    Odrv4 I__9425 (
            .O(N__42749),
            .I(n20599));
    Odrv4 I__9424 (
            .O(N__42746),
            .I(n20599));
    Odrv4 I__9423 (
            .O(N__42741),
            .I(n20599));
    CascadeMux I__9422 (
            .O(N__42734),
            .I(n12108_cascade_));
    InMux I__9421 (
            .O(N__42731),
            .I(N__42728));
    LocalMux I__9420 (
            .O(N__42728),
            .I(n4_adj_1616));
    CEMux I__9419 (
            .O(N__42725),
            .I(N__42718));
    CEMux I__9418 (
            .O(N__42724),
            .I(N__42714));
    CEMux I__9417 (
            .O(N__42723),
            .I(N__42711));
    CEMux I__9416 (
            .O(N__42722),
            .I(N__42708));
    CEMux I__9415 (
            .O(N__42721),
            .I(N__42705));
    LocalMux I__9414 (
            .O(N__42718),
            .I(N__42702));
    CEMux I__9413 (
            .O(N__42717),
            .I(N__42699));
    LocalMux I__9412 (
            .O(N__42714),
            .I(N__42696));
    LocalMux I__9411 (
            .O(N__42711),
            .I(N__42693));
    LocalMux I__9410 (
            .O(N__42708),
            .I(N__42690));
    LocalMux I__9409 (
            .O(N__42705),
            .I(N__42686));
    Span12Mux_v I__9408 (
            .O(N__42702),
            .I(N__42683));
    LocalMux I__9407 (
            .O(N__42699),
            .I(N__42676));
    Span4Mux_v I__9406 (
            .O(N__42696),
            .I(N__42676));
    Span4Mux_v I__9405 (
            .O(N__42693),
            .I(N__42676));
    Sp12to4 I__9404 (
            .O(N__42690),
            .I(N__42673));
    InMux I__9403 (
            .O(N__42689),
            .I(N__42670));
    Odrv4 I__9402 (
            .O(N__42686),
            .I(n11977));
    Odrv12 I__9401 (
            .O(N__42683),
            .I(n11977));
    Odrv4 I__9400 (
            .O(N__42676),
            .I(n11977));
    Odrv12 I__9399 (
            .O(N__42673),
            .I(n11977));
    LocalMux I__9398 (
            .O(N__42670),
            .I(n11977));
    InMux I__9397 (
            .O(N__42659),
            .I(N__42656));
    LocalMux I__9396 (
            .O(N__42656),
            .I(N__42653));
    Span4Mux_h I__9395 (
            .O(N__42653),
            .I(N__42650));
    Odrv4 I__9394 (
            .O(N__42650),
            .I(comm_buf_3_6));
    InMux I__9393 (
            .O(N__42647),
            .I(N__42644));
    LocalMux I__9392 (
            .O(N__42644),
            .I(N__42641));
    Odrv12 I__9391 (
            .O(N__42641),
            .I(comm_buf_2_6));
    InMux I__9390 (
            .O(N__42638),
            .I(N__42635));
    LocalMux I__9389 (
            .O(N__42635),
            .I(N__42632));
    Odrv12 I__9388 (
            .O(N__42632),
            .I(buf_data_iac_22));
    InMux I__9387 (
            .O(N__42629),
            .I(N__42626));
    LocalMux I__9386 (
            .O(N__42626),
            .I(N__42623));
    Span4Mux_v I__9385 (
            .O(N__42623),
            .I(N__42620));
    Odrv4 I__9384 (
            .O(N__42620),
            .I(n21038));
    InMux I__9383 (
            .O(N__42617),
            .I(N__42614));
    LocalMux I__9382 (
            .O(N__42614),
            .I(N__42611));
    Span4Mux_v I__9381 (
            .O(N__42611),
            .I(N__42600));
    InMux I__9380 (
            .O(N__42610),
            .I(N__42597));
    InMux I__9379 (
            .O(N__42609),
            .I(N__42582));
    InMux I__9378 (
            .O(N__42608),
            .I(N__42582));
    InMux I__9377 (
            .O(N__42607),
            .I(N__42582));
    InMux I__9376 (
            .O(N__42606),
            .I(N__42582));
    InMux I__9375 (
            .O(N__42605),
            .I(N__42582));
    InMux I__9374 (
            .O(N__42604),
            .I(N__42582));
    InMux I__9373 (
            .O(N__42603),
            .I(N__42582));
    Odrv4 I__9372 (
            .O(N__42600),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__9371 (
            .O(N__42597),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__9370 (
            .O(N__42582),
            .I(\comm_spi.bit_cnt_3 ));
    InMux I__9369 (
            .O(N__42575),
            .I(N__42568));
    InMux I__9368 (
            .O(N__42574),
            .I(N__42568));
    InMux I__9367 (
            .O(N__42573),
            .I(N__42565));
    LocalMux I__9366 (
            .O(N__42568),
            .I(\comm_spi.bit_cnt_2 ));
    LocalMux I__9365 (
            .O(N__42565),
            .I(\comm_spi.bit_cnt_2 ));
    InMux I__9364 (
            .O(N__42560),
            .I(N__42550));
    InMux I__9363 (
            .O(N__42559),
            .I(N__42550));
    InMux I__9362 (
            .O(N__42558),
            .I(N__42550));
    InMux I__9361 (
            .O(N__42557),
            .I(N__42547));
    LocalMux I__9360 (
            .O(N__42550),
            .I(\comm_spi.bit_cnt_1 ));
    LocalMux I__9359 (
            .O(N__42547),
            .I(\comm_spi.bit_cnt_1 ));
    CascadeMux I__9358 (
            .O(N__42542),
            .I(N__42539));
    InMux I__9357 (
            .O(N__42539),
            .I(N__42526));
    InMux I__9356 (
            .O(N__42538),
            .I(N__42526));
    InMux I__9355 (
            .O(N__42537),
            .I(N__42526));
    InMux I__9354 (
            .O(N__42536),
            .I(N__42526));
    InMux I__9353 (
            .O(N__42535),
            .I(N__42523));
    LocalMux I__9352 (
            .O(N__42526),
            .I(\comm_spi.bit_cnt_0 ));
    LocalMux I__9351 (
            .O(N__42523),
            .I(\comm_spi.bit_cnt_0 ));
    InMux I__9350 (
            .O(N__42518),
            .I(n19507));
    InMux I__9349 (
            .O(N__42515),
            .I(n19508));
    InMux I__9348 (
            .O(N__42512),
            .I(N__42508));
    InMux I__9347 (
            .O(N__42511),
            .I(N__42505));
    LocalMux I__9346 (
            .O(N__42508),
            .I(clk_cnt_0));
    LocalMux I__9345 (
            .O(N__42505),
            .I(clk_cnt_0));
    InMux I__9344 (
            .O(N__42500),
            .I(N__42496));
    InMux I__9343 (
            .O(N__42499),
            .I(N__42493));
    LocalMux I__9342 (
            .O(N__42496),
            .I(clk_cnt_4));
    LocalMux I__9341 (
            .O(N__42493),
            .I(clk_cnt_4));
    InMux I__9340 (
            .O(N__42488),
            .I(N__42484));
    InMux I__9339 (
            .O(N__42487),
            .I(N__42481));
    LocalMux I__9338 (
            .O(N__42484),
            .I(N__42478));
    LocalMux I__9337 (
            .O(N__42481),
            .I(clk_cnt_1));
    Odrv4 I__9336 (
            .O(N__42478),
            .I(clk_cnt_1));
    InMux I__9335 (
            .O(N__42473),
            .I(N__42469));
    InMux I__9334 (
            .O(N__42472),
            .I(N__42466));
    LocalMux I__9333 (
            .O(N__42469),
            .I(clk_cnt_3));
    LocalMux I__9332 (
            .O(N__42466),
            .I(clk_cnt_3));
    CascadeMux I__9331 (
            .O(N__42461),
            .I(n6_cascade_));
    InMux I__9330 (
            .O(N__42458),
            .I(N__42454));
    InMux I__9329 (
            .O(N__42457),
            .I(N__42451));
    LocalMux I__9328 (
            .O(N__42454),
            .I(N__42448));
    LocalMux I__9327 (
            .O(N__42451),
            .I(clk_cnt_2));
    Odrv4 I__9326 (
            .O(N__42448),
            .I(clk_cnt_2));
    InMux I__9325 (
            .O(N__42443),
            .I(N__42440));
    LocalMux I__9324 (
            .O(N__42440),
            .I(N__42435));
    CascadeMux I__9323 (
            .O(N__42439),
            .I(N__42432));
    CascadeMux I__9322 (
            .O(N__42438),
            .I(N__42429));
    Span4Mux_h I__9321 (
            .O(N__42435),
            .I(N__42426));
    InMux I__9320 (
            .O(N__42432),
            .I(N__42421));
    InMux I__9319 (
            .O(N__42429),
            .I(N__42421));
    Odrv4 I__9318 (
            .O(N__42426),
            .I(acadc_skipCount_11));
    LocalMux I__9317 (
            .O(N__42421),
            .I(acadc_skipCount_11));
    InMux I__9316 (
            .O(N__42416),
            .I(N__42412));
    InMux I__9315 (
            .O(N__42415),
            .I(N__42409));
    LocalMux I__9314 (
            .O(N__42412),
            .I(dds0_mclkcnt_3));
    LocalMux I__9313 (
            .O(N__42409),
            .I(dds0_mclkcnt_3));
    InMux I__9312 (
            .O(N__42404),
            .I(N__42400));
    InMux I__9311 (
            .O(N__42403),
            .I(N__42397));
    LocalMux I__9310 (
            .O(N__42400),
            .I(dds0_mclkcnt_5));
    LocalMux I__9309 (
            .O(N__42397),
            .I(dds0_mclkcnt_5));
    CascadeMux I__9308 (
            .O(N__42392),
            .I(N__42388));
    InMux I__9307 (
            .O(N__42391),
            .I(N__42385));
    InMux I__9306 (
            .O(N__42388),
            .I(N__42382));
    LocalMux I__9305 (
            .O(N__42385),
            .I(dds0_mclkcnt_1));
    LocalMux I__9304 (
            .O(N__42382),
            .I(dds0_mclkcnt_1));
    InMux I__9303 (
            .O(N__42377),
            .I(N__42373));
    InMux I__9302 (
            .O(N__42376),
            .I(N__42370));
    LocalMux I__9301 (
            .O(N__42373),
            .I(dds0_mclkcnt_4));
    LocalMux I__9300 (
            .O(N__42370),
            .I(dds0_mclkcnt_4));
    InMux I__9299 (
            .O(N__42365),
            .I(N__42361));
    InMux I__9298 (
            .O(N__42364),
            .I(N__42358));
    LocalMux I__9297 (
            .O(N__42361),
            .I(dds0_mclkcnt_2));
    LocalMux I__9296 (
            .O(N__42358),
            .I(dds0_mclkcnt_2));
    InMux I__9295 (
            .O(N__42353),
            .I(N__42349));
    InMux I__9294 (
            .O(N__42352),
            .I(N__42346));
    LocalMux I__9293 (
            .O(N__42349),
            .I(dds0_mclkcnt_0));
    LocalMux I__9292 (
            .O(N__42346),
            .I(dds0_mclkcnt_0));
    CascadeMux I__9291 (
            .O(N__42341),
            .I(n12_cascade_));
    InMux I__9290 (
            .O(N__42338),
            .I(N__42334));
    InMux I__9289 (
            .O(N__42337),
            .I(N__42331));
    LocalMux I__9288 (
            .O(N__42334),
            .I(dds0_mclkcnt_7));
    LocalMux I__9287 (
            .O(N__42331),
            .I(dds0_mclkcnt_7));
    InMux I__9286 (
            .O(N__42326),
            .I(N__42323));
    LocalMux I__9285 (
            .O(N__42323),
            .I(n20543));
    CascadeMux I__9284 (
            .O(N__42320),
            .I(n20543_cascade_));
    InMux I__9283 (
            .O(N__42317),
            .I(N__42313));
    InMux I__9282 (
            .O(N__42316),
            .I(N__42310));
    LocalMux I__9281 (
            .O(N__42313),
            .I(dds0_mclkcnt_6));
    LocalMux I__9280 (
            .O(N__42310),
            .I(dds0_mclkcnt_6));
    CascadeMux I__9279 (
            .O(N__42305),
            .I(n8_adj_1559_cascade_));
    CascadeMux I__9278 (
            .O(N__42302),
            .I(N__42299));
    CascadeBuf I__9277 (
            .O(N__42299),
            .I(N__42296));
    CascadeMux I__9276 (
            .O(N__42296),
            .I(N__42293));
    CascadeBuf I__9275 (
            .O(N__42293),
            .I(N__42290));
    CascadeMux I__9274 (
            .O(N__42290),
            .I(N__42287));
    CascadeBuf I__9273 (
            .O(N__42287),
            .I(N__42284));
    CascadeMux I__9272 (
            .O(N__42284),
            .I(N__42281));
    CascadeBuf I__9271 (
            .O(N__42281),
            .I(N__42278));
    CascadeMux I__9270 (
            .O(N__42278),
            .I(N__42275));
    CascadeBuf I__9269 (
            .O(N__42275),
            .I(N__42272));
    CascadeMux I__9268 (
            .O(N__42272),
            .I(N__42269));
    CascadeBuf I__9267 (
            .O(N__42269),
            .I(N__42266));
    CascadeMux I__9266 (
            .O(N__42266),
            .I(N__42263));
    CascadeBuf I__9265 (
            .O(N__42263),
            .I(N__42260));
    CascadeMux I__9264 (
            .O(N__42260),
            .I(N__42256));
    CascadeMux I__9263 (
            .O(N__42259),
            .I(N__42253));
    CascadeBuf I__9262 (
            .O(N__42256),
            .I(N__42250));
    CascadeBuf I__9261 (
            .O(N__42253),
            .I(N__42247));
    CascadeMux I__9260 (
            .O(N__42250),
            .I(N__42244));
    CascadeMux I__9259 (
            .O(N__42247),
            .I(N__42241));
    CascadeBuf I__9258 (
            .O(N__42244),
            .I(N__42238));
    InMux I__9257 (
            .O(N__42241),
            .I(N__42235));
    CascadeMux I__9256 (
            .O(N__42238),
            .I(N__42232));
    LocalMux I__9255 (
            .O(N__42235),
            .I(N__42229));
    InMux I__9254 (
            .O(N__42232),
            .I(N__42226));
    Span12Mux_h I__9253 (
            .O(N__42229),
            .I(N__42223));
    LocalMux I__9252 (
            .O(N__42226),
            .I(N__42220));
    Span12Mux_v I__9251 (
            .O(N__42223),
            .I(N__42215));
    Span12Mux_s11_v I__9250 (
            .O(N__42220),
            .I(N__42215));
    Odrv12 I__9249 (
            .O(N__42215),
            .I(data_index_9_N_216_6));
    InMux I__9248 (
            .O(N__42212),
            .I(N__42209));
    LocalMux I__9247 (
            .O(N__42209),
            .I(N__42206));
    Span4Mux_v I__9246 (
            .O(N__42206),
            .I(N__42203));
    Odrv4 I__9245 (
            .O(N__42203),
            .I(n8_adj_1567));
    InMux I__9244 (
            .O(N__42200),
            .I(N__42196));
    InMux I__9243 (
            .O(N__42199),
            .I(N__42193));
    LocalMux I__9242 (
            .O(N__42196),
            .I(N__42190));
    LocalMux I__9241 (
            .O(N__42193),
            .I(N__42187));
    Span4Mux_v I__9240 (
            .O(N__42190),
            .I(N__42182));
    Span4Mux_h I__9239 (
            .O(N__42187),
            .I(N__42182));
    Span4Mux_h I__9238 (
            .O(N__42182),
            .I(N__42179));
    Odrv4 I__9237 (
            .O(N__42179),
            .I(n7_adj_1566));
    CascadeMux I__9236 (
            .O(N__42176),
            .I(N__42173));
    CascadeBuf I__9235 (
            .O(N__42173),
            .I(N__42170));
    CascadeMux I__9234 (
            .O(N__42170),
            .I(N__42167));
    CascadeBuf I__9233 (
            .O(N__42167),
            .I(N__42164));
    CascadeMux I__9232 (
            .O(N__42164),
            .I(N__42161));
    CascadeBuf I__9231 (
            .O(N__42161),
            .I(N__42158));
    CascadeMux I__9230 (
            .O(N__42158),
            .I(N__42155));
    CascadeBuf I__9229 (
            .O(N__42155),
            .I(N__42152));
    CascadeMux I__9228 (
            .O(N__42152),
            .I(N__42149));
    CascadeBuf I__9227 (
            .O(N__42149),
            .I(N__42146));
    CascadeMux I__9226 (
            .O(N__42146),
            .I(N__42143));
    CascadeBuf I__9225 (
            .O(N__42143),
            .I(N__42140));
    CascadeMux I__9224 (
            .O(N__42140),
            .I(N__42137));
    CascadeBuf I__9223 (
            .O(N__42137),
            .I(N__42134));
    CascadeMux I__9222 (
            .O(N__42134),
            .I(N__42131));
    CascadeBuf I__9221 (
            .O(N__42131),
            .I(N__42127));
    CascadeMux I__9220 (
            .O(N__42130),
            .I(N__42124));
    CascadeMux I__9219 (
            .O(N__42127),
            .I(N__42121));
    CascadeBuf I__9218 (
            .O(N__42124),
            .I(N__42118));
    CascadeBuf I__9217 (
            .O(N__42121),
            .I(N__42115));
    CascadeMux I__9216 (
            .O(N__42118),
            .I(N__42112));
    CascadeMux I__9215 (
            .O(N__42115),
            .I(N__42109));
    InMux I__9214 (
            .O(N__42112),
            .I(N__42106));
    InMux I__9213 (
            .O(N__42109),
            .I(N__42103));
    LocalMux I__9212 (
            .O(N__42106),
            .I(N__42100));
    LocalMux I__9211 (
            .O(N__42103),
            .I(N__42097));
    Span12Mux_s11_h I__9210 (
            .O(N__42100),
            .I(N__42094));
    Span4Mux_h I__9209 (
            .O(N__42097),
            .I(N__42091));
    Span12Mux_v I__9208 (
            .O(N__42094),
            .I(N__42088));
    Span4Mux_v I__9207 (
            .O(N__42091),
            .I(N__42085));
    Odrv12 I__9206 (
            .O(N__42088),
            .I(data_index_9_N_216_1));
    Odrv4 I__9205 (
            .O(N__42085),
            .I(data_index_9_N_216_1));
    InMux I__9204 (
            .O(N__42080),
            .I(N__42076));
    InMux I__9203 (
            .O(N__42079),
            .I(N__42073));
    LocalMux I__9202 (
            .O(N__42076),
            .I(data_cntvec_12));
    LocalMux I__9201 (
            .O(N__42073),
            .I(data_cntvec_12));
    InMux I__9200 (
            .O(N__42068),
            .I(N__42065));
    LocalMux I__9199 (
            .O(N__42065),
            .I(N__42062));
    Span4Mux_h I__9198 (
            .O(N__42062),
            .I(N__42057));
    InMux I__9197 (
            .O(N__42061),
            .I(N__42054));
    InMux I__9196 (
            .O(N__42060),
            .I(N__42051));
    Span4Mux_v I__9195 (
            .O(N__42057),
            .I(N__42048));
    LocalMux I__9194 (
            .O(N__42054),
            .I(data_cntvec_10));
    LocalMux I__9193 (
            .O(N__42051),
            .I(data_cntvec_10));
    Odrv4 I__9192 (
            .O(N__42048),
            .I(data_cntvec_10));
    InMux I__9191 (
            .O(N__42041),
            .I(N__42036));
    CascadeMux I__9190 (
            .O(N__42040),
            .I(N__42033));
    InMux I__9189 (
            .O(N__42039),
            .I(N__42030));
    LocalMux I__9188 (
            .O(N__42036),
            .I(N__42027));
    InMux I__9187 (
            .O(N__42033),
            .I(N__42024));
    LocalMux I__9186 (
            .O(N__42030),
            .I(req_data_cnt_12));
    Odrv4 I__9185 (
            .O(N__42027),
            .I(req_data_cnt_12));
    LocalMux I__9184 (
            .O(N__42024),
            .I(req_data_cnt_12));
    InMux I__9183 (
            .O(N__42017),
            .I(N__42014));
    LocalMux I__9182 (
            .O(N__42014),
            .I(N__42010));
    InMux I__9181 (
            .O(N__42013),
            .I(N__42006));
    Span4Mux_v I__9180 (
            .O(N__42010),
            .I(N__42003));
    InMux I__9179 (
            .O(N__42009),
            .I(N__42000));
    LocalMux I__9178 (
            .O(N__42006),
            .I(req_data_cnt_10));
    Odrv4 I__9177 (
            .O(N__42003),
            .I(req_data_cnt_10));
    LocalMux I__9176 (
            .O(N__42000),
            .I(req_data_cnt_10));
    InMux I__9175 (
            .O(N__41993),
            .I(N__41990));
    LocalMux I__9174 (
            .O(N__41990),
            .I(n8_adj_1559));
    CascadeMux I__9173 (
            .O(N__41987),
            .I(N__41984));
    InMux I__9172 (
            .O(N__41984),
            .I(N__41978));
    InMux I__9171 (
            .O(N__41983),
            .I(N__41978));
    LocalMux I__9170 (
            .O(N__41978),
            .I(N__41975));
    Span4Mux_v I__9169 (
            .O(N__41975),
            .I(N__41972));
    Span4Mux_v I__9168 (
            .O(N__41972),
            .I(N__41969));
    Span4Mux_h I__9167 (
            .O(N__41969),
            .I(N__41966));
    Odrv4 I__9166 (
            .O(N__41966),
            .I(n7_adj_1558));
    InMux I__9165 (
            .O(N__41963),
            .I(N__41959));
    InMux I__9164 (
            .O(N__41962),
            .I(N__41956));
    LocalMux I__9163 (
            .O(N__41959),
            .I(N__41953));
    LocalMux I__9162 (
            .O(N__41956),
            .I(N__41950));
    Span4Mux_h I__9161 (
            .O(N__41953),
            .I(N__41946));
    Span4Mux_h I__9160 (
            .O(N__41950),
            .I(N__41943));
    InMux I__9159 (
            .O(N__41949),
            .I(N__41940));
    Span4Mux_h I__9158 (
            .O(N__41946),
            .I(N__41935));
    Span4Mux_h I__9157 (
            .O(N__41943),
            .I(N__41935));
    LocalMux I__9156 (
            .O(N__41940),
            .I(data_index_6));
    Odrv4 I__9155 (
            .O(N__41935),
            .I(data_index_6));
    SRMux I__9154 (
            .O(N__41930),
            .I(N__41927));
    LocalMux I__9153 (
            .O(N__41927),
            .I(N__41924));
    Span4Mux_h I__9152 (
            .O(N__41924),
            .I(N__41921));
    Span4Mux_v I__9151 (
            .O(N__41921),
            .I(N__41918));
    Odrv4 I__9150 (
            .O(N__41918),
            .I(\comm_spi.data_tx_7__N_771 ));
    InMux I__9149 (
            .O(N__41915),
            .I(bfn_15_16_0_));
    InMux I__9148 (
            .O(N__41912),
            .I(n19505));
    InMux I__9147 (
            .O(N__41909),
            .I(n19506));
    InMux I__9146 (
            .O(N__41906),
            .I(n19363));
    InMux I__9145 (
            .O(N__41903),
            .I(n19364));
    InMux I__9144 (
            .O(N__41900),
            .I(n19365));
    InMux I__9143 (
            .O(N__41897),
            .I(n19366));
    InMux I__9142 (
            .O(N__41894),
            .I(n19367));
    InMux I__9141 (
            .O(N__41891),
            .I(n19368));
    CEMux I__9140 (
            .O(N__41888),
            .I(N__41882));
    CEMux I__9139 (
            .O(N__41887),
            .I(N__41879));
    CEMux I__9138 (
            .O(N__41886),
            .I(N__41876));
    InMux I__9137 (
            .O(N__41885),
            .I(N__41872));
    LocalMux I__9136 (
            .O(N__41882),
            .I(N__41869));
    LocalMux I__9135 (
            .O(N__41879),
            .I(N__41866));
    LocalMux I__9134 (
            .O(N__41876),
            .I(N__41863));
    CEMux I__9133 (
            .O(N__41875),
            .I(N__41860));
    LocalMux I__9132 (
            .O(N__41872),
            .I(N__41857));
    Span4Mux_v I__9131 (
            .O(N__41869),
            .I(N__41848));
    Span4Mux_v I__9130 (
            .O(N__41866),
            .I(N__41848));
    Span4Mux_v I__9129 (
            .O(N__41863),
            .I(N__41848));
    LocalMux I__9128 (
            .O(N__41860),
            .I(N__41848));
    Span4Mux_h I__9127 (
            .O(N__41857),
            .I(N__41845));
    Odrv4 I__9126 (
            .O(N__41848),
            .I(n13473));
    Odrv4 I__9125 (
            .O(N__41845),
            .I(n13473));
    SRMux I__9124 (
            .O(N__41840),
            .I(N__41836));
    SRMux I__9123 (
            .O(N__41839),
            .I(N__41833));
    LocalMux I__9122 (
            .O(N__41836),
            .I(N__41829));
    LocalMux I__9121 (
            .O(N__41833),
            .I(N__41825));
    SRMux I__9120 (
            .O(N__41832),
            .I(N__41822));
    Span4Mux_h I__9119 (
            .O(N__41829),
            .I(N__41819));
    SRMux I__9118 (
            .O(N__41828),
            .I(N__41816));
    Span4Mux_v I__9117 (
            .O(N__41825),
            .I(N__41811));
    LocalMux I__9116 (
            .O(N__41822),
            .I(N__41811));
    Sp12to4 I__9115 (
            .O(N__41819),
            .I(N__41806));
    LocalMux I__9114 (
            .O(N__41816),
            .I(N__41806));
    Span4Mux_h I__9113 (
            .O(N__41811),
            .I(N__41803));
    Odrv12 I__9112 (
            .O(N__41806),
            .I(n14663));
    Odrv4 I__9111 (
            .O(N__41803),
            .I(n14663));
    InMux I__9110 (
            .O(N__41798),
            .I(N__41794));
    InMux I__9109 (
            .O(N__41797),
            .I(N__41791));
    LocalMux I__9108 (
            .O(N__41794),
            .I(data_cntvec_14));
    LocalMux I__9107 (
            .O(N__41791),
            .I(data_cntvec_14));
    InMux I__9106 (
            .O(N__41786),
            .I(N__41781));
    InMux I__9105 (
            .O(N__41785),
            .I(N__41778));
    InMux I__9104 (
            .O(N__41784),
            .I(N__41775));
    LocalMux I__9103 (
            .O(N__41781),
            .I(N__41772));
    LocalMux I__9102 (
            .O(N__41778),
            .I(data_cntvec_11));
    LocalMux I__9101 (
            .O(N__41775),
            .I(data_cntvec_11));
    Odrv12 I__9100 (
            .O(N__41772),
            .I(data_cntvec_11));
    InMux I__9099 (
            .O(N__41765),
            .I(N__41758));
    InMux I__9098 (
            .O(N__41764),
            .I(N__41758));
    InMux I__9097 (
            .O(N__41763),
            .I(N__41755));
    LocalMux I__9096 (
            .O(N__41758),
            .I(req_data_cnt_14));
    LocalMux I__9095 (
            .O(N__41755),
            .I(req_data_cnt_14));
    InMux I__9094 (
            .O(N__41750),
            .I(N__41743));
    InMux I__9093 (
            .O(N__41749),
            .I(N__41740));
    InMux I__9092 (
            .O(N__41748),
            .I(N__41737));
    InMux I__9091 (
            .O(N__41747),
            .I(N__41734));
    InMux I__9090 (
            .O(N__41746),
            .I(N__41731));
    LocalMux I__9089 (
            .O(N__41743),
            .I(N__41725));
    LocalMux I__9088 (
            .O(N__41740),
            .I(N__41722));
    LocalMux I__9087 (
            .O(N__41737),
            .I(N__41715));
    LocalMux I__9086 (
            .O(N__41734),
            .I(N__41715));
    LocalMux I__9085 (
            .O(N__41731),
            .I(N__41715));
    InMux I__9084 (
            .O(N__41730),
            .I(N__41710));
    InMux I__9083 (
            .O(N__41729),
            .I(N__41710));
    InMux I__9082 (
            .O(N__41728),
            .I(N__41705));
    Span4Mux_h I__9081 (
            .O(N__41725),
            .I(N__41696));
    Span4Mux_h I__9080 (
            .O(N__41722),
            .I(N__41696));
    Span4Mux_v I__9079 (
            .O(N__41715),
            .I(N__41696));
    LocalMux I__9078 (
            .O(N__41710),
            .I(N__41696));
    InMux I__9077 (
            .O(N__41709),
            .I(N__41691));
    InMux I__9076 (
            .O(N__41708),
            .I(N__41691));
    LocalMux I__9075 (
            .O(N__41705),
            .I(n8828));
    Odrv4 I__9074 (
            .O(N__41696),
            .I(n8828));
    LocalMux I__9073 (
            .O(N__41691),
            .I(n8828));
    InMux I__9072 (
            .O(N__41684),
            .I(n19354));
    InMux I__9071 (
            .O(N__41681),
            .I(n19355));
    InMux I__9070 (
            .O(N__41678),
            .I(n19356));
    InMux I__9069 (
            .O(N__41675),
            .I(n19357));
    InMux I__9068 (
            .O(N__41672),
            .I(n19358));
    InMux I__9067 (
            .O(N__41669),
            .I(n19359));
    InMux I__9066 (
            .O(N__41666),
            .I(n19360));
    InMux I__9065 (
            .O(N__41663),
            .I(bfn_15_14_0_));
    InMux I__9064 (
            .O(N__41660),
            .I(n19362));
    InMux I__9063 (
            .O(N__41657),
            .I(N__41653));
    CascadeMux I__9062 (
            .O(N__41656),
            .I(N__41650));
    LocalMux I__9061 (
            .O(N__41653),
            .I(N__41647));
    InMux I__9060 (
            .O(N__41650),
            .I(N__41643));
    Span4Mux_h I__9059 (
            .O(N__41647),
            .I(N__41640));
    InMux I__9058 (
            .O(N__41646),
            .I(N__41637));
    LocalMux I__9057 (
            .O(N__41643),
            .I(acadc_skipCount_8));
    Odrv4 I__9056 (
            .O(N__41640),
            .I(acadc_skipCount_8));
    LocalMux I__9055 (
            .O(N__41637),
            .I(acadc_skipCount_8));
    InMux I__9054 (
            .O(N__41630),
            .I(N__41627));
    LocalMux I__9053 (
            .O(N__41627),
            .I(N__41620));
    InMux I__9052 (
            .O(N__41626),
            .I(N__41615));
    InMux I__9051 (
            .O(N__41625),
            .I(N__41615));
    InMux I__9050 (
            .O(N__41624),
            .I(N__41612));
    InMux I__9049 (
            .O(N__41623),
            .I(N__41609));
    Span4Mux_v I__9048 (
            .O(N__41620),
            .I(N__41606));
    LocalMux I__9047 (
            .O(N__41615),
            .I(N__41603));
    LocalMux I__9046 (
            .O(N__41612),
            .I(N__41600));
    LocalMux I__9045 (
            .O(N__41609),
            .I(eis_start));
    Odrv4 I__9044 (
            .O(N__41606),
            .I(eis_start));
    Odrv4 I__9043 (
            .O(N__41603),
            .I(eis_start));
    Odrv4 I__9042 (
            .O(N__41600),
            .I(eis_start));
    InMux I__9041 (
            .O(N__41591),
            .I(N__41588));
    LocalMux I__9040 (
            .O(N__41588),
            .I(n21992));
    InMux I__9039 (
            .O(N__41585),
            .I(N__41581));
    CascadeMux I__9038 (
            .O(N__41584),
            .I(N__41578));
    LocalMux I__9037 (
            .O(N__41581),
            .I(N__41575));
    InMux I__9036 (
            .O(N__41578),
            .I(N__41572));
    Span4Mux_h I__9035 (
            .O(N__41575),
            .I(N__41569));
    LocalMux I__9034 (
            .O(N__41572),
            .I(data_idxvec_8));
    Odrv4 I__9033 (
            .O(N__41569),
            .I(data_idxvec_8));
    InMux I__9032 (
            .O(N__41564),
            .I(N__41561));
    LocalMux I__9031 (
            .O(N__41561),
            .I(N__41558));
    Odrv12 I__9030 (
            .O(N__41558),
            .I(buf_data_iac_16));
    CascadeMux I__9029 (
            .O(N__41555),
            .I(n20917_cascade_));
    InMux I__9028 (
            .O(N__41552),
            .I(N__41549));
    LocalMux I__9027 (
            .O(N__41549),
            .I(n21995));
    CascadeMux I__9026 (
            .O(N__41546),
            .I(n20919_cascade_));
    InMux I__9025 (
            .O(N__41543),
            .I(N__41540));
    LocalMux I__9024 (
            .O(N__41540),
            .I(N__41537));
    Span12Mux_h I__9023 (
            .O(N__41537),
            .I(N__41534));
    Odrv12 I__9022 (
            .O(N__41534),
            .I(n22043));
    InMux I__9021 (
            .O(N__41531),
            .I(N__41528));
    LocalMux I__9020 (
            .O(N__41528),
            .I(N__41525));
    Span4Mux_v I__9019 (
            .O(N__41525),
            .I(N__41522));
    Span4Mux_h I__9018 (
            .O(N__41522),
            .I(N__41519));
    Odrv4 I__9017 (
            .O(N__41519),
            .I(n22019));
    CascadeMux I__9016 (
            .O(N__41516),
            .I(n22220_cascade_));
    CascadeMux I__9015 (
            .O(N__41513),
            .I(n22223_cascade_));
    CascadeMux I__9014 (
            .O(N__41510),
            .I(N__41507));
    InMux I__9013 (
            .O(N__41507),
            .I(N__41501));
    InMux I__9012 (
            .O(N__41506),
            .I(N__41501));
    LocalMux I__9011 (
            .O(N__41501),
            .I(N__41495));
    InMux I__9010 (
            .O(N__41500),
            .I(N__41490));
    InMux I__9009 (
            .O(N__41499),
            .I(N__41487));
    InMux I__9008 (
            .O(N__41498),
            .I(N__41484));
    Span4Mux_v I__9007 (
            .O(N__41495),
            .I(N__41481));
    InMux I__9006 (
            .O(N__41494),
            .I(N__41478));
    InMux I__9005 (
            .O(N__41493),
            .I(N__41475));
    LocalMux I__9004 (
            .O(N__41490),
            .I(N__41472));
    LocalMux I__9003 (
            .O(N__41487),
            .I(N__41469));
    LocalMux I__9002 (
            .O(N__41484),
            .I(N__41466));
    Span4Mux_h I__9001 (
            .O(N__41481),
            .I(N__41461));
    LocalMux I__9000 (
            .O(N__41478),
            .I(N__41461));
    LocalMux I__8999 (
            .O(N__41475),
            .I(N__41456));
    Span4Mux_v I__8998 (
            .O(N__41472),
            .I(N__41456));
    Span4Mux_h I__8997 (
            .O(N__41469),
            .I(N__41451));
    Span4Mux_v I__8996 (
            .O(N__41466),
            .I(N__41451));
    Span4Mux_v I__8995 (
            .O(N__41461),
            .I(N__41444));
    Span4Mux_v I__8994 (
            .O(N__41456),
            .I(N__41444));
    Span4Mux_h I__8993 (
            .O(N__41451),
            .I(N__41444));
    Odrv4 I__8992 (
            .O(N__41444),
            .I(comm_buf_0_0));
    CascadeMux I__8991 (
            .O(N__41441),
            .I(N__41438));
    InMux I__8990 (
            .O(N__41438),
            .I(N__41434));
    InMux I__8989 (
            .O(N__41437),
            .I(N__41429));
    LocalMux I__8988 (
            .O(N__41434),
            .I(N__41426));
    InMux I__8987 (
            .O(N__41433),
            .I(N__41423));
    InMux I__8986 (
            .O(N__41432),
            .I(N__41420));
    LocalMux I__8985 (
            .O(N__41429),
            .I(N__41415));
    Span4Mux_v I__8984 (
            .O(N__41426),
            .I(N__41412));
    LocalMux I__8983 (
            .O(N__41423),
            .I(N__41407));
    LocalMux I__8982 (
            .O(N__41420),
            .I(N__41407));
    InMux I__8981 (
            .O(N__41419),
            .I(N__41402));
    InMux I__8980 (
            .O(N__41418),
            .I(N__41402));
    Span4Mux_v I__8979 (
            .O(N__41415),
            .I(N__41395));
    Span4Mux_h I__8978 (
            .O(N__41412),
            .I(N__41395));
    Span4Mux_v I__8977 (
            .O(N__41407),
            .I(N__41395));
    LocalMux I__8976 (
            .O(N__41402),
            .I(iac_raw_buf_N_737));
    Odrv4 I__8975 (
            .O(N__41395),
            .I(iac_raw_buf_N_737));
    InMux I__8974 (
            .O(N__41390),
            .I(N__41383));
    InMux I__8973 (
            .O(N__41389),
            .I(N__41383));
    InMux I__8972 (
            .O(N__41388),
            .I(N__41379));
    LocalMux I__8971 (
            .O(N__41383),
            .I(N__41376));
    CascadeMux I__8970 (
            .O(N__41382),
            .I(N__41372));
    LocalMux I__8969 (
            .O(N__41379),
            .I(N__41367));
    Span4Mux_h I__8968 (
            .O(N__41376),
            .I(N__41364));
    InMux I__8967 (
            .O(N__41375),
            .I(N__41361));
    InMux I__8966 (
            .O(N__41372),
            .I(N__41358));
    InMux I__8965 (
            .O(N__41371),
            .I(N__41353));
    InMux I__8964 (
            .O(N__41370),
            .I(N__41353));
    Span4Mux_h I__8963 (
            .O(N__41367),
            .I(N__41348));
    Span4Mux_h I__8962 (
            .O(N__41364),
            .I(N__41348));
    LocalMux I__8961 (
            .O(N__41361),
            .I(n12397));
    LocalMux I__8960 (
            .O(N__41358),
            .I(n12397));
    LocalMux I__8959 (
            .O(N__41353),
            .I(n12397));
    Odrv4 I__8958 (
            .O(N__41348),
            .I(n12397));
    IoInMux I__8957 (
            .O(N__41339),
            .I(N__41336));
    LocalMux I__8956 (
            .O(N__41336),
            .I(N__41333));
    Span4Mux_s2_h I__8955 (
            .O(N__41333),
            .I(N__41330));
    Span4Mux_h I__8954 (
            .O(N__41330),
            .I(N__41327));
    Sp12to4 I__8953 (
            .O(N__41327),
            .I(N__41324));
    Span12Mux_s10_v I__8952 (
            .O(N__41324),
            .I(N__41319));
    InMux I__8951 (
            .O(N__41323),
            .I(N__41316));
    InMux I__8950 (
            .O(N__41322),
            .I(N__41313));
    Span12Mux_h I__8949 (
            .O(N__41319),
            .I(N__41308));
    LocalMux I__8948 (
            .O(N__41316),
            .I(N__41308));
    LocalMux I__8947 (
            .O(N__41313),
            .I(VAC_OSR0));
    Odrv12 I__8946 (
            .O(N__41308),
            .I(VAC_OSR0));
    InMux I__8945 (
            .O(N__41303),
            .I(N__41300));
    LocalMux I__8944 (
            .O(N__41300),
            .I(N__41297));
    Span4Mux_v I__8943 (
            .O(N__41297),
            .I(N__41294));
    Odrv4 I__8942 (
            .O(N__41294),
            .I(n21046));
    InMux I__8941 (
            .O(N__41291),
            .I(N__41288));
    LocalMux I__8940 (
            .O(N__41288),
            .I(N__41285));
    Span4Mux_h I__8939 (
            .O(N__41285),
            .I(N__41280));
    InMux I__8938 (
            .O(N__41284),
            .I(N__41275));
    InMux I__8937 (
            .O(N__41283),
            .I(N__41275));
    Odrv4 I__8936 (
            .O(N__41280),
            .I(acadc_skipCount_0));
    LocalMux I__8935 (
            .O(N__41275),
            .I(acadc_skipCount_0));
    InMux I__8934 (
            .O(N__41270),
            .I(N__41267));
    LocalMux I__8933 (
            .O(N__41267),
            .I(N__41264));
    Span4Mux_h I__8932 (
            .O(N__41264),
            .I(N__41261));
    Odrv4 I__8931 (
            .O(N__41261),
            .I(n19_adj_1487));
    CascadeMux I__8930 (
            .O(N__41258),
            .I(N__41255));
    InMux I__8929 (
            .O(N__41255),
            .I(N__41252));
    LocalMux I__8928 (
            .O(N__41252),
            .I(N__41248));
    CascadeMux I__8927 (
            .O(N__41251),
            .I(N__41245));
    Span12Mux_h I__8926 (
            .O(N__41248),
            .I(N__41242));
    InMux I__8925 (
            .O(N__41245),
            .I(N__41239));
    Odrv12 I__8924 (
            .O(N__41242),
            .I(buf_readRTD_0));
    LocalMux I__8923 (
            .O(N__41239),
            .I(buf_readRTD_0));
    CascadeMux I__8922 (
            .O(N__41234),
            .I(N__41230));
    InMux I__8921 (
            .O(N__41233),
            .I(N__41227));
    InMux I__8920 (
            .O(N__41230),
            .I(N__41224));
    LocalMux I__8919 (
            .O(N__41227),
            .I(N__41221));
    LocalMux I__8918 (
            .O(N__41224),
            .I(data_idxvec_0));
    Odrv12 I__8917 (
            .O(N__41221),
            .I(data_idxvec_0));
    InMux I__8916 (
            .O(N__41216),
            .I(N__41213));
    LocalMux I__8915 (
            .O(N__41213),
            .I(N__41210));
    Odrv4 I__8914 (
            .O(N__41210),
            .I(n20973));
    CascadeMux I__8913 (
            .O(N__41207),
            .I(n26_cascade_));
    InMux I__8912 (
            .O(N__41204),
            .I(N__41201));
    LocalMux I__8911 (
            .O(N__41201),
            .I(n21998));
    InMux I__8910 (
            .O(N__41198),
            .I(N__41195));
    LocalMux I__8909 (
            .O(N__41195),
            .I(N__41192));
    Span4Mux_h I__8908 (
            .O(N__41192),
            .I(N__41189));
    Odrv4 I__8907 (
            .O(N__41189),
            .I(n16_adj_1488));
    InMux I__8906 (
            .O(N__41186),
            .I(N__41183));
    LocalMux I__8905 (
            .O(N__41183),
            .I(n22004));
    CascadeMux I__8904 (
            .O(N__41180),
            .I(n22007_cascade_));
    InMux I__8903 (
            .O(N__41177),
            .I(N__41174));
    LocalMux I__8902 (
            .O(N__41174),
            .I(n22001));
    CascadeMux I__8901 (
            .O(N__41171),
            .I(n30_adj_1486_cascade_));
    CascadeMux I__8900 (
            .O(N__41168),
            .I(N__41164));
    CascadeMux I__8899 (
            .O(N__41167),
            .I(N__41159));
    InMux I__8898 (
            .O(N__41164),
            .I(N__41150));
    InMux I__8897 (
            .O(N__41163),
            .I(N__41150));
    InMux I__8896 (
            .O(N__41162),
            .I(N__41150));
    InMux I__8895 (
            .O(N__41159),
            .I(N__41147));
    InMux I__8894 (
            .O(N__41158),
            .I(N__41144));
    InMux I__8893 (
            .O(N__41157),
            .I(N__41141));
    LocalMux I__8892 (
            .O(N__41150),
            .I(N__41138));
    LocalMux I__8891 (
            .O(N__41147),
            .I(N__41133));
    LocalMux I__8890 (
            .O(N__41144),
            .I(N__41133));
    LocalMux I__8889 (
            .O(N__41141),
            .I(N__41130));
    Span4Mux_h I__8888 (
            .O(N__41138),
            .I(N__41127));
    Span4Mux_h I__8887 (
            .O(N__41133),
            .I(N__41124));
    Span4Mux_v I__8886 (
            .O(N__41130),
            .I(N__41121));
    Span4Mux_h I__8885 (
            .O(N__41127),
            .I(N__41118));
    Span4Mux_v I__8884 (
            .O(N__41124),
            .I(N__41115));
    Odrv4 I__8883 (
            .O(N__41121),
            .I(comm_buf_1_0));
    Odrv4 I__8882 (
            .O(N__41118),
            .I(comm_buf_1_0));
    Odrv4 I__8881 (
            .O(N__41115),
            .I(comm_buf_1_0));
    CascadeMux I__8880 (
            .O(N__41108),
            .I(n12242_cascade_));
    CascadeMux I__8879 (
            .O(N__41105),
            .I(n20599_cascade_));
    InMux I__8878 (
            .O(N__41102),
            .I(N__41099));
    LocalMux I__8877 (
            .O(N__41099),
            .I(N__41096));
    Odrv12 I__8876 (
            .O(N__41096),
            .I(n5));
    IoInMux I__8875 (
            .O(N__41093),
            .I(N__41090));
    LocalMux I__8874 (
            .O(N__41090),
            .I(N__41087));
    IoSpan4Mux I__8873 (
            .O(N__41087),
            .I(N__41084));
    Span4Mux_s3_v I__8872 (
            .O(N__41084),
            .I(N__41081));
    Span4Mux_v I__8871 (
            .O(N__41081),
            .I(N__41078));
    Sp12to4 I__8870 (
            .O(N__41078),
            .I(N__41074));
    InMux I__8869 (
            .O(N__41077),
            .I(N__41070));
    Span12Mux_h I__8868 (
            .O(N__41074),
            .I(N__41067));
    InMux I__8867 (
            .O(N__41073),
            .I(N__41064));
    LocalMux I__8866 (
            .O(N__41070),
            .I(N__41061));
    Odrv12 I__8865 (
            .O(N__41067),
            .I(IAC_FLT1));
    LocalMux I__8864 (
            .O(N__41064),
            .I(IAC_FLT1));
    Odrv4 I__8863 (
            .O(N__41061),
            .I(IAC_FLT1));
    CascadeMux I__8862 (
            .O(N__41054),
            .I(N__41046));
    InMux I__8861 (
            .O(N__41053),
            .I(N__41042));
    InMux I__8860 (
            .O(N__41052),
            .I(N__41037));
    InMux I__8859 (
            .O(N__41051),
            .I(N__41037));
    CascadeMux I__8858 (
            .O(N__41050),
            .I(N__41032));
    InMux I__8857 (
            .O(N__41049),
            .I(N__41027));
    InMux I__8856 (
            .O(N__41046),
            .I(N__41027));
    InMux I__8855 (
            .O(N__41045),
            .I(N__41024));
    LocalMux I__8854 (
            .O(N__41042),
            .I(N__41017));
    LocalMux I__8853 (
            .O(N__41037),
            .I(N__41014));
    InMux I__8852 (
            .O(N__41036),
            .I(N__41011));
    InMux I__8851 (
            .O(N__41035),
            .I(N__41006));
    InMux I__8850 (
            .O(N__41032),
            .I(N__41006));
    LocalMux I__8849 (
            .O(N__41027),
            .I(N__41003));
    LocalMux I__8848 (
            .O(N__41024),
            .I(N__41000));
    InMux I__8847 (
            .O(N__41023),
            .I(N__40997));
    InMux I__8846 (
            .O(N__41022),
            .I(N__40994));
    InMux I__8845 (
            .O(N__41021),
            .I(N__40991));
    InMux I__8844 (
            .O(N__41020),
            .I(N__40988));
    Span4Mux_h I__8843 (
            .O(N__41017),
            .I(N__40985));
    Span4Mux_v I__8842 (
            .O(N__41014),
            .I(N__40982));
    LocalMux I__8841 (
            .O(N__41011),
            .I(N__40973));
    LocalMux I__8840 (
            .O(N__41006),
            .I(N__40973));
    Span4Mux_h I__8839 (
            .O(N__41003),
            .I(N__40973));
    Span4Mux_h I__8838 (
            .O(N__41000),
            .I(N__40973));
    LocalMux I__8837 (
            .O(N__40997),
            .I(eis_state_1));
    LocalMux I__8836 (
            .O(N__40994),
            .I(eis_state_1));
    LocalMux I__8835 (
            .O(N__40991),
            .I(eis_state_1));
    LocalMux I__8834 (
            .O(N__40988),
            .I(eis_state_1));
    Odrv4 I__8833 (
            .O(N__40985),
            .I(eis_state_1));
    Odrv4 I__8832 (
            .O(N__40982),
            .I(eis_state_1));
    Odrv4 I__8831 (
            .O(N__40973),
            .I(eis_state_1));
    InMux I__8830 (
            .O(N__40958),
            .I(N__40955));
    LocalMux I__8829 (
            .O(N__40955),
            .I(N__40952));
    Span12Mux_h I__8828 (
            .O(N__40952),
            .I(N__40949));
    Odrv12 I__8827 (
            .O(N__40949),
            .I(buf_data_iac_8));
    InMux I__8826 (
            .O(N__40946),
            .I(N__40942));
    CascadeMux I__8825 (
            .O(N__40945),
            .I(N__40939));
    LocalMux I__8824 (
            .O(N__40942),
            .I(N__40936));
    InMux I__8823 (
            .O(N__40939),
            .I(N__40933));
    Span4Mux_h I__8822 (
            .O(N__40936),
            .I(N__40930));
    LocalMux I__8821 (
            .O(N__40933),
            .I(data_idxvec_12));
    Odrv4 I__8820 (
            .O(N__40930),
            .I(data_idxvec_12));
    CascadeMux I__8819 (
            .O(N__40925),
            .I(N__40922));
    InMux I__8818 (
            .O(N__40922),
            .I(N__40919));
    LocalMux I__8817 (
            .O(N__40919),
            .I(N__40916));
    Odrv12 I__8816 (
            .O(N__40916),
            .I(n20983));
    InMux I__8815 (
            .O(N__40913),
            .I(N__40910));
    LocalMux I__8814 (
            .O(N__40910),
            .I(N__40906));
    CascadeMux I__8813 (
            .O(N__40909),
            .I(N__40903));
    Span4Mux_h I__8812 (
            .O(N__40906),
            .I(N__40900));
    InMux I__8811 (
            .O(N__40903),
            .I(N__40897));
    Span4Mux_v I__8810 (
            .O(N__40900),
            .I(N__40894));
    LocalMux I__8809 (
            .O(N__40897),
            .I(N__40890));
    Span4Mux_h I__8808 (
            .O(N__40894),
            .I(N__40887));
    InMux I__8807 (
            .O(N__40893),
            .I(N__40884));
    Span12Mux_v I__8806 (
            .O(N__40890),
            .I(N__40881));
    Span4Mux_h I__8805 (
            .O(N__40887),
            .I(N__40878));
    LocalMux I__8804 (
            .O(N__40884),
            .I(buf_adcdata_iac_19));
    Odrv12 I__8803 (
            .O(N__40881),
            .I(buf_adcdata_iac_19));
    Odrv4 I__8802 (
            .O(N__40878),
            .I(buf_adcdata_iac_19));
    InMux I__8801 (
            .O(N__40871),
            .I(N__40868));
    LocalMux I__8800 (
            .O(N__40868),
            .I(n22082));
    InMux I__8799 (
            .O(N__40865),
            .I(N__40861));
    CascadeMux I__8798 (
            .O(N__40864),
            .I(N__40858));
    LocalMux I__8797 (
            .O(N__40861),
            .I(N__40855));
    InMux I__8796 (
            .O(N__40858),
            .I(N__40852));
    Span4Mux_h I__8795 (
            .O(N__40855),
            .I(N__40849));
    LocalMux I__8794 (
            .O(N__40852),
            .I(data_idxvec_11));
    Odrv4 I__8793 (
            .O(N__40849),
            .I(data_idxvec_11));
    InMux I__8792 (
            .O(N__40844),
            .I(N__40841));
    LocalMux I__8791 (
            .O(N__40841),
            .I(N__40838));
    Span4Mux_h I__8790 (
            .O(N__40838),
            .I(N__40835));
    Span4Mux_h I__8789 (
            .O(N__40835),
            .I(N__40832));
    Odrv4 I__8788 (
            .O(N__40832),
            .I(buf_data_iac_19));
    CascadeMux I__8787 (
            .O(N__40829),
            .I(n26_adj_1541_cascade_));
    CascadeMux I__8786 (
            .O(N__40826),
            .I(n20837_cascade_));
    InMux I__8785 (
            .O(N__40823),
            .I(N__40820));
    LocalMux I__8784 (
            .O(N__40820),
            .I(n22085));
    CascadeMux I__8783 (
            .O(N__40817),
            .I(n22094_cascade_));
    InMux I__8782 (
            .O(N__40814),
            .I(N__40811));
    LocalMux I__8781 (
            .O(N__40811),
            .I(N__40808));
    Span12Mux_v I__8780 (
            .O(N__40808),
            .I(N__40805));
    Odrv12 I__8779 (
            .O(N__40805),
            .I(n20828));
    InMux I__8778 (
            .O(N__40802),
            .I(N__40798));
    CascadeMux I__8777 (
            .O(N__40801),
            .I(N__40794));
    LocalMux I__8776 (
            .O(N__40798),
            .I(N__40789));
    InMux I__8775 (
            .O(N__40797),
            .I(N__40786));
    InMux I__8774 (
            .O(N__40794),
            .I(N__40783));
    InMux I__8773 (
            .O(N__40793),
            .I(N__40780));
    InMux I__8772 (
            .O(N__40792),
            .I(N__40777));
    Span4Mux_v I__8771 (
            .O(N__40789),
            .I(N__40773));
    LocalMux I__8770 (
            .O(N__40786),
            .I(N__40770));
    LocalMux I__8769 (
            .O(N__40783),
            .I(N__40765));
    LocalMux I__8768 (
            .O(N__40780),
            .I(N__40765));
    LocalMux I__8767 (
            .O(N__40777),
            .I(N__40762));
    InMux I__8766 (
            .O(N__40776),
            .I(N__40759));
    Span4Mux_v I__8765 (
            .O(N__40773),
            .I(N__40754));
    Span4Mux_v I__8764 (
            .O(N__40770),
            .I(N__40751));
    Span4Mux_v I__8763 (
            .O(N__40765),
            .I(N__40748));
    Span4Mux_v I__8762 (
            .O(N__40762),
            .I(N__40743));
    LocalMux I__8761 (
            .O(N__40759),
            .I(N__40743));
    InMux I__8760 (
            .O(N__40758),
            .I(N__40740));
    InMux I__8759 (
            .O(N__40757),
            .I(N__40737));
    Span4Mux_h I__8758 (
            .O(N__40754),
            .I(N__40733));
    Span4Mux_v I__8757 (
            .O(N__40751),
            .I(N__40730));
    Span4Mux_h I__8756 (
            .O(N__40748),
            .I(N__40727));
    Span4Mux_h I__8755 (
            .O(N__40743),
            .I(N__40724));
    LocalMux I__8754 (
            .O(N__40740),
            .I(N__40721));
    LocalMux I__8753 (
            .O(N__40737),
            .I(N__40718));
    InMux I__8752 (
            .O(N__40736),
            .I(N__40715));
    Odrv4 I__8751 (
            .O(N__40733),
            .I(comm_rx_buf_3));
    Odrv4 I__8750 (
            .O(N__40730),
            .I(comm_rx_buf_3));
    Odrv4 I__8749 (
            .O(N__40727),
            .I(comm_rx_buf_3));
    Odrv4 I__8748 (
            .O(N__40724),
            .I(comm_rx_buf_3));
    Odrv12 I__8747 (
            .O(N__40721),
            .I(comm_rx_buf_3));
    Odrv4 I__8746 (
            .O(N__40718),
            .I(comm_rx_buf_3));
    LocalMux I__8745 (
            .O(N__40715),
            .I(comm_rx_buf_3));
    CascadeMux I__8744 (
            .O(N__40700),
            .I(n22097_cascade_));
    SRMux I__8743 (
            .O(N__40697),
            .I(N__40693));
    SRMux I__8742 (
            .O(N__40696),
            .I(N__40690));
    LocalMux I__8741 (
            .O(N__40693),
            .I(N__40687));
    LocalMux I__8740 (
            .O(N__40690),
            .I(N__40684));
    Span4Mux_v I__8739 (
            .O(N__40687),
            .I(N__40681));
    Span4Mux_h I__8738 (
            .O(N__40684),
            .I(N__40678));
    Span4Mux_h I__8737 (
            .O(N__40681),
            .I(N__40673));
    Span4Mux_h I__8736 (
            .O(N__40678),
            .I(N__40673));
    Sp12to4 I__8735 (
            .O(N__40673),
            .I(N__40670));
    Odrv12 I__8734 (
            .O(N__40670),
            .I(flagcntwd));
    CEMux I__8733 (
            .O(N__40667),
            .I(N__40664));
    LocalMux I__8732 (
            .O(N__40664),
            .I(n11406));
    CascadeMux I__8731 (
            .O(N__40661),
            .I(N__40658));
    InMux I__8730 (
            .O(N__40658),
            .I(N__40655));
    LocalMux I__8729 (
            .O(N__40655),
            .I(N__40651));
    InMux I__8728 (
            .O(N__40654),
            .I(N__40647));
    Span4Mux_v I__8727 (
            .O(N__40651),
            .I(N__40642));
    InMux I__8726 (
            .O(N__40650),
            .I(N__40639));
    LocalMux I__8725 (
            .O(N__40647),
            .I(N__40635));
    InMux I__8724 (
            .O(N__40646),
            .I(N__40632));
    InMux I__8723 (
            .O(N__40645),
            .I(N__40629));
    Span4Mux_h I__8722 (
            .O(N__40642),
            .I(N__40624));
    LocalMux I__8721 (
            .O(N__40639),
            .I(N__40624));
    InMux I__8720 (
            .O(N__40638),
            .I(N__40621));
    Span4Mux_v I__8719 (
            .O(N__40635),
            .I(N__40614));
    LocalMux I__8718 (
            .O(N__40632),
            .I(N__40614));
    LocalMux I__8717 (
            .O(N__40629),
            .I(N__40611));
    Span4Mux_v I__8716 (
            .O(N__40624),
            .I(N__40606));
    LocalMux I__8715 (
            .O(N__40621),
            .I(N__40606));
    InMux I__8714 (
            .O(N__40620),
            .I(N__40603));
    InMux I__8713 (
            .O(N__40619),
            .I(N__40600));
    Span4Mux_v I__8712 (
            .O(N__40614),
            .I(N__40596));
    Span12Mux_h I__8711 (
            .O(N__40611),
            .I(N__40593));
    Span4Mux_v I__8710 (
            .O(N__40606),
            .I(N__40586));
    LocalMux I__8709 (
            .O(N__40603),
            .I(N__40586));
    LocalMux I__8708 (
            .O(N__40600),
            .I(N__40586));
    InMux I__8707 (
            .O(N__40599),
            .I(N__40583));
    Odrv4 I__8706 (
            .O(N__40596),
            .I(comm_rx_buf_4));
    Odrv12 I__8705 (
            .O(N__40593),
            .I(comm_rx_buf_4));
    Odrv4 I__8704 (
            .O(N__40586),
            .I(comm_rx_buf_4));
    LocalMux I__8703 (
            .O(N__40583),
            .I(comm_rx_buf_4));
    CascadeMux I__8702 (
            .O(N__40574),
            .I(n30_adj_1539_cascade_));
    InMux I__8701 (
            .O(N__40571),
            .I(N__40564));
    InMux I__8700 (
            .O(N__40570),
            .I(N__40564));
    CascadeMux I__8699 (
            .O(N__40569),
            .I(N__40559));
    LocalMux I__8698 (
            .O(N__40564),
            .I(N__40556));
    InMux I__8697 (
            .O(N__40563),
            .I(N__40551));
    InMux I__8696 (
            .O(N__40562),
            .I(N__40551));
    InMux I__8695 (
            .O(N__40559),
            .I(N__40548));
    Span4Mux_v I__8694 (
            .O(N__40556),
            .I(N__40543));
    LocalMux I__8693 (
            .O(N__40551),
            .I(N__40543));
    LocalMux I__8692 (
            .O(N__40548),
            .I(N__40538));
    Span4Mux_h I__8691 (
            .O(N__40543),
            .I(N__40538));
    Odrv4 I__8690 (
            .O(N__40538),
            .I(comm_cmd_7));
    CascadeMux I__8689 (
            .O(N__40535),
            .I(n20621_cascade_));
    CascadeMux I__8688 (
            .O(N__40532),
            .I(n25_adj_1619_cascade_));
    InMux I__8687 (
            .O(N__40529),
            .I(N__40526));
    LocalMux I__8686 (
            .O(N__40526),
            .I(N__40516));
    InMux I__8685 (
            .O(N__40525),
            .I(N__40501));
    InMux I__8684 (
            .O(N__40524),
            .I(N__40501));
    InMux I__8683 (
            .O(N__40523),
            .I(N__40501));
    InMux I__8682 (
            .O(N__40522),
            .I(N__40501));
    InMux I__8681 (
            .O(N__40521),
            .I(N__40501));
    InMux I__8680 (
            .O(N__40520),
            .I(N__40501));
    InMux I__8679 (
            .O(N__40519),
            .I(N__40501));
    Odrv12 I__8678 (
            .O(N__40516),
            .I(\comm_spi.n16869 ));
    LocalMux I__8677 (
            .O(N__40501),
            .I(\comm_spi.n16869 ));
    InMux I__8676 (
            .O(N__40496),
            .I(N__40493));
    LocalMux I__8675 (
            .O(N__40493),
            .I(N__40490));
    Span4Mux_h I__8674 (
            .O(N__40490),
            .I(N__40487));
    Odrv4 I__8673 (
            .O(N__40487),
            .I(n7_adj_1609));
    InMux I__8672 (
            .O(N__40484),
            .I(N__40480));
    InMux I__8671 (
            .O(N__40483),
            .I(N__40476));
    LocalMux I__8670 (
            .O(N__40480),
            .I(N__40473));
    InMux I__8669 (
            .O(N__40479),
            .I(N__40470));
    LocalMux I__8668 (
            .O(N__40476),
            .I(N__40467));
    Span12Mux_h I__8667 (
            .O(N__40473),
            .I(N__40464));
    LocalMux I__8666 (
            .O(N__40470),
            .I(buf_dds1_11));
    Odrv4 I__8665 (
            .O(N__40467),
            .I(buf_dds1_11));
    Odrv12 I__8664 (
            .O(N__40464),
            .I(buf_dds1_11));
    InMux I__8663 (
            .O(N__40457),
            .I(N__40453));
    CascadeMux I__8662 (
            .O(N__40456),
            .I(N__40450));
    LocalMux I__8661 (
            .O(N__40453),
            .I(N__40446));
    InMux I__8660 (
            .O(N__40450),
            .I(N__40443));
    InMux I__8659 (
            .O(N__40449),
            .I(N__40440));
    Span4Mux_v I__8658 (
            .O(N__40446),
            .I(N__40437));
    LocalMux I__8657 (
            .O(N__40443),
            .I(N__40434));
    LocalMux I__8656 (
            .O(N__40440),
            .I(N__40427));
    Span4Mux_h I__8655 (
            .O(N__40437),
            .I(N__40427));
    Span4Mux_v I__8654 (
            .O(N__40434),
            .I(N__40427));
    Odrv4 I__8653 (
            .O(N__40427),
            .I(buf_dds0_11));
    CascadeMux I__8652 (
            .O(N__40424),
            .I(n21506_cascade_));
    InMux I__8651 (
            .O(N__40421),
            .I(N__40418));
    LocalMux I__8650 (
            .O(N__40418),
            .I(N__40415));
    Span12Mux_h I__8649 (
            .O(N__40415),
            .I(N__40412));
    Span12Mux_v I__8648 (
            .O(N__40412),
            .I(N__40409));
    Odrv12 I__8647 (
            .O(N__40409),
            .I(n21067));
    CascadeMux I__8646 (
            .O(N__40406),
            .I(N__40403));
    InMux I__8645 (
            .O(N__40403),
            .I(N__40400));
    LocalMux I__8644 (
            .O(N__40400),
            .I(N__40397));
    Span4Mux_h I__8643 (
            .O(N__40397),
            .I(N__40394));
    Span4Mux_v I__8642 (
            .O(N__40394),
            .I(N__40391));
    Odrv4 I__8641 (
            .O(N__40391),
            .I(n23_adj_1538));
    InMux I__8640 (
            .O(N__40388),
            .I(N__40385));
    LocalMux I__8639 (
            .O(N__40385),
            .I(n22028));
    InMux I__8638 (
            .O(N__40382),
            .I(N__40378));
    CascadeMux I__8637 (
            .O(N__40381),
            .I(N__40375));
    LocalMux I__8636 (
            .O(N__40378),
            .I(N__40372));
    InMux I__8635 (
            .O(N__40375),
            .I(N__40369));
    Span4Mux_v I__8634 (
            .O(N__40372),
            .I(N__40366));
    LocalMux I__8633 (
            .O(N__40369),
            .I(N__40363));
    Sp12to4 I__8632 (
            .O(N__40366),
            .I(N__40359));
    Span4Mux_h I__8631 (
            .O(N__40363),
            .I(N__40356));
    InMux I__8630 (
            .O(N__40362),
            .I(N__40353));
    Span12Mux_h I__8629 (
            .O(N__40359),
            .I(N__40350));
    Span4Mux_h I__8628 (
            .O(N__40356),
            .I(N__40347));
    LocalMux I__8627 (
            .O(N__40353),
            .I(buf_adcdata_iac_20));
    Odrv12 I__8626 (
            .O(N__40350),
            .I(buf_adcdata_iac_20));
    Odrv4 I__8625 (
            .O(N__40347),
            .I(buf_adcdata_iac_20));
    InMux I__8624 (
            .O(N__40340),
            .I(N__40337));
    LocalMux I__8623 (
            .O(N__40337),
            .I(N__40334));
    Span4Mux_h I__8622 (
            .O(N__40334),
            .I(N__40330));
    InMux I__8621 (
            .O(N__40333),
            .I(N__40327));
    Span4Mux_v I__8620 (
            .O(N__40330),
            .I(N__40323));
    LocalMux I__8619 (
            .O(N__40327),
            .I(N__40320));
    InMux I__8618 (
            .O(N__40326),
            .I(N__40317));
    Span4Mux_v I__8617 (
            .O(N__40323),
            .I(N__40314));
    Odrv4 I__8616 (
            .O(N__40320),
            .I(buf_dds0_12));
    LocalMux I__8615 (
            .O(N__40317),
            .I(buf_dds0_12));
    Odrv4 I__8614 (
            .O(N__40314),
            .I(buf_dds0_12));
    CascadeMux I__8613 (
            .O(N__40307),
            .I(n22088_cascade_));
    InMux I__8612 (
            .O(N__40304),
            .I(N__40301));
    LocalMux I__8611 (
            .O(N__40301),
            .I(N__40298));
    Span4Mux_h I__8610 (
            .O(N__40298),
            .I(N__40295));
    Span4Mux_v I__8609 (
            .O(N__40295),
            .I(N__40290));
    InMux I__8608 (
            .O(N__40294),
            .I(N__40287));
    InMux I__8607 (
            .O(N__40293),
            .I(N__40284));
    Span4Mux_h I__8606 (
            .O(N__40290),
            .I(N__40281));
    LocalMux I__8605 (
            .O(N__40287),
            .I(buf_dds1_12));
    LocalMux I__8604 (
            .O(N__40284),
            .I(buf_dds1_12));
    Odrv4 I__8603 (
            .O(N__40281),
            .I(buf_dds1_12));
    CascadeMux I__8602 (
            .O(N__40274),
            .I(n22091_cascade_));
    InMux I__8601 (
            .O(N__40271),
            .I(N__40268));
    LocalMux I__8600 (
            .O(N__40268),
            .I(N__40265));
    Span4Mux_v I__8599 (
            .O(N__40265),
            .I(N__40262));
    Sp12to4 I__8598 (
            .O(N__40262),
            .I(N__40259));
    Odrv12 I__8597 (
            .O(N__40259),
            .I(n22205));
    InMux I__8596 (
            .O(N__40256),
            .I(N__40253));
    LocalMux I__8595 (
            .O(N__40253),
            .I(n22031));
    CascadeMux I__8594 (
            .O(N__40250),
            .I(n20844_cascade_));
    InMux I__8593 (
            .O(N__40247),
            .I(N__40241));
    InMux I__8592 (
            .O(N__40246),
            .I(N__40238));
    InMux I__8591 (
            .O(N__40245),
            .I(N__40235));
    InMux I__8590 (
            .O(N__40244),
            .I(N__40230));
    LocalMux I__8589 (
            .O(N__40241),
            .I(N__40225));
    LocalMux I__8588 (
            .O(N__40238),
            .I(N__40225));
    LocalMux I__8587 (
            .O(N__40235),
            .I(N__40222));
    InMux I__8586 (
            .O(N__40234),
            .I(N__40219));
    InMux I__8585 (
            .O(N__40233),
            .I(N__40216));
    LocalMux I__8584 (
            .O(N__40230),
            .I(N__40212));
    Span4Mux_v I__8583 (
            .O(N__40225),
            .I(N__40205));
    Span4Mux_v I__8582 (
            .O(N__40222),
            .I(N__40205));
    LocalMux I__8581 (
            .O(N__40219),
            .I(N__40205));
    LocalMux I__8580 (
            .O(N__40216),
            .I(N__40202));
    InMux I__8579 (
            .O(N__40215),
            .I(N__40199));
    Span4Mux_v I__8578 (
            .O(N__40212),
            .I(N__40188));
    Span4Mux_h I__8577 (
            .O(N__40205),
            .I(N__40188));
    Span4Mux_v I__8576 (
            .O(N__40202),
            .I(N__40188));
    LocalMux I__8575 (
            .O(N__40199),
            .I(N__40188));
    InMux I__8574 (
            .O(N__40198),
            .I(N__40185));
    InMux I__8573 (
            .O(N__40197),
            .I(N__40182));
    Odrv4 I__8572 (
            .O(N__40188),
            .I(comm_rx_buf_6));
    LocalMux I__8571 (
            .O(N__40185),
            .I(comm_rx_buf_6));
    LocalMux I__8570 (
            .O(N__40182),
            .I(comm_rx_buf_6));
    InMux I__8569 (
            .O(N__40175),
            .I(N__40172));
    LocalMux I__8568 (
            .O(N__40172),
            .I(N__40167));
    InMux I__8567 (
            .O(N__40171),
            .I(N__40164));
    InMux I__8566 (
            .O(N__40170),
            .I(N__40157));
    Span4Mux_v I__8565 (
            .O(N__40167),
            .I(N__40152));
    LocalMux I__8564 (
            .O(N__40164),
            .I(N__40152));
    InMux I__8563 (
            .O(N__40163),
            .I(N__40143));
    InMux I__8562 (
            .O(N__40162),
            .I(N__40143));
    InMux I__8561 (
            .O(N__40161),
            .I(N__40143));
    InMux I__8560 (
            .O(N__40160),
            .I(N__40143));
    LocalMux I__8559 (
            .O(N__40157),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__8558 (
            .O(N__40152),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__8557 (
            .O(N__40143),
            .I(\ADC_VDC.genclk.div_state_1 ));
    ClkMux I__8556 (
            .O(N__40136),
            .I(N__40128));
    ClkMux I__8555 (
            .O(N__40135),
            .I(N__40125));
    ClkMux I__8554 (
            .O(N__40134),
            .I(N__40122));
    ClkMux I__8553 (
            .O(N__40133),
            .I(N__40113));
    ClkMux I__8552 (
            .O(N__40132),
            .I(N__40104));
    ClkMux I__8551 (
            .O(N__40131),
            .I(N__40101));
    LocalMux I__8550 (
            .O(N__40128),
            .I(N__40098));
    LocalMux I__8549 (
            .O(N__40125),
            .I(N__40093));
    LocalMux I__8548 (
            .O(N__40122),
            .I(N__40093));
    ClkMux I__8547 (
            .O(N__40121),
            .I(N__40090));
    ClkMux I__8546 (
            .O(N__40120),
            .I(N__40085));
    ClkMux I__8545 (
            .O(N__40119),
            .I(N__40082));
    ClkMux I__8544 (
            .O(N__40118),
            .I(N__40079));
    ClkMux I__8543 (
            .O(N__40117),
            .I(N__40076));
    ClkMux I__8542 (
            .O(N__40116),
            .I(N__40073));
    LocalMux I__8541 (
            .O(N__40113),
            .I(N__40070));
    ClkMux I__8540 (
            .O(N__40112),
            .I(N__40067));
    ClkMux I__8539 (
            .O(N__40111),
            .I(N__40064));
    ClkMux I__8538 (
            .O(N__40110),
            .I(N__40061));
    ClkMux I__8537 (
            .O(N__40109),
            .I(N__40057));
    ClkMux I__8536 (
            .O(N__40108),
            .I(N__40054));
    ClkMux I__8535 (
            .O(N__40107),
            .I(N__40050));
    LocalMux I__8534 (
            .O(N__40104),
            .I(N__40045));
    LocalMux I__8533 (
            .O(N__40101),
            .I(N__40042));
    Span4Mux_v I__8532 (
            .O(N__40098),
            .I(N__40035));
    Span4Mux_h I__8531 (
            .O(N__40093),
            .I(N__40035));
    LocalMux I__8530 (
            .O(N__40090),
            .I(N__40035));
    IoInMux I__8529 (
            .O(N__40089),
            .I(N__40031));
    ClkMux I__8528 (
            .O(N__40088),
            .I(N__40028));
    LocalMux I__8527 (
            .O(N__40085),
            .I(N__40025));
    LocalMux I__8526 (
            .O(N__40082),
            .I(N__40018));
    LocalMux I__8525 (
            .O(N__40079),
            .I(N__40018));
    LocalMux I__8524 (
            .O(N__40076),
            .I(N__40018));
    LocalMux I__8523 (
            .O(N__40073),
            .I(N__40015));
    Span4Mux_v I__8522 (
            .O(N__40070),
            .I(N__40010));
    LocalMux I__8521 (
            .O(N__40067),
            .I(N__40010));
    LocalMux I__8520 (
            .O(N__40064),
            .I(N__40007));
    LocalMux I__8519 (
            .O(N__40061),
            .I(N__40004));
    ClkMux I__8518 (
            .O(N__40060),
            .I(N__40001));
    LocalMux I__8517 (
            .O(N__40057),
            .I(N__39996));
    LocalMux I__8516 (
            .O(N__40054),
            .I(N__39996));
    ClkMux I__8515 (
            .O(N__40053),
            .I(N__39993));
    LocalMux I__8514 (
            .O(N__40050),
            .I(N__39990));
    ClkMux I__8513 (
            .O(N__40049),
            .I(N__39987));
    ClkMux I__8512 (
            .O(N__40048),
            .I(N__39984));
    Span4Mux_v I__8511 (
            .O(N__40045),
            .I(N__39981));
    Span4Mux_v I__8510 (
            .O(N__40042),
            .I(N__39976));
    Span4Mux_h I__8509 (
            .O(N__40035),
            .I(N__39976));
    ClkMux I__8508 (
            .O(N__40034),
            .I(N__39973));
    LocalMux I__8507 (
            .O(N__40031),
            .I(N__39970));
    LocalMux I__8506 (
            .O(N__40028),
            .I(N__39967));
    Span4Mux_v I__8505 (
            .O(N__40025),
            .I(N__39962));
    Span4Mux_v I__8504 (
            .O(N__40018),
            .I(N__39962));
    Span4Mux_v I__8503 (
            .O(N__40015),
            .I(N__39957));
    Span4Mux_h I__8502 (
            .O(N__40010),
            .I(N__39957));
    Span4Mux_v I__8501 (
            .O(N__40007),
            .I(N__39946));
    Span4Mux_h I__8500 (
            .O(N__40004),
            .I(N__39946));
    LocalMux I__8499 (
            .O(N__40001),
            .I(N__39946));
    Span4Mux_v I__8498 (
            .O(N__39996),
            .I(N__39946));
    LocalMux I__8497 (
            .O(N__39993),
            .I(N__39946));
    Span4Mux_v I__8496 (
            .O(N__39990),
            .I(N__39939));
    LocalMux I__8495 (
            .O(N__39987),
            .I(N__39939));
    LocalMux I__8494 (
            .O(N__39984),
            .I(N__39939));
    Span4Mux_h I__8493 (
            .O(N__39981),
            .I(N__39932));
    Span4Mux_h I__8492 (
            .O(N__39976),
            .I(N__39932));
    LocalMux I__8491 (
            .O(N__39973),
            .I(N__39932));
    Span12Mux_s6_h I__8490 (
            .O(N__39970),
            .I(N__39929));
    Span4Mux_v I__8489 (
            .O(N__39967),
            .I(N__39926));
    Span4Mux_h I__8488 (
            .O(N__39962),
            .I(N__39923));
    Span4Mux_v I__8487 (
            .O(N__39957),
            .I(N__39918));
    Span4Mux_h I__8486 (
            .O(N__39946),
            .I(N__39918));
    Span4Mux_v I__8485 (
            .O(N__39939),
            .I(N__39915));
    Span4Mux_h I__8484 (
            .O(N__39932),
            .I(N__39912));
    Span12Mux_h I__8483 (
            .O(N__39929),
            .I(N__39909));
    Span4Mux_h I__8482 (
            .O(N__39926),
            .I(N__39904));
    Span4Mux_h I__8481 (
            .O(N__39923),
            .I(N__39904));
    Span4Mux_h I__8480 (
            .O(N__39918),
            .I(N__39899));
    Span4Mux_h I__8479 (
            .O(N__39915),
            .I(N__39899));
    Span4Mux_v I__8478 (
            .O(N__39912),
            .I(N__39896));
    Odrv12 I__8477 (
            .O(N__39909),
            .I(VDC_CLK));
    Odrv4 I__8476 (
            .O(N__39904),
            .I(VDC_CLK));
    Odrv4 I__8475 (
            .O(N__39899),
            .I(VDC_CLK));
    Odrv4 I__8474 (
            .O(N__39896),
            .I(VDC_CLK));
    InMux I__8473 (
            .O(N__39887),
            .I(N__39883));
    InMux I__8472 (
            .O(N__39886),
            .I(N__39880));
    LocalMux I__8471 (
            .O(N__39883),
            .I(secclk_cnt_15));
    LocalMux I__8470 (
            .O(N__39880),
            .I(secclk_cnt_15));
    InMux I__8469 (
            .O(N__39875),
            .I(n19523));
    InMux I__8468 (
            .O(N__39872),
            .I(N__39868));
    InMux I__8467 (
            .O(N__39871),
            .I(N__39865));
    LocalMux I__8466 (
            .O(N__39868),
            .I(secclk_cnt_16));
    LocalMux I__8465 (
            .O(N__39865),
            .I(secclk_cnt_16));
    InMux I__8464 (
            .O(N__39860),
            .I(bfn_14_20_0_));
    InMux I__8463 (
            .O(N__39857),
            .I(N__39853));
    InMux I__8462 (
            .O(N__39856),
            .I(N__39850));
    LocalMux I__8461 (
            .O(N__39853),
            .I(secclk_cnt_17));
    LocalMux I__8460 (
            .O(N__39850),
            .I(secclk_cnt_17));
    InMux I__8459 (
            .O(N__39845),
            .I(n19525));
    CascadeMux I__8458 (
            .O(N__39842),
            .I(N__39838));
    InMux I__8457 (
            .O(N__39841),
            .I(N__39835));
    InMux I__8456 (
            .O(N__39838),
            .I(N__39832));
    LocalMux I__8455 (
            .O(N__39835),
            .I(secclk_cnt_18));
    LocalMux I__8454 (
            .O(N__39832),
            .I(secclk_cnt_18));
    InMux I__8453 (
            .O(N__39827),
            .I(n19526));
    InMux I__8452 (
            .O(N__39824),
            .I(N__39820));
    InMux I__8451 (
            .O(N__39823),
            .I(N__39817));
    LocalMux I__8450 (
            .O(N__39820),
            .I(secclk_cnt_19));
    LocalMux I__8449 (
            .O(N__39817),
            .I(secclk_cnt_19));
    InMux I__8448 (
            .O(N__39812),
            .I(n19527));
    InMux I__8447 (
            .O(N__39809),
            .I(N__39805));
    InMux I__8446 (
            .O(N__39808),
            .I(N__39802));
    LocalMux I__8445 (
            .O(N__39805),
            .I(secclk_cnt_20));
    LocalMux I__8444 (
            .O(N__39802),
            .I(secclk_cnt_20));
    InMux I__8443 (
            .O(N__39797),
            .I(n19528));
    InMux I__8442 (
            .O(N__39794),
            .I(N__39790));
    InMux I__8441 (
            .O(N__39793),
            .I(N__39787));
    LocalMux I__8440 (
            .O(N__39790),
            .I(secclk_cnt_21));
    LocalMux I__8439 (
            .O(N__39787),
            .I(secclk_cnt_21));
    InMux I__8438 (
            .O(N__39782),
            .I(n19529));
    InMux I__8437 (
            .O(N__39779),
            .I(n19530));
    InMux I__8436 (
            .O(N__39776),
            .I(N__39772));
    InMux I__8435 (
            .O(N__39775),
            .I(N__39769));
    LocalMux I__8434 (
            .O(N__39772),
            .I(secclk_cnt_22));
    LocalMux I__8433 (
            .O(N__39769),
            .I(secclk_cnt_22));
    SRMux I__8432 (
            .O(N__39764),
            .I(N__39760));
    SRMux I__8431 (
            .O(N__39763),
            .I(N__39757));
    LocalMux I__8430 (
            .O(N__39760),
            .I(N__39753));
    LocalMux I__8429 (
            .O(N__39757),
            .I(N__39750));
    SRMux I__8428 (
            .O(N__39756),
            .I(N__39747));
    Span4Mux_h I__8427 (
            .O(N__39753),
            .I(N__39743));
    Span4Mux_h I__8426 (
            .O(N__39750),
            .I(N__39740));
    LocalMux I__8425 (
            .O(N__39747),
            .I(N__39737));
    InMux I__8424 (
            .O(N__39746),
            .I(N__39734));
    Odrv4 I__8423 (
            .O(N__39743),
            .I(n14731));
    Odrv4 I__8422 (
            .O(N__39740),
            .I(n14731));
    Odrv4 I__8421 (
            .O(N__39737),
            .I(n14731));
    LocalMux I__8420 (
            .O(N__39734),
            .I(n14731));
    InMux I__8419 (
            .O(N__39725),
            .I(N__39721));
    InMux I__8418 (
            .O(N__39724),
            .I(N__39718));
    LocalMux I__8417 (
            .O(N__39721),
            .I(secclk_cnt_7));
    LocalMux I__8416 (
            .O(N__39718),
            .I(secclk_cnt_7));
    InMux I__8415 (
            .O(N__39713),
            .I(n19515));
    InMux I__8414 (
            .O(N__39710),
            .I(N__39706));
    InMux I__8413 (
            .O(N__39709),
            .I(N__39703));
    LocalMux I__8412 (
            .O(N__39706),
            .I(secclk_cnt_8));
    LocalMux I__8411 (
            .O(N__39703),
            .I(secclk_cnt_8));
    InMux I__8410 (
            .O(N__39698),
            .I(bfn_14_19_0_));
    InMux I__8409 (
            .O(N__39695),
            .I(N__39691));
    InMux I__8408 (
            .O(N__39694),
            .I(N__39688));
    LocalMux I__8407 (
            .O(N__39691),
            .I(secclk_cnt_9));
    LocalMux I__8406 (
            .O(N__39688),
            .I(secclk_cnt_9));
    InMux I__8405 (
            .O(N__39683),
            .I(n19517));
    CascadeMux I__8404 (
            .O(N__39680),
            .I(N__39676));
    InMux I__8403 (
            .O(N__39679),
            .I(N__39673));
    InMux I__8402 (
            .O(N__39676),
            .I(N__39670));
    LocalMux I__8401 (
            .O(N__39673),
            .I(secclk_cnt_10));
    LocalMux I__8400 (
            .O(N__39670),
            .I(secclk_cnt_10));
    InMux I__8399 (
            .O(N__39665),
            .I(n19518));
    InMux I__8398 (
            .O(N__39662),
            .I(N__39658));
    InMux I__8397 (
            .O(N__39661),
            .I(N__39655));
    LocalMux I__8396 (
            .O(N__39658),
            .I(secclk_cnt_11));
    LocalMux I__8395 (
            .O(N__39655),
            .I(secclk_cnt_11));
    InMux I__8394 (
            .O(N__39650),
            .I(n19519));
    CascadeMux I__8393 (
            .O(N__39647),
            .I(N__39643));
    InMux I__8392 (
            .O(N__39646),
            .I(N__39640));
    InMux I__8391 (
            .O(N__39643),
            .I(N__39637));
    LocalMux I__8390 (
            .O(N__39640),
            .I(secclk_cnt_12));
    LocalMux I__8389 (
            .O(N__39637),
            .I(secclk_cnt_12));
    InMux I__8388 (
            .O(N__39632),
            .I(n19520));
    CascadeMux I__8387 (
            .O(N__39629),
            .I(N__39625));
    InMux I__8386 (
            .O(N__39628),
            .I(N__39622));
    InMux I__8385 (
            .O(N__39625),
            .I(N__39619));
    LocalMux I__8384 (
            .O(N__39622),
            .I(secclk_cnt_13));
    LocalMux I__8383 (
            .O(N__39619),
            .I(secclk_cnt_13));
    InMux I__8382 (
            .O(N__39614),
            .I(n19521));
    InMux I__8381 (
            .O(N__39611),
            .I(N__39607));
    InMux I__8380 (
            .O(N__39610),
            .I(N__39604));
    LocalMux I__8379 (
            .O(N__39607),
            .I(secclk_cnt_14));
    LocalMux I__8378 (
            .O(N__39604),
            .I(secclk_cnt_14));
    InMux I__8377 (
            .O(N__39599),
            .I(n19522));
    InMux I__8376 (
            .O(N__39596),
            .I(n19503));
    InMux I__8375 (
            .O(N__39593),
            .I(n19504));
    InMux I__8374 (
            .O(N__39590),
            .I(N__39586));
    InMux I__8373 (
            .O(N__39589),
            .I(N__39583));
    LocalMux I__8372 (
            .O(N__39586),
            .I(secclk_cnt_0));
    LocalMux I__8371 (
            .O(N__39583),
            .I(secclk_cnt_0));
    InMux I__8370 (
            .O(N__39578),
            .I(bfn_14_18_0_));
    CascadeMux I__8369 (
            .O(N__39575),
            .I(N__39571));
    InMux I__8368 (
            .O(N__39574),
            .I(N__39568));
    InMux I__8367 (
            .O(N__39571),
            .I(N__39565));
    LocalMux I__8366 (
            .O(N__39568),
            .I(secclk_cnt_1));
    LocalMux I__8365 (
            .O(N__39565),
            .I(secclk_cnt_1));
    InMux I__8364 (
            .O(N__39560),
            .I(n19509));
    InMux I__8363 (
            .O(N__39557),
            .I(N__39553));
    InMux I__8362 (
            .O(N__39556),
            .I(N__39550));
    LocalMux I__8361 (
            .O(N__39553),
            .I(secclk_cnt_2));
    LocalMux I__8360 (
            .O(N__39550),
            .I(secclk_cnt_2));
    InMux I__8359 (
            .O(N__39545),
            .I(n19510));
    InMux I__8358 (
            .O(N__39542),
            .I(N__39538));
    InMux I__8357 (
            .O(N__39541),
            .I(N__39535));
    LocalMux I__8356 (
            .O(N__39538),
            .I(secclk_cnt_3));
    LocalMux I__8355 (
            .O(N__39535),
            .I(secclk_cnt_3));
    InMux I__8354 (
            .O(N__39530),
            .I(n19511));
    InMux I__8353 (
            .O(N__39527),
            .I(N__39523));
    InMux I__8352 (
            .O(N__39526),
            .I(N__39520));
    LocalMux I__8351 (
            .O(N__39523),
            .I(secclk_cnt_4));
    LocalMux I__8350 (
            .O(N__39520),
            .I(secclk_cnt_4));
    InMux I__8349 (
            .O(N__39515),
            .I(n19512));
    InMux I__8348 (
            .O(N__39512),
            .I(N__39508));
    InMux I__8347 (
            .O(N__39511),
            .I(N__39505));
    LocalMux I__8346 (
            .O(N__39508),
            .I(secclk_cnt_5));
    LocalMux I__8345 (
            .O(N__39505),
            .I(secclk_cnt_5));
    InMux I__8344 (
            .O(N__39500),
            .I(n19513));
    InMux I__8343 (
            .O(N__39497),
            .I(N__39493));
    InMux I__8342 (
            .O(N__39496),
            .I(N__39490));
    LocalMux I__8341 (
            .O(N__39493),
            .I(secclk_cnt_6));
    LocalMux I__8340 (
            .O(N__39490),
            .I(secclk_cnt_6));
    InMux I__8339 (
            .O(N__39485),
            .I(n19514));
    InMux I__8338 (
            .O(N__39482),
            .I(N__39479));
    LocalMux I__8337 (
            .O(N__39479),
            .I(N__39476));
    Odrv12 I__8336 (
            .O(N__39476),
            .I(n10_adj_1613));
    InMux I__8335 (
            .O(N__39473),
            .I(bfn_14_17_0_));
    InMux I__8334 (
            .O(N__39470),
            .I(n19498));
    InMux I__8333 (
            .O(N__39467),
            .I(n19499));
    InMux I__8332 (
            .O(N__39464),
            .I(n19500));
    InMux I__8331 (
            .O(N__39461),
            .I(n19501));
    InMux I__8330 (
            .O(N__39458),
            .I(n19502));
    InMux I__8329 (
            .O(N__39455),
            .I(N__39452));
    LocalMux I__8328 (
            .O(N__39452),
            .I(n10));
    CascadeMux I__8327 (
            .O(N__39449),
            .I(N__39446));
    InMux I__8326 (
            .O(N__39446),
            .I(N__39443));
    LocalMux I__8325 (
            .O(N__39443),
            .I(N__39439));
    InMux I__8324 (
            .O(N__39442),
            .I(N__39436));
    Odrv4 I__8323 (
            .O(N__39439),
            .I(n8_adj_1565));
    LocalMux I__8322 (
            .O(N__39436),
            .I(n8_adj_1565));
    InMux I__8321 (
            .O(N__39431),
            .I(N__39428));
    LocalMux I__8320 (
            .O(N__39428),
            .I(N__39424));
    InMux I__8319 (
            .O(N__39427),
            .I(N__39421));
    Span4Mux_h I__8318 (
            .O(N__39424),
            .I(N__39418));
    LocalMux I__8317 (
            .O(N__39421),
            .I(n7_adj_1564));
    Odrv4 I__8316 (
            .O(N__39418),
            .I(n7_adj_1564));
    CascadeMux I__8315 (
            .O(N__39413),
            .I(N__39410));
    CascadeBuf I__8314 (
            .O(N__39410),
            .I(N__39407));
    CascadeMux I__8313 (
            .O(N__39407),
            .I(N__39404));
    CascadeBuf I__8312 (
            .O(N__39404),
            .I(N__39401));
    CascadeMux I__8311 (
            .O(N__39401),
            .I(N__39398));
    CascadeBuf I__8310 (
            .O(N__39398),
            .I(N__39395));
    CascadeMux I__8309 (
            .O(N__39395),
            .I(N__39392));
    CascadeBuf I__8308 (
            .O(N__39392),
            .I(N__39389));
    CascadeMux I__8307 (
            .O(N__39389),
            .I(N__39386));
    CascadeBuf I__8306 (
            .O(N__39386),
            .I(N__39383));
    CascadeMux I__8305 (
            .O(N__39383),
            .I(N__39380));
    CascadeBuf I__8304 (
            .O(N__39380),
            .I(N__39377));
    CascadeMux I__8303 (
            .O(N__39377),
            .I(N__39374));
    CascadeBuf I__8302 (
            .O(N__39374),
            .I(N__39371));
    CascadeMux I__8301 (
            .O(N__39371),
            .I(N__39368));
    CascadeBuf I__8300 (
            .O(N__39368),
            .I(N__39364));
    CascadeMux I__8299 (
            .O(N__39367),
            .I(N__39361));
    CascadeMux I__8298 (
            .O(N__39364),
            .I(N__39358));
    CascadeBuf I__8297 (
            .O(N__39361),
            .I(N__39355));
    CascadeBuf I__8296 (
            .O(N__39358),
            .I(N__39352));
    CascadeMux I__8295 (
            .O(N__39355),
            .I(N__39349));
    CascadeMux I__8294 (
            .O(N__39352),
            .I(N__39346));
    InMux I__8293 (
            .O(N__39349),
            .I(N__39343));
    InMux I__8292 (
            .O(N__39346),
            .I(N__39340));
    LocalMux I__8291 (
            .O(N__39343),
            .I(N__39337));
    LocalMux I__8290 (
            .O(N__39340),
            .I(N__39334));
    Span12Mux_s10_h I__8289 (
            .O(N__39337),
            .I(N__39331));
    Span4Mux_v I__8288 (
            .O(N__39334),
            .I(N__39328));
    Span12Mux_v I__8287 (
            .O(N__39331),
            .I(N__39325));
    Span4Mux_h I__8286 (
            .O(N__39328),
            .I(N__39322));
    Odrv12 I__8285 (
            .O(N__39325),
            .I(data_index_9_N_216_2));
    Odrv4 I__8284 (
            .O(N__39322),
            .I(data_index_9_N_216_2));
    InMux I__8283 (
            .O(N__39317),
            .I(N__39314));
    LocalMux I__8282 (
            .O(N__39314),
            .I(N__39310));
    InMux I__8281 (
            .O(N__39313),
            .I(N__39307));
    Span4Mux_v I__8280 (
            .O(N__39310),
            .I(N__39304));
    LocalMux I__8279 (
            .O(N__39307),
            .I(N__39301));
    Span4Mux_h I__8278 (
            .O(N__39304),
            .I(N__39298));
    Span4Mux_v I__8277 (
            .O(N__39301),
            .I(N__39295));
    Span4Mux_v I__8276 (
            .O(N__39298),
            .I(N__39292));
    Span4Mux_h I__8275 (
            .O(N__39295),
            .I(N__39289));
    Odrv4 I__8274 (
            .O(N__39292),
            .I(n14_adj_1573));
    Odrv4 I__8273 (
            .O(N__39289),
            .I(n14_adj_1573));
    InMux I__8272 (
            .O(N__39284),
            .I(N__39281));
    LocalMux I__8271 (
            .O(N__39281),
            .I(N__39278));
    Span4Mux_h I__8270 (
            .O(N__39278),
            .I(N__39275));
    Span4Mux_h I__8269 (
            .O(N__39275),
            .I(N__39271));
    InMux I__8268 (
            .O(N__39274),
            .I(N__39268));
    Sp12to4 I__8267 (
            .O(N__39271),
            .I(N__39263));
    LocalMux I__8266 (
            .O(N__39268),
            .I(N__39263));
    Span12Mux_v I__8265 (
            .O(N__39263),
            .I(N__39260));
    Odrv12 I__8264 (
            .O(N__39260),
            .I(n14_adj_1572));
    InMux I__8263 (
            .O(N__39257),
            .I(N__39254));
    LocalMux I__8262 (
            .O(N__39254),
            .I(N__39250));
    InMux I__8261 (
            .O(N__39253),
            .I(N__39247));
    Span4Mux_h I__8260 (
            .O(N__39250),
            .I(N__39244));
    LocalMux I__8259 (
            .O(N__39247),
            .I(acadc_skipcnt_7));
    Odrv4 I__8258 (
            .O(N__39244),
            .I(acadc_skipcnt_7));
    InMux I__8257 (
            .O(N__39239),
            .I(N__39236));
    LocalMux I__8256 (
            .O(N__39236),
            .I(N__39232));
    InMux I__8255 (
            .O(N__39235),
            .I(N__39229));
    Span4Mux_h I__8254 (
            .O(N__39232),
            .I(N__39226));
    LocalMux I__8253 (
            .O(N__39229),
            .I(acadc_skipcnt_2));
    Odrv4 I__8252 (
            .O(N__39226),
            .I(acadc_skipcnt_2));
    InMux I__8251 (
            .O(N__39221),
            .I(N__39218));
    LocalMux I__8250 (
            .O(N__39218),
            .I(n22_adj_1620));
    CascadeMux I__8249 (
            .O(N__39215),
            .I(N__39212));
    InMux I__8248 (
            .O(N__39212),
            .I(N__39209));
    LocalMux I__8247 (
            .O(N__39209),
            .I(N__39206));
    Span4Mux_h I__8246 (
            .O(N__39206),
            .I(N__39203));
    Odrv4 I__8245 (
            .O(N__39203),
            .I(n9_adj_1415));
    CascadeMux I__8244 (
            .O(N__39200),
            .I(N__39197));
    InMux I__8243 (
            .O(N__39197),
            .I(N__39194));
    LocalMux I__8242 (
            .O(N__39194),
            .I(N__39191));
    Span4Mux_h I__8241 (
            .O(N__39191),
            .I(N__39187));
    InMux I__8240 (
            .O(N__39190),
            .I(N__39184));
    Span4Mux_v I__8239 (
            .O(N__39187),
            .I(N__39179));
    LocalMux I__8238 (
            .O(N__39184),
            .I(N__39179));
    Span4Mux_v I__8237 (
            .O(N__39179),
            .I(N__39176));
    Span4Mux_h I__8236 (
            .O(N__39176),
            .I(N__39173));
    Odrv4 I__8235 (
            .O(N__39173),
            .I(n14_adj_1570));
    InMux I__8234 (
            .O(N__39170),
            .I(N__39167));
    LocalMux I__8233 (
            .O(N__39167),
            .I(N__39164));
    Span12Mux_v I__8232 (
            .O(N__39164),
            .I(N__39161));
    Odrv12 I__8231 (
            .O(N__39161),
            .I(n21048));
    CascadeMux I__8230 (
            .O(N__39158),
            .I(N__39154));
    InMux I__8229 (
            .O(N__39157),
            .I(N__39150));
    InMux I__8228 (
            .O(N__39154),
            .I(N__39147));
    CascadeMux I__8227 (
            .O(N__39153),
            .I(N__39144));
    LocalMux I__8226 (
            .O(N__39150),
            .I(N__39133));
    LocalMux I__8225 (
            .O(N__39147),
            .I(N__39130));
    InMux I__8224 (
            .O(N__39144),
            .I(N__39127));
    CascadeMux I__8223 (
            .O(N__39143),
            .I(N__39124));
    CascadeMux I__8222 (
            .O(N__39142),
            .I(N__39121));
    CascadeMux I__8221 (
            .O(N__39141),
            .I(N__39118));
    CascadeMux I__8220 (
            .O(N__39140),
            .I(N__39115));
    CascadeMux I__8219 (
            .O(N__39139),
            .I(N__39112));
    CascadeMux I__8218 (
            .O(N__39138),
            .I(N__39109));
    CascadeMux I__8217 (
            .O(N__39137),
            .I(N__39106));
    CascadeMux I__8216 (
            .O(N__39136),
            .I(N__39103));
    Span4Mux_h I__8215 (
            .O(N__39133),
            .I(N__39100));
    Span4Mux_v I__8214 (
            .O(N__39130),
            .I(N__39097));
    LocalMux I__8213 (
            .O(N__39127),
            .I(N__39094));
    InMux I__8212 (
            .O(N__39124),
            .I(N__39085));
    InMux I__8211 (
            .O(N__39121),
            .I(N__39085));
    InMux I__8210 (
            .O(N__39118),
            .I(N__39085));
    InMux I__8209 (
            .O(N__39115),
            .I(N__39085));
    InMux I__8208 (
            .O(N__39112),
            .I(N__39076));
    InMux I__8207 (
            .O(N__39109),
            .I(N__39076));
    InMux I__8206 (
            .O(N__39106),
            .I(N__39076));
    InMux I__8205 (
            .O(N__39103),
            .I(N__39076));
    Odrv4 I__8204 (
            .O(N__39100),
            .I(n10614));
    Odrv4 I__8203 (
            .O(N__39097),
            .I(n10614));
    Odrv12 I__8202 (
            .O(N__39094),
            .I(n10614));
    LocalMux I__8201 (
            .O(N__39085),
            .I(n10614));
    LocalMux I__8200 (
            .O(N__39076),
            .I(n10614));
    CEMux I__8199 (
            .O(N__39065),
            .I(N__39062));
    LocalMux I__8198 (
            .O(N__39062),
            .I(N__39058));
    CEMux I__8197 (
            .O(N__39061),
            .I(N__39055));
    Span4Mux_h I__8196 (
            .O(N__39058),
            .I(N__39052));
    LocalMux I__8195 (
            .O(N__39055),
            .I(N__39049));
    Span4Mux_v I__8194 (
            .O(N__39052),
            .I(N__39046));
    Span4Mux_h I__8193 (
            .O(N__39049),
            .I(N__39043));
    Sp12to4 I__8192 (
            .O(N__39046),
            .I(N__39040));
    Odrv4 I__8191 (
            .O(N__39043),
            .I(n12312));
    Odrv12 I__8190 (
            .O(N__39040),
            .I(n12312));
    IoInMux I__8189 (
            .O(N__39035),
            .I(N__39032));
    LocalMux I__8188 (
            .O(N__39032),
            .I(N__39029));
    IoSpan4Mux I__8187 (
            .O(N__39029),
            .I(N__39026));
    Span4Mux_s2_h I__8186 (
            .O(N__39026),
            .I(N__39023));
    Sp12to4 I__8185 (
            .O(N__39023),
            .I(N__39020));
    Span12Mux_h I__8184 (
            .O(N__39020),
            .I(N__39017));
    Span12Mux_v I__8183 (
            .O(N__39017),
            .I(N__39012));
    InMux I__8182 (
            .O(N__39016),
            .I(N__39009));
    InMux I__8181 (
            .O(N__39015),
            .I(N__39006));
    Odrv12 I__8180 (
            .O(N__39012),
            .I(VDC_RNG0));
    LocalMux I__8179 (
            .O(N__39009),
            .I(VDC_RNG0));
    LocalMux I__8178 (
            .O(N__39006),
            .I(VDC_RNG0));
    InMux I__8177 (
            .O(N__38999),
            .I(N__38996));
    LocalMux I__8176 (
            .O(N__38996),
            .I(N__38991));
    CascadeMux I__8175 (
            .O(N__38995),
            .I(N__38988));
    InMux I__8174 (
            .O(N__38994),
            .I(N__38985));
    Span4Mux_h I__8173 (
            .O(N__38991),
            .I(N__38982));
    InMux I__8172 (
            .O(N__38988),
            .I(N__38979));
    LocalMux I__8171 (
            .O(N__38985),
            .I(acadc_skipCount_12));
    Odrv4 I__8170 (
            .O(N__38982),
            .I(acadc_skipCount_12));
    LocalMux I__8169 (
            .O(N__38979),
            .I(acadc_skipCount_12));
    InMux I__8168 (
            .O(N__38972),
            .I(N__38969));
    LocalMux I__8167 (
            .O(N__38969),
            .I(N__38961));
    InMux I__8166 (
            .O(N__38968),
            .I(N__38958));
    InMux I__8165 (
            .O(N__38967),
            .I(N__38951));
    InMux I__8164 (
            .O(N__38966),
            .I(N__38947));
    InMux I__8163 (
            .O(N__38965),
            .I(N__38944));
    InMux I__8162 (
            .O(N__38964),
            .I(N__38941));
    Span4Mux_h I__8161 (
            .O(N__38961),
            .I(N__38936));
    LocalMux I__8160 (
            .O(N__38958),
            .I(N__38936));
    InMux I__8159 (
            .O(N__38957),
            .I(N__38925));
    InMux I__8158 (
            .O(N__38956),
            .I(N__38925));
    InMux I__8157 (
            .O(N__38955),
            .I(N__38925));
    InMux I__8156 (
            .O(N__38954),
            .I(N__38922));
    LocalMux I__8155 (
            .O(N__38951),
            .I(N__38919));
    InMux I__8154 (
            .O(N__38950),
            .I(N__38916));
    LocalMux I__8153 (
            .O(N__38947),
            .I(N__38913));
    LocalMux I__8152 (
            .O(N__38944),
            .I(N__38908));
    LocalMux I__8151 (
            .O(N__38941),
            .I(N__38908));
    Span4Mux_h I__8150 (
            .O(N__38936),
            .I(N__38905));
    InMux I__8149 (
            .O(N__38935),
            .I(N__38902));
    InMux I__8148 (
            .O(N__38934),
            .I(N__38897));
    InMux I__8147 (
            .O(N__38933),
            .I(N__38897));
    InMux I__8146 (
            .O(N__38932),
            .I(N__38894));
    LocalMux I__8145 (
            .O(N__38925),
            .I(N__38889));
    LocalMux I__8144 (
            .O(N__38922),
            .I(N__38889));
    Span4Mux_h I__8143 (
            .O(N__38919),
            .I(N__38886));
    LocalMux I__8142 (
            .O(N__38916),
            .I(N__38883));
    Span4Mux_h I__8141 (
            .O(N__38913),
            .I(N__38876));
    Span4Mux_v I__8140 (
            .O(N__38908),
            .I(N__38876));
    Span4Mux_h I__8139 (
            .O(N__38905),
            .I(N__38876));
    LocalMux I__8138 (
            .O(N__38902),
            .I(n12383));
    LocalMux I__8137 (
            .O(N__38897),
            .I(n12383));
    LocalMux I__8136 (
            .O(N__38894),
            .I(n12383));
    Odrv4 I__8135 (
            .O(N__38889),
            .I(n12383));
    Odrv4 I__8134 (
            .O(N__38886),
            .I(n12383));
    Odrv12 I__8133 (
            .O(N__38883),
            .I(n12383));
    Odrv4 I__8132 (
            .O(N__38876),
            .I(n12383));
    InMux I__8131 (
            .O(N__38861),
            .I(N__38858));
    LocalMux I__8130 (
            .O(N__38858),
            .I(N__38854));
    InMux I__8129 (
            .O(N__38857),
            .I(N__38851));
    Span4Mux_h I__8128 (
            .O(N__38854),
            .I(N__38848));
    LocalMux I__8127 (
            .O(N__38851),
            .I(acadc_skipcnt_13));
    Odrv4 I__8126 (
            .O(N__38848),
            .I(acadc_skipcnt_13));
    InMux I__8125 (
            .O(N__38843),
            .I(N__38840));
    LocalMux I__8124 (
            .O(N__38840),
            .I(N__38836));
    InMux I__8123 (
            .O(N__38839),
            .I(N__38832));
    Span4Mux_v I__8122 (
            .O(N__38836),
            .I(N__38829));
    InMux I__8121 (
            .O(N__38835),
            .I(N__38826));
    LocalMux I__8120 (
            .O(N__38832),
            .I(acadc_skipCount_13));
    Odrv4 I__8119 (
            .O(N__38829),
            .I(acadc_skipCount_13));
    LocalMux I__8118 (
            .O(N__38826),
            .I(acadc_skipCount_13));
    InMux I__8117 (
            .O(N__38819),
            .I(N__38816));
    LocalMux I__8116 (
            .O(N__38816),
            .I(n14));
    InMux I__8115 (
            .O(N__38813),
            .I(N__38810));
    LocalMux I__8114 (
            .O(N__38810),
            .I(N__38806));
    InMux I__8113 (
            .O(N__38809),
            .I(N__38803));
    Span4Mux_h I__8112 (
            .O(N__38806),
            .I(N__38800));
    LocalMux I__8111 (
            .O(N__38803),
            .I(acadc_skipcnt_1));
    Odrv4 I__8110 (
            .O(N__38800),
            .I(acadc_skipcnt_1));
    CascadeMux I__8109 (
            .O(N__38795),
            .I(N__38792));
    InMux I__8108 (
            .O(N__38792),
            .I(N__38789));
    LocalMux I__8107 (
            .O(N__38789),
            .I(N__38785));
    InMux I__8106 (
            .O(N__38788),
            .I(N__38782));
    Span4Mux_v I__8105 (
            .O(N__38785),
            .I(N__38779));
    LocalMux I__8104 (
            .O(N__38782),
            .I(acadc_skipcnt_4));
    Odrv4 I__8103 (
            .O(N__38779),
            .I(acadc_skipcnt_4));
    InMux I__8102 (
            .O(N__38774),
            .I(N__38771));
    LocalMux I__8101 (
            .O(N__38771),
            .I(n18_adj_1611));
    InMux I__8100 (
            .O(N__38768),
            .I(N__38764));
    InMux I__8099 (
            .O(N__38767),
            .I(N__38761));
    LocalMux I__8098 (
            .O(N__38764),
            .I(N__38756));
    LocalMux I__8097 (
            .O(N__38761),
            .I(N__38756));
    Span4Mux_v I__8096 (
            .O(N__38756),
            .I(N__38752));
    InMux I__8095 (
            .O(N__38755),
            .I(N__38749));
    Span4Mux_h I__8094 (
            .O(N__38752),
            .I(N__38746));
    LocalMux I__8093 (
            .O(N__38749),
            .I(data_index_4));
    Odrv4 I__8092 (
            .O(N__38746),
            .I(data_index_4));
    InMux I__8091 (
            .O(N__38741),
            .I(N__38735));
    InMux I__8090 (
            .O(N__38740),
            .I(N__38735));
    LocalMux I__8089 (
            .O(N__38735),
            .I(N__38732));
    Span4Mux_v I__8088 (
            .O(N__38732),
            .I(N__38729));
    Odrv4 I__8087 (
            .O(N__38729),
            .I(n7_adj_1560));
    CascadeMux I__8086 (
            .O(N__38726),
            .I(N__38722));
    InMux I__8085 (
            .O(N__38725),
            .I(N__38717));
    InMux I__8084 (
            .O(N__38722),
            .I(N__38717));
    LocalMux I__8083 (
            .O(N__38717),
            .I(n8_adj_1561));
    CascadeMux I__8082 (
            .O(N__38714),
            .I(N__38711));
    CascadeBuf I__8081 (
            .O(N__38711),
            .I(N__38708));
    CascadeMux I__8080 (
            .O(N__38708),
            .I(N__38705));
    CascadeBuf I__8079 (
            .O(N__38705),
            .I(N__38702));
    CascadeMux I__8078 (
            .O(N__38702),
            .I(N__38699));
    CascadeBuf I__8077 (
            .O(N__38699),
            .I(N__38696));
    CascadeMux I__8076 (
            .O(N__38696),
            .I(N__38693));
    CascadeBuf I__8075 (
            .O(N__38693),
            .I(N__38690));
    CascadeMux I__8074 (
            .O(N__38690),
            .I(N__38687));
    CascadeBuf I__8073 (
            .O(N__38687),
            .I(N__38684));
    CascadeMux I__8072 (
            .O(N__38684),
            .I(N__38681));
    CascadeBuf I__8071 (
            .O(N__38681),
            .I(N__38678));
    CascadeMux I__8070 (
            .O(N__38678),
            .I(N__38675));
    CascadeBuf I__8069 (
            .O(N__38675),
            .I(N__38672));
    CascadeMux I__8068 (
            .O(N__38672),
            .I(N__38669));
    CascadeBuf I__8067 (
            .O(N__38669),
            .I(N__38665));
    CascadeMux I__8066 (
            .O(N__38668),
            .I(N__38662));
    CascadeMux I__8065 (
            .O(N__38665),
            .I(N__38659));
    CascadeBuf I__8064 (
            .O(N__38662),
            .I(N__38656));
    CascadeBuf I__8063 (
            .O(N__38659),
            .I(N__38653));
    CascadeMux I__8062 (
            .O(N__38656),
            .I(N__38650));
    CascadeMux I__8061 (
            .O(N__38653),
            .I(N__38647));
    InMux I__8060 (
            .O(N__38650),
            .I(N__38644));
    InMux I__8059 (
            .O(N__38647),
            .I(N__38641));
    LocalMux I__8058 (
            .O(N__38644),
            .I(N__38638));
    LocalMux I__8057 (
            .O(N__38641),
            .I(N__38635));
    Span12Mux_s11_h I__8056 (
            .O(N__38638),
            .I(N__38632));
    Span4Mux_v I__8055 (
            .O(N__38635),
            .I(N__38629));
    Span12Mux_v I__8054 (
            .O(N__38632),
            .I(N__38626));
    Span4Mux_h I__8053 (
            .O(N__38629),
            .I(N__38623));
    Odrv12 I__8052 (
            .O(N__38626),
            .I(data_index_9_N_216_4));
    Odrv4 I__8051 (
            .O(N__38623),
            .I(data_index_9_N_216_4));
    InMux I__8050 (
            .O(N__38618),
            .I(N__38615));
    LocalMux I__8049 (
            .O(N__38615),
            .I(n22013));
    CascadeMux I__8048 (
            .O(N__38612),
            .I(n12441_cascade_));
    CascadeMux I__8047 (
            .O(N__38609),
            .I(n8_adj_1567_cascade_));
    InMux I__8046 (
            .O(N__38606),
            .I(N__38602));
    InMux I__8045 (
            .O(N__38605),
            .I(N__38599));
    LocalMux I__8044 (
            .O(N__38602),
            .I(N__38594));
    LocalMux I__8043 (
            .O(N__38599),
            .I(N__38594));
    Span4Mux_v I__8042 (
            .O(N__38594),
            .I(N__38590));
    InMux I__8041 (
            .O(N__38593),
            .I(N__38587));
    Span4Mux_h I__8040 (
            .O(N__38590),
            .I(N__38584));
    LocalMux I__8039 (
            .O(N__38587),
            .I(data_index_1));
    Odrv4 I__8038 (
            .O(N__38584),
            .I(data_index_1));
    CascadeMux I__8037 (
            .O(N__38579),
            .I(N__38575));
    InMux I__8036 (
            .O(N__38578),
            .I(N__38568));
    InMux I__8035 (
            .O(N__38575),
            .I(N__38564));
    InMux I__8034 (
            .O(N__38574),
            .I(N__38552));
    InMux I__8033 (
            .O(N__38573),
            .I(N__38549));
    InMux I__8032 (
            .O(N__38572),
            .I(N__38544));
    InMux I__8031 (
            .O(N__38571),
            .I(N__38544));
    LocalMux I__8030 (
            .O(N__38568),
            .I(N__38541));
    InMux I__8029 (
            .O(N__38567),
            .I(N__38538));
    LocalMux I__8028 (
            .O(N__38564),
            .I(N__38535));
    InMux I__8027 (
            .O(N__38563),
            .I(N__38532));
    InMux I__8026 (
            .O(N__38562),
            .I(N__38529));
    InMux I__8025 (
            .O(N__38561),
            .I(N__38524));
    InMux I__8024 (
            .O(N__38560),
            .I(N__38524));
    InMux I__8023 (
            .O(N__38559),
            .I(N__38521));
    InMux I__8022 (
            .O(N__38558),
            .I(N__38516));
    InMux I__8021 (
            .O(N__38557),
            .I(N__38516));
    InMux I__8020 (
            .O(N__38556),
            .I(N__38511));
    InMux I__8019 (
            .O(N__38555),
            .I(N__38511));
    LocalMux I__8018 (
            .O(N__38552),
            .I(N__38502));
    LocalMux I__8017 (
            .O(N__38549),
            .I(N__38502));
    LocalMux I__8016 (
            .O(N__38544),
            .I(N__38502));
    Span4Mux_h I__8015 (
            .O(N__38541),
            .I(N__38502));
    LocalMux I__8014 (
            .O(N__38538),
            .I(N__38497));
    Span4Mux_v I__8013 (
            .O(N__38535),
            .I(N__38497));
    LocalMux I__8012 (
            .O(N__38532),
            .I(n11835));
    LocalMux I__8011 (
            .O(N__38529),
            .I(n11835));
    LocalMux I__8010 (
            .O(N__38524),
            .I(n11835));
    LocalMux I__8009 (
            .O(N__38521),
            .I(n11835));
    LocalMux I__8008 (
            .O(N__38516),
            .I(n11835));
    LocalMux I__8007 (
            .O(N__38511),
            .I(n11835));
    Odrv4 I__8006 (
            .O(N__38502),
            .I(n11835));
    Odrv4 I__8005 (
            .O(N__38497),
            .I(n11835));
    InMux I__8004 (
            .O(N__38480),
            .I(N__38476));
    InMux I__8003 (
            .O(N__38479),
            .I(N__38473));
    LocalMux I__8002 (
            .O(N__38476),
            .I(N__38467));
    LocalMux I__8001 (
            .O(N__38473),
            .I(N__38464));
    InMux I__8000 (
            .O(N__38472),
            .I(N__38461));
    InMux I__7999 (
            .O(N__38471),
            .I(N__38456));
    InMux I__7998 (
            .O(N__38470),
            .I(N__38456));
    Span4Mux_h I__7997 (
            .O(N__38467),
            .I(N__38445));
    Span4Mux_h I__7996 (
            .O(N__38464),
            .I(N__38440));
    LocalMux I__7995 (
            .O(N__38461),
            .I(N__38440));
    LocalMux I__7994 (
            .O(N__38456),
            .I(N__38437));
    InMux I__7993 (
            .O(N__38455),
            .I(N__38434));
    InMux I__7992 (
            .O(N__38454),
            .I(N__38431));
    InMux I__7991 (
            .O(N__38453),
            .I(N__38426));
    InMux I__7990 (
            .O(N__38452),
            .I(N__38426));
    InMux I__7989 (
            .O(N__38451),
            .I(N__38423));
    InMux I__7988 (
            .O(N__38450),
            .I(N__38416));
    InMux I__7987 (
            .O(N__38449),
            .I(N__38416));
    InMux I__7986 (
            .O(N__38448),
            .I(N__38416));
    Odrv4 I__7985 (
            .O(N__38445),
            .I(n16763));
    Odrv4 I__7984 (
            .O(N__38440),
            .I(n16763));
    Odrv12 I__7983 (
            .O(N__38437),
            .I(n16763));
    LocalMux I__7982 (
            .O(N__38434),
            .I(n16763));
    LocalMux I__7981 (
            .O(N__38431),
            .I(n16763));
    LocalMux I__7980 (
            .O(N__38426),
            .I(n16763));
    LocalMux I__7979 (
            .O(N__38423),
            .I(n16763));
    LocalMux I__7978 (
            .O(N__38416),
            .I(n16763));
    InMux I__7977 (
            .O(N__38399),
            .I(N__38395));
    InMux I__7976 (
            .O(N__38398),
            .I(N__38392));
    LocalMux I__7975 (
            .O(N__38395),
            .I(N__38389));
    LocalMux I__7974 (
            .O(N__38392),
            .I(N__38385));
    Span4Mux_h I__7973 (
            .O(N__38389),
            .I(N__38382));
    InMux I__7972 (
            .O(N__38388),
            .I(N__38379));
    Span12Mux_h I__7971 (
            .O(N__38385),
            .I(N__38376));
    Span4Mux_h I__7970 (
            .O(N__38382),
            .I(N__38373));
    LocalMux I__7969 (
            .O(N__38379),
            .I(buf_dds1_1));
    Odrv12 I__7968 (
            .O(N__38376),
            .I(buf_dds1_1));
    Odrv4 I__7967 (
            .O(N__38373),
            .I(buf_dds1_1));
    InMux I__7966 (
            .O(N__38366),
            .I(N__38363));
    LocalMux I__7965 (
            .O(N__38363),
            .I(N__38360));
    Span4Mux_h I__7964 (
            .O(N__38360),
            .I(N__38356));
    InMux I__7963 (
            .O(N__38359),
            .I(N__38353));
    Span4Mux_h I__7962 (
            .O(N__38356),
            .I(N__38347));
    LocalMux I__7961 (
            .O(N__38353),
            .I(N__38347));
    InMux I__7960 (
            .O(N__38352),
            .I(N__38344));
    Span4Mux_h I__7959 (
            .O(N__38347),
            .I(N__38341));
    LocalMux I__7958 (
            .O(N__38344),
            .I(buf_adcdata_iac_14));
    Odrv4 I__7957 (
            .O(N__38341),
            .I(buf_adcdata_iac_14));
    InMux I__7956 (
            .O(N__38336),
            .I(N__38333));
    LocalMux I__7955 (
            .O(N__38333),
            .I(N__38330));
    Span4Mux_h I__7954 (
            .O(N__38330),
            .I(N__38327));
    Odrv4 I__7953 (
            .O(N__38327),
            .I(n16));
    InMux I__7952 (
            .O(N__38324),
            .I(N__38321));
    LocalMux I__7951 (
            .O(N__38321),
            .I(N__38318));
    Odrv12 I__7950 (
            .O(N__38318),
            .I(n20953));
    InMux I__7949 (
            .O(N__38315),
            .I(N__38312));
    LocalMux I__7948 (
            .O(N__38312),
            .I(N__38308));
    InMux I__7947 (
            .O(N__38311),
            .I(N__38305));
    Odrv12 I__7946 (
            .O(N__38308),
            .I(buf_readRTD_3));
    LocalMux I__7945 (
            .O(N__38305),
            .I(buf_readRTD_3));
    InMux I__7944 (
            .O(N__38300),
            .I(N__38297));
    LocalMux I__7943 (
            .O(N__38297),
            .I(n20879));
    InMux I__7942 (
            .O(N__38294),
            .I(N__38291));
    LocalMux I__7941 (
            .O(N__38291),
            .I(N__38287));
    CascadeMux I__7940 (
            .O(N__38290),
            .I(N__38283));
    Span4Mux_h I__7939 (
            .O(N__38287),
            .I(N__38280));
    InMux I__7938 (
            .O(N__38286),
            .I(N__38277));
    InMux I__7937 (
            .O(N__38283),
            .I(N__38274));
    Span4Mux_h I__7936 (
            .O(N__38280),
            .I(N__38271));
    LocalMux I__7935 (
            .O(N__38277),
            .I(N__38268));
    LocalMux I__7934 (
            .O(N__38274),
            .I(N__38263));
    Span4Mux_v I__7933 (
            .O(N__38271),
            .I(N__38263));
    Odrv4 I__7932 (
            .O(N__38268),
            .I(buf_adcdata_vac_11));
    Odrv4 I__7931 (
            .O(N__38263),
            .I(buf_adcdata_vac_11));
    InMux I__7930 (
            .O(N__38258),
            .I(N__38255));
    LocalMux I__7929 (
            .O(N__38255),
            .I(N__38252));
    Span4Mux_v I__7928 (
            .O(N__38252),
            .I(N__38249));
    Span4Mux_h I__7927 (
            .O(N__38249),
            .I(N__38245));
    InMux I__7926 (
            .O(N__38248),
            .I(N__38242));
    Odrv4 I__7925 (
            .O(N__38245),
            .I(buf_adcdata_vdc_11));
    LocalMux I__7924 (
            .O(N__38242),
            .I(buf_adcdata_vdc_11));
    InMux I__7923 (
            .O(N__38237),
            .I(N__38234));
    LocalMux I__7922 (
            .O(N__38234),
            .I(n19_adj_1513));
    CascadeMux I__7921 (
            .O(N__38231),
            .I(n22178_cascade_));
    CascadeMux I__7920 (
            .O(N__38228),
            .I(n22181_cascade_));
    CascadeMux I__7919 (
            .O(N__38225),
            .I(n30_adj_1511_cascade_));
    InMux I__7918 (
            .O(N__38222),
            .I(N__38219));
    LocalMux I__7917 (
            .O(N__38219),
            .I(N__38215));
    CascadeMux I__7916 (
            .O(N__38218),
            .I(N__38212));
    Span4Mux_v I__7915 (
            .O(N__38215),
            .I(N__38209));
    InMux I__7914 (
            .O(N__38212),
            .I(N__38206));
    Sp12to4 I__7913 (
            .O(N__38209),
            .I(N__38203));
    LocalMux I__7912 (
            .O(N__38206),
            .I(data_idxvec_4));
    Odrv12 I__7911 (
            .O(N__38203),
            .I(data_idxvec_4));
    InMux I__7910 (
            .O(N__38198),
            .I(N__38195));
    LocalMux I__7909 (
            .O(N__38195),
            .I(n26_adj_1510));
    InMux I__7908 (
            .O(N__38192),
            .I(N__38189));
    LocalMux I__7907 (
            .O(N__38189),
            .I(n19_adj_1509));
    InMux I__7906 (
            .O(N__38186),
            .I(N__38183));
    LocalMux I__7905 (
            .O(N__38183),
            .I(N__38179));
    CascadeMux I__7904 (
            .O(N__38182),
            .I(N__38176));
    Sp12to4 I__7903 (
            .O(N__38179),
            .I(N__38173));
    InMux I__7902 (
            .O(N__38176),
            .I(N__38170));
    Odrv12 I__7901 (
            .O(N__38173),
            .I(buf_readRTD_4));
    LocalMux I__7900 (
            .O(N__38170),
            .I(buf_readRTD_4));
    InMux I__7899 (
            .O(N__38165),
            .I(N__38162));
    LocalMux I__7898 (
            .O(N__38162),
            .I(N__38158));
    InMux I__7897 (
            .O(N__38161),
            .I(N__38155));
    Span4Mux_h I__7896 (
            .O(N__38158),
            .I(N__38152));
    LocalMux I__7895 (
            .O(N__38155),
            .I(N__38149));
    Span4Mux_h I__7894 (
            .O(N__38152),
            .I(N__38145));
    Span4Mux_v I__7893 (
            .O(N__38149),
            .I(N__38142));
    InMux I__7892 (
            .O(N__38148),
            .I(N__38139));
    Span4Mux_h I__7891 (
            .O(N__38145),
            .I(N__38136));
    Span4Mux_h I__7890 (
            .O(N__38142),
            .I(N__38133));
    LocalMux I__7889 (
            .O(N__38139),
            .I(buf_adcdata_iac_12));
    Odrv4 I__7888 (
            .O(N__38136),
            .I(buf_adcdata_iac_12));
    Odrv4 I__7887 (
            .O(N__38133),
            .I(buf_adcdata_iac_12));
    CascadeMux I__7886 (
            .O(N__38126),
            .I(n22010_cascade_));
    InMux I__7885 (
            .O(N__38123),
            .I(N__38120));
    LocalMux I__7884 (
            .O(N__38120),
            .I(N__38117));
    Span4Mux_h I__7883 (
            .O(N__38117),
            .I(N__38114));
    Span4Mux_h I__7882 (
            .O(N__38114),
            .I(N__38111));
    Odrv4 I__7881 (
            .O(N__38111),
            .I(n16_adj_1508));
    InMux I__7880 (
            .O(N__38108),
            .I(N__38105));
    LocalMux I__7879 (
            .O(N__38105),
            .I(N__38102));
    Span4Mux_v I__7878 (
            .O(N__38102),
            .I(N__38098));
    CascadeMux I__7877 (
            .O(N__38101),
            .I(N__38095));
    Span4Mux_h I__7876 (
            .O(N__38098),
            .I(N__38092));
    InMux I__7875 (
            .O(N__38095),
            .I(N__38089));
    Odrv4 I__7874 (
            .O(N__38092),
            .I(buf_adcdata_vdc_14));
    LocalMux I__7873 (
            .O(N__38089),
            .I(buf_adcdata_vdc_14));
    InMux I__7872 (
            .O(N__38084),
            .I(N__38081));
    LocalMux I__7871 (
            .O(N__38081),
            .I(N__38078));
    Span4Mux_h I__7870 (
            .O(N__38078),
            .I(N__38073));
    CascadeMux I__7869 (
            .O(N__38077),
            .I(N__38070));
    InMux I__7868 (
            .O(N__38076),
            .I(N__38067));
    Span4Mux_v I__7867 (
            .O(N__38073),
            .I(N__38064));
    InMux I__7866 (
            .O(N__38070),
            .I(N__38061));
    LocalMux I__7865 (
            .O(N__38067),
            .I(N__38056));
    Span4Mux_h I__7864 (
            .O(N__38064),
            .I(N__38056));
    LocalMux I__7863 (
            .O(N__38061),
            .I(buf_adcdata_vac_14));
    Odrv4 I__7862 (
            .O(N__38056),
            .I(buf_adcdata_vac_14));
    InMux I__7861 (
            .O(N__38051),
            .I(N__38048));
    LocalMux I__7860 (
            .O(N__38048),
            .I(N__38045));
    Span12Mux_h I__7859 (
            .O(N__38045),
            .I(N__38041));
    InMux I__7858 (
            .O(N__38044),
            .I(N__38038));
    Odrv12 I__7857 (
            .O(N__38041),
            .I(buf_readRTD_6));
    LocalMux I__7856 (
            .O(N__38038),
            .I(buf_readRTD_6));
    CascadeMux I__7855 (
            .O(N__38033),
            .I(n19_cascade_));
    InMux I__7854 (
            .O(N__38030),
            .I(N__38027));
    LocalMux I__7853 (
            .O(N__38027),
            .I(N__38024));
    Odrv4 I__7852 (
            .O(N__38024),
            .I(n20954));
    CascadeMux I__7851 (
            .O(N__38021),
            .I(N__38018));
    InMux I__7850 (
            .O(N__38018),
            .I(N__38015));
    LocalMux I__7849 (
            .O(N__38015),
            .I(N__38010));
    InMux I__7848 (
            .O(N__38014),
            .I(N__38007));
    InMux I__7847 (
            .O(N__38013),
            .I(N__38004));
    Span4Mux_v I__7846 (
            .O(N__38010),
            .I(N__38001));
    LocalMux I__7845 (
            .O(N__38007),
            .I(N__37998));
    LocalMux I__7844 (
            .O(N__38004),
            .I(acadc_skipCount_6));
    Odrv4 I__7843 (
            .O(N__38001),
            .I(acadc_skipCount_6));
    Odrv12 I__7842 (
            .O(N__37998),
            .I(acadc_skipCount_6));
    InMux I__7841 (
            .O(N__37991),
            .I(N__37988));
    LocalMux I__7840 (
            .O(N__37988),
            .I(n20929));
    CascadeMux I__7839 (
            .O(N__37985),
            .I(N__37982));
    InMux I__7838 (
            .O(N__37982),
            .I(N__37978));
    InMux I__7837 (
            .O(N__37981),
            .I(N__37975));
    LocalMux I__7836 (
            .O(N__37978),
            .I(N__37972));
    LocalMux I__7835 (
            .O(N__37975),
            .I(N__37966));
    Span4Mux_h I__7834 (
            .O(N__37972),
            .I(N__37963));
    InMux I__7833 (
            .O(N__37971),
            .I(N__37958));
    InMux I__7832 (
            .O(N__37970),
            .I(N__37958));
    InMux I__7831 (
            .O(N__37969),
            .I(N__37955));
    Span4Mux_h I__7830 (
            .O(N__37966),
            .I(N__37952));
    Span4Mux_h I__7829 (
            .O(N__37963),
            .I(N__37947));
    LocalMux I__7828 (
            .O(N__37958),
            .I(N__37947));
    LocalMux I__7827 (
            .O(N__37955),
            .I(N__37944));
    Span4Mux_h I__7826 (
            .O(N__37952),
            .I(N__37941));
    Span4Mux_v I__7825 (
            .O(N__37947),
            .I(N__37938));
    Odrv4 I__7824 (
            .O(N__37944),
            .I(comm_buf_1_3));
    Odrv4 I__7823 (
            .O(N__37941),
            .I(comm_buf_1_3));
    Odrv4 I__7822 (
            .O(N__37938),
            .I(comm_buf_1_3));
    InMux I__7821 (
            .O(N__37931),
            .I(N__37926));
    CascadeMux I__7820 (
            .O(N__37930),
            .I(N__37923));
    CascadeMux I__7819 (
            .O(N__37929),
            .I(N__37920));
    LocalMux I__7818 (
            .O(N__37926),
            .I(N__37917));
    InMux I__7817 (
            .O(N__37923),
            .I(N__37912));
    InMux I__7816 (
            .O(N__37920),
            .I(N__37912));
    Odrv4 I__7815 (
            .O(N__37917),
            .I(acadc_skipCount_3));
    LocalMux I__7814 (
            .O(N__37912),
            .I(acadc_skipCount_3));
    CascadeMux I__7813 (
            .O(N__37907),
            .I(n20884_cascade_));
    InMux I__7812 (
            .O(N__37904),
            .I(N__37901));
    LocalMux I__7811 (
            .O(N__37901),
            .I(N__37898));
    Span4Mux_h I__7810 (
            .O(N__37898),
            .I(N__37895));
    Span4Mux_h I__7809 (
            .O(N__37895),
            .I(N__37892));
    Odrv4 I__7808 (
            .O(N__37892),
            .I(n20878));
    CascadeMux I__7807 (
            .O(N__37889),
            .I(n22124_cascade_));
    InMux I__7806 (
            .O(N__37886),
            .I(N__37883));
    LocalMux I__7805 (
            .O(N__37883),
            .I(n22127));
    CascadeMux I__7804 (
            .O(N__37880),
            .I(N__37877));
    InMux I__7803 (
            .O(N__37877),
            .I(N__37873));
    InMux I__7802 (
            .O(N__37876),
            .I(N__37870));
    LocalMux I__7801 (
            .O(N__37873),
            .I(N__37865));
    LocalMux I__7800 (
            .O(N__37870),
            .I(N__37865));
    Odrv4 I__7799 (
            .O(N__37865),
            .I(data_idxvec_3));
    InMux I__7798 (
            .O(N__37862),
            .I(N__37859));
    LocalMux I__7797 (
            .O(N__37859),
            .I(N__37856));
    Span4Mux_v I__7796 (
            .O(N__37856),
            .I(N__37853));
    Span4Mux_h I__7795 (
            .O(N__37853),
            .I(N__37850));
    Span4Mux_h I__7794 (
            .O(N__37850),
            .I(N__37847));
    Span4Mux_h I__7793 (
            .O(N__37847),
            .I(N__37844));
    Odrv4 I__7792 (
            .O(N__37844),
            .I(buf_data_iac_11));
    CascadeMux I__7791 (
            .O(N__37841),
            .I(n26_adj_1514_cascade_));
    InMux I__7790 (
            .O(N__37838),
            .I(N__37835));
    LocalMux I__7789 (
            .O(N__37835),
            .I(n20885));
    InMux I__7788 (
            .O(N__37832),
            .I(N__37829));
    LocalMux I__7787 (
            .O(N__37829),
            .I(N__37826));
    Odrv12 I__7786 (
            .O(N__37826),
            .I(comm_buf_3_3));
    InMux I__7785 (
            .O(N__37823),
            .I(N__37820));
    LocalMux I__7784 (
            .O(N__37820),
            .I(N__37817));
    Span4Mux_h I__7783 (
            .O(N__37817),
            .I(N__37814));
    Sp12to4 I__7782 (
            .O(N__37814),
            .I(N__37811));
    Odrv12 I__7781 (
            .O(N__37811),
            .I(comm_buf_2_3));
    InMux I__7780 (
            .O(N__37808),
            .I(N__37805));
    LocalMux I__7779 (
            .O(N__37805),
            .I(n2_adj_1590));
    CascadeMux I__7778 (
            .O(N__37802),
            .I(n21102_cascade_));
    InMux I__7777 (
            .O(N__37799),
            .I(N__37796));
    LocalMux I__7776 (
            .O(N__37796),
            .I(n21_adj_1618));
    InMux I__7775 (
            .O(N__37793),
            .I(N__37790));
    LocalMux I__7774 (
            .O(N__37790),
            .I(n16_adj_1599));
    InMux I__7773 (
            .O(N__37787),
            .I(N__37783));
    CascadeMux I__7772 (
            .O(N__37786),
            .I(N__37780));
    LocalMux I__7771 (
            .O(N__37783),
            .I(N__37777));
    InMux I__7770 (
            .O(N__37780),
            .I(N__37774));
    Span4Mux_h I__7769 (
            .O(N__37777),
            .I(N__37771));
    LocalMux I__7768 (
            .O(N__37774),
            .I(data_idxvec_6));
    Odrv4 I__7767 (
            .O(N__37771),
            .I(data_idxvec_6));
    InMux I__7766 (
            .O(N__37766),
            .I(N__37763));
    LocalMux I__7765 (
            .O(N__37763),
            .I(N__37760));
    Span4Mux_h I__7764 (
            .O(N__37760),
            .I(N__37757));
    Span4Mux_h I__7763 (
            .O(N__37757),
            .I(N__37754));
    Odrv4 I__7762 (
            .O(N__37754),
            .I(buf_data_iac_14));
    CascadeMux I__7761 (
            .O(N__37751),
            .I(n26_adj_1505_cascade_));
    CascadeMux I__7760 (
            .O(N__37748),
            .I(n20930_cascade_));
    CascadeMux I__7759 (
            .O(N__37745),
            .I(n21962_cascade_));
    CascadeMux I__7758 (
            .O(N__37742),
            .I(n21965_cascade_));
    InMux I__7757 (
            .O(N__37739),
            .I(N__37736));
    LocalMux I__7756 (
            .O(N__37736),
            .I(N__37733));
    Span4Mux_h I__7755 (
            .O(N__37733),
            .I(N__37730));
    Span4Mux_v I__7754 (
            .O(N__37730),
            .I(N__37727));
    Span4Mux_v I__7753 (
            .O(N__37727),
            .I(N__37724));
    Odrv4 I__7752 (
            .O(N__37724),
            .I(buf_data_vac_12));
    InMux I__7751 (
            .O(N__37721),
            .I(N__37718));
    LocalMux I__7750 (
            .O(N__37718),
            .I(N__37715));
    Span4Mux_h I__7749 (
            .O(N__37715),
            .I(N__37712));
    Odrv4 I__7748 (
            .O(N__37712),
            .I(comm_buf_4_4));
    InMux I__7747 (
            .O(N__37709),
            .I(N__37706));
    LocalMux I__7746 (
            .O(N__37706),
            .I(N__37703));
    Span4Mux_v I__7745 (
            .O(N__37703),
            .I(N__37700));
    Span4Mux_v I__7744 (
            .O(N__37700),
            .I(N__37697));
    Span4Mux_h I__7743 (
            .O(N__37697),
            .I(N__37694));
    Span4Mux_h I__7742 (
            .O(N__37694),
            .I(N__37691));
    Odrv4 I__7741 (
            .O(N__37691),
            .I(buf_data_vac_11));
    InMux I__7740 (
            .O(N__37688),
            .I(N__37685));
    LocalMux I__7739 (
            .O(N__37685),
            .I(N__37682));
    Span4Mux_h I__7738 (
            .O(N__37682),
            .I(N__37679));
    Span4Mux_h I__7737 (
            .O(N__37679),
            .I(N__37676));
    Span4Mux_v I__7736 (
            .O(N__37676),
            .I(N__37673));
    Span4Mux_v I__7735 (
            .O(N__37673),
            .I(N__37670));
    Odrv4 I__7734 (
            .O(N__37670),
            .I(buf_data_vac_10));
    InMux I__7733 (
            .O(N__37667),
            .I(N__37664));
    LocalMux I__7732 (
            .O(N__37664),
            .I(N__37661));
    Span4Mux_h I__7731 (
            .O(N__37661),
            .I(N__37658));
    Span4Mux_h I__7730 (
            .O(N__37658),
            .I(N__37655));
    Span4Mux_v I__7729 (
            .O(N__37655),
            .I(N__37652));
    Span4Mux_v I__7728 (
            .O(N__37652),
            .I(N__37649));
    Odrv4 I__7727 (
            .O(N__37649),
            .I(buf_data_vac_9));
    CEMux I__7726 (
            .O(N__37646),
            .I(N__37643));
    LocalMux I__7725 (
            .O(N__37643),
            .I(N__37640));
    Span4Mux_h I__7724 (
            .O(N__37640),
            .I(N__37637));
    Odrv4 I__7723 (
            .O(N__37637),
            .I(n12194));
    SRMux I__7722 (
            .O(N__37634),
            .I(N__37631));
    LocalMux I__7721 (
            .O(N__37631),
            .I(N__37628));
    Span4Mux_h I__7720 (
            .O(N__37628),
            .I(N__37625));
    Odrv4 I__7719 (
            .O(N__37625),
            .I(n14794));
    CascadeMux I__7718 (
            .O(N__37622),
            .I(n1_adj_1589_cascade_));
    InMux I__7717 (
            .O(N__37619),
            .I(N__37615));
    InMux I__7716 (
            .O(N__37618),
            .I(N__37612));
    LocalMux I__7715 (
            .O(N__37615),
            .I(N__37609));
    LocalMux I__7714 (
            .O(N__37612),
            .I(comm_buf_6_3));
    Odrv4 I__7713 (
            .O(N__37609),
            .I(comm_buf_6_3));
    CascadeMux I__7712 (
            .O(N__37604),
            .I(n21296_cascade_));
    InMux I__7711 (
            .O(N__37601),
            .I(N__37598));
    LocalMux I__7710 (
            .O(N__37598),
            .I(n22154));
    InMux I__7709 (
            .O(N__37595),
            .I(N__37592));
    LocalMux I__7708 (
            .O(N__37592),
            .I(comm_buf_4_3));
    InMux I__7707 (
            .O(N__37589),
            .I(N__37586));
    LocalMux I__7706 (
            .O(N__37586),
            .I(N__37583));
    Span4Mux_v I__7705 (
            .O(N__37583),
            .I(N__37580));
    Odrv4 I__7704 (
            .O(N__37580),
            .I(comm_buf_5_3));
    InMux I__7703 (
            .O(N__37577),
            .I(N__37574));
    LocalMux I__7702 (
            .O(N__37574),
            .I(n4_adj_1591));
    CascadeMux I__7701 (
            .O(N__37571),
            .I(N__37568));
    InMux I__7700 (
            .O(N__37568),
            .I(N__37565));
    LocalMux I__7699 (
            .O(N__37565),
            .I(comm_buf_2_0));
    InMux I__7698 (
            .O(N__37562),
            .I(N__37559));
    LocalMux I__7697 (
            .O(N__37559),
            .I(N__37556));
    Odrv12 I__7696 (
            .O(N__37556),
            .I(comm_buf_3_0));
    InMux I__7695 (
            .O(N__37553),
            .I(N__37550));
    LocalMux I__7694 (
            .O(N__37550),
            .I(n2));
    InMux I__7693 (
            .O(N__37547),
            .I(N__37544));
    LocalMux I__7692 (
            .O(N__37544),
            .I(N__37541));
    Span4Mux_v I__7691 (
            .O(N__37541),
            .I(N__37538));
    Odrv4 I__7690 (
            .O(N__37538),
            .I(comm_buf_5_0));
    InMux I__7689 (
            .O(N__37535),
            .I(N__37532));
    LocalMux I__7688 (
            .O(N__37532),
            .I(n20970));
    CascadeMux I__7687 (
            .O(N__37529),
            .I(n4_adj_1507_cascade_));
    InMux I__7686 (
            .O(N__37526),
            .I(N__37523));
    LocalMux I__7685 (
            .O(N__37523),
            .I(n21980));
    CascadeMux I__7684 (
            .O(N__37520),
            .I(n21116_cascade_));
    InMux I__7683 (
            .O(N__37517),
            .I(N__37513));
    InMux I__7682 (
            .O(N__37516),
            .I(N__37509));
    LocalMux I__7681 (
            .O(N__37513),
            .I(N__37506));
    InMux I__7680 (
            .O(N__37512),
            .I(N__37503));
    LocalMux I__7679 (
            .O(N__37509),
            .I(N__37500));
    Span4Mux_h I__7678 (
            .O(N__37506),
            .I(N__37495));
    LocalMux I__7677 (
            .O(N__37503),
            .I(N__37495));
    Span12Mux_h I__7676 (
            .O(N__37500),
            .I(N__37492));
    Span4Mux_v I__7675 (
            .O(N__37495),
            .I(N__37489));
    Span12Mux_v I__7674 (
            .O(N__37492),
            .I(N__37486));
    Span4Mux_v I__7673 (
            .O(N__37489),
            .I(N__37483));
    Odrv12 I__7672 (
            .O(N__37486),
            .I(n10713));
    Odrv4 I__7671 (
            .O(N__37483),
            .I(n10713));
    InMux I__7670 (
            .O(N__37478),
            .I(N__37475));
    LocalMux I__7669 (
            .O(N__37475),
            .I(n12_adj_1602));
    InMux I__7668 (
            .O(N__37472),
            .I(N__37469));
    LocalMux I__7667 (
            .O(N__37469),
            .I(N__37466));
    Span12Mux_h I__7666 (
            .O(N__37466),
            .I(N__37463));
    Span12Mux_v I__7665 (
            .O(N__37463),
            .I(N__37460));
    Odrv12 I__7664 (
            .O(N__37460),
            .I(buf_data_vac_8));
    InMux I__7663 (
            .O(N__37457),
            .I(N__37454));
    LocalMux I__7662 (
            .O(N__37454),
            .I(comm_buf_4_0));
    InMux I__7661 (
            .O(N__37451),
            .I(N__37448));
    LocalMux I__7660 (
            .O(N__37448),
            .I(N__37445));
    Span4Mux_h I__7659 (
            .O(N__37445),
            .I(N__37442));
    Span4Mux_h I__7658 (
            .O(N__37442),
            .I(N__37439));
    Span4Mux_v I__7657 (
            .O(N__37439),
            .I(N__37436));
    Odrv4 I__7656 (
            .O(N__37436),
            .I(buf_data_vac_15));
    InMux I__7655 (
            .O(N__37433),
            .I(N__37430));
    LocalMux I__7654 (
            .O(N__37430),
            .I(N__37427));
    Span12Mux_h I__7653 (
            .O(N__37427),
            .I(N__37424));
    Odrv12 I__7652 (
            .O(N__37424),
            .I(buf_data_vac_14));
    InMux I__7651 (
            .O(N__37421),
            .I(N__37418));
    LocalMux I__7650 (
            .O(N__37418),
            .I(N__37415));
    Span4Mux_h I__7649 (
            .O(N__37415),
            .I(N__37412));
    Span4Mux_v I__7648 (
            .O(N__37412),
            .I(N__37409));
    Span4Mux_h I__7647 (
            .O(N__37409),
            .I(N__37406));
    Odrv4 I__7646 (
            .O(N__37406),
            .I(buf_data_vac_13));
    InMux I__7645 (
            .O(N__37403),
            .I(N__37400));
    LocalMux I__7644 (
            .O(N__37400),
            .I(N__37397));
    Span4Mux_v I__7643 (
            .O(N__37397),
            .I(N__37394));
    Span4Mux_h I__7642 (
            .O(N__37394),
            .I(N__37391));
    Span4Mux_h I__7641 (
            .O(N__37391),
            .I(N__37388));
    Odrv4 I__7640 (
            .O(N__37388),
            .I(buf_data_vac_23));
    InMux I__7639 (
            .O(N__37385),
            .I(N__37382));
    LocalMux I__7638 (
            .O(N__37382),
            .I(N__37379));
    Span4Mux_v I__7637 (
            .O(N__37379),
            .I(N__37376));
    Span4Mux_h I__7636 (
            .O(N__37376),
            .I(N__37373));
    Odrv4 I__7635 (
            .O(N__37373),
            .I(buf_data_vac_22));
    InMux I__7634 (
            .O(N__37370),
            .I(N__37367));
    LocalMux I__7633 (
            .O(N__37367),
            .I(N__37364));
    Span4Mux_h I__7632 (
            .O(N__37364),
            .I(N__37361));
    Span4Mux_h I__7631 (
            .O(N__37361),
            .I(N__37358));
    Odrv4 I__7630 (
            .O(N__37358),
            .I(buf_data_vac_21));
    InMux I__7629 (
            .O(N__37355),
            .I(N__37352));
    LocalMux I__7628 (
            .O(N__37352),
            .I(N__37349));
    Span4Mux_h I__7627 (
            .O(N__37349),
            .I(N__37346));
    Span4Mux_h I__7626 (
            .O(N__37346),
            .I(N__37343));
    Odrv4 I__7625 (
            .O(N__37343),
            .I(buf_data_vac_19));
    InMux I__7624 (
            .O(N__37340),
            .I(N__37337));
    LocalMux I__7623 (
            .O(N__37337),
            .I(N__37334));
    Span4Mux_h I__7622 (
            .O(N__37334),
            .I(N__37331));
    Span4Mux_v I__7621 (
            .O(N__37331),
            .I(N__37328));
    Span4Mux_h I__7620 (
            .O(N__37328),
            .I(N__37325));
    Odrv4 I__7619 (
            .O(N__37325),
            .I(buf_data_vac_18));
    InMux I__7618 (
            .O(N__37322),
            .I(N__37319));
    LocalMux I__7617 (
            .O(N__37319),
            .I(N__37316));
    Span4Mux_h I__7616 (
            .O(N__37316),
            .I(N__37313));
    Span4Mux_v I__7615 (
            .O(N__37313),
            .I(N__37310));
    Span4Mux_h I__7614 (
            .O(N__37310),
            .I(N__37307));
    Odrv4 I__7613 (
            .O(N__37307),
            .I(buf_data_vac_17));
    CEMux I__7612 (
            .O(N__37304),
            .I(N__37301));
    LocalMux I__7611 (
            .O(N__37301),
            .I(N__37298));
    Span4Mux_v I__7610 (
            .O(N__37298),
            .I(N__37295));
    Odrv4 I__7609 (
            .O(N__37295),
            .I(n12152));
    SRMux I__7608 (
            .O(N__37292),
            .I(N__37289));
    LocalMux I__7607 (
            .O(N__37289),
            .I(n14787));
    CascadeMux I__7606 (
            .O(N__37286),
            .I(n1_cascade_));
    CascadeMux I__7605 (
            .O(N__37283),
            .I(n30_adj_1535_cascade_));
    CascadeMux I__7604 (
            .O(N__37280),
            .I(N__37277));
    InMux I__7603 (
            .O(N__37277),
            .I(N__37273));
    InMux I__7602 (
            .O(N__37276),
            .I(N__37270));
    LocalMux I__7601 (
            .O(N__37273),
            .I(\ADC_VDC.genclk.t0on_6 ));
    LocalMux I__7600 (
            .O(N__37270),
            .I(\ADC_VDC.genclk.t0on_6 ));
    InMux I__7599 (
            .O(N__37265),
            .I(N__37261));
    InMux I__7598 (
            .O(N__37264),
            .I(N__37258));
    LocalMux I__7597 (
            .O(N__37261),
            .I(\ADC_VDC.genclk.t0on_1 ));
    LocalMux I__7596 (
            .O(N__37258),
            .I(\ADC_VDC.genclk.t0on_1 ));
    CascadeMux I__7595 (
            .O(N__37253),
            .I(N__37249));
    CascadeMux I__7594 (
            .O(N__37252),
            .I(N__37246));
    InMux I__7593 (
            .O(N__37249),
            .I(N__37243));
    InMux I__7592 (
            .O(N__37246),
            .I(N__37240));
    LocalMux I__7591 (
            .O(N__37243),
            .I(N__37237));
    LocalMux I__7590 (
            .O(N__37240),
            .I(\ADC_VDC.genclk.t0on_4 ));
    Odrv4 I__7589 (
            .O(N__37237),
            .I(\ADC_VDC.genclk.t0on_4 ));
    InMux I__7588 (
            .O(N__37232),
            .I(N__37228));
    InMux I__7587 (
            .O(N__37231),
            .I(N__37225));
    LocalMux I__7586 (
            .O(N__37228),
            .I(\ADC_VDC.genclk.t0on_0 ));
    LocalMux I__7585 (
            .O(N__37225),
            .I(\ADC_VDC.genclk.t0on_0 ));
    CascadeMux I__7584 (
            .O(N__37220),
            .I(\ADC_VDC.genclk.n21211_cascade_ ));
    CascadeMux I__7583 (
            .O(N__37217),
            .I(N__37213));
    InMux I__7582 (
            .O(N__37216),
            .I(N__37210));
    InMux I__7581 (
            .O(N__37213),
            .I(N__37207));
    LocalMux I__7580 (
            .O(N__37210),
            .I(N__37202));
    LocalMux I__7579 (
            .O(N__37207),
            .I(N__37202));
    Odrv4 I__7578 (
            .O(N__37202),
            .I(\ADC_VDC.genclk.n21205 ));
    InMux I__7577 (
            .O(N__37199),
            .I(N__37195));
    InMux I__7576 (
            .O(N__37198),
            .I(N__37192));
    LocalMux I__7575 (
            .O(N__37195),
            .I(\ADC_VDC.genclk.t0on_13 ));
    LocalMux I__7574 (
            .O(N__37192),
            .I(\ADC_VDC.genclk.t0on_13 ));
    InMux I__7573 (
            .O(N__37187),
            .I(N__37183));
    InMux I__7572 (
            .O(N__37186),
            .I(N__37180));
    LocalMux I__7571 (
            .O(N__37183),
            .I(\ADC_VDC.genclk.t0on_3 ));
    LocalMux I__7570 (
            .O(N__37180),
            .I(\ADC_VDC.genclk.t0on_3 ));
    CascadeMux I__7569 (
            .O(N__37175),
            .I(N__37171));
    InMux I__7568 (
            .O(N__37174),
            .I(N__37168));
    InMux I__7567 (
            .O(N__37171),
            .I(N__37165));
    LocalMux I__7566 (
            .O(N__37168),
            .I(\ADC_VDC.genclk.t0on_5 ));
    LocalMux I__7565 (
            .O(N__37165),
            .I(\ADC_VDC.genclk.t0on_5 ));
    CascadeMux I__7564 (
            .O(N__37160),
            .I(N__37157));
    InMux I__7563 (
            .O(N__37157),
            .I(N__37153));
    InMux I__7562 (
            .O(N__37156),
            .I(N__37150));
    LocalMux I__7561 (
            .O(N__37153),
            .I(\ADC_VDC.genclk.t0on_8 ));
    LocalMux I__7560 (
            .O(N__37150),
            .I(\ADC_VDC.genclk.t0on_8 ));
    InMux I__7559 (
            .O(N__37145),
            .I(N__37142));
    LocalMux I__7558 (
            .O(N__37142),
            .I(\ADC_VDC.genclk.n26_adj_1408 ));
    CascadeMux I__7557 (
            .O(N__37139),
            .I(N__37136));
    InMux I__7556 (
            .O(N__37136),
            .I(N__37132));
    InMux I__7555 (
            .O(N__37135),
            .I(N__37129));
    LocalMux I__7554 (
            .O(N__37132),
            .I(\ADC_VDC.genclk.t0on_14 ));
    LocalMux I__7553 (
            .O(N__37129),
            .I(\ADC_VDC.genclk.t0on_14 ));
    InMux I__7552 (
            .O(N__37124),
            .I(N__37120));
    InMux I__7551 (
            .O(N__37123),
            .I(N__37117));
    LocalMux I__7550 (
            .O(N__37120),
            .I(\ADC_VDC.genclk.t0on_9 ));
    LocalMux I__7549 (
            .O(N__37117),
            .I(\ADC_VDC.genclk.t0on_9 ));
    CascadeMux I__7548 (
            .O(N__37112),
            .I(N__37108));
    InMux I__7547 (
            .O(N__37111),
            .I(N__37105));
    InMux I__7546 (
            .O(N__37108),
            .I(N__37102));
    LocalMux I__7545 (
            .O(N__37105),
            .I(\ADC_VDC.genclk.t0on_15 ));
    LocalMux I__7544 (
            .O(N__37102),
            .I(\ADC_VDC.genclk.t0on_15 ));
    InMux I__7543 (
            .O(N__37097),
            .I(N__37093));
    InMux I__7542 (
            .O(N__37096),
            .I(N__37090));
    LocalMux I__7541 (
            .O(N__37093),
            .I(\ADC_VDC.genclk.t0on_11 ));
    LocalMux I__7540 (
            .O(N__37090),
            .I(\ADC_VDC.genclk.t0on_11 ));
    InMux I__7539 (
            .O(N__37085),
            .I(N__37082));
    LocalMux I__7538 (
            .O(N__37082),
            .I(\ADC_VDC.genclk.n28_adj_1407 ));
    CascadeMux I__7537 (
            .O(N__37079),
            .I(N__37076));
    InMux I__7536 (
            .O(N__37076),
            .I(N__37072));
    InMux I__7535 (
            .O(N__37075),
            .I(N__37069));
    LocalMux I__7534 (
            .O(N__37072),
            .I(\ADC_VDC.genclk.t0on_12 ));
    LocalMux I__7533 (
            .O(N__37069),
            .I(\ADC_VDC.genclk.t0on_12 ));
    CascadeMux I__7532 (
            .O(N__37064),
            .I(N__37061));
    InMux I__7531 (
            .O(N__37061),
            .I(N__37057));
    InMux I__7530 (
            .O(N__37060),
            .I(N__37054));
    LocalMux I__7529 (
            .O(N__37057),
            .I(\ADC_VDC.genclk.t0on_2 ));
    LocalMux I__7528 (
            .O(N__37054),
            .I(\ADC_VDC.genclk.t0on_2 ));
    CascadeMux I__7527 (
            .O(N__37049),
            .I(N__37045));
    InMux I__7526 (
            .O(N__37048),
            .I(N__37042));
    InMux I__7525 (
            .O(N__37045),
            .I(N__37039));
    LocalMux I__7524 (
            .O(N__37042),
            .I(\ADC_VDC.genclk.t0on_7 ));
    LocalMux I__7523 (
            .O(N__37039),
            .I(\ADC_VDC.genclk.t0on_7 ));
    CascadeMux I__7522 (
            .O(N__37034),
            .I(N__37031));
    InMux I__7521 (
            .O(N__37031),
            .I(N__37027));
    InMux I__7520 (
            .O(N__37030),
            .I(N__37024));
    LocalMux I__7519 (
            .O(N__37027),
            .I(\ADC_VDC.genclk.t0on_10 ));
    LocalMux I__7518 (
            .O(N__37024),
            .I(\ADC_VDC.genclk.t0on_10 ));
    InMux I__7517 (
            .O(N__37019),
            .I(N__37016));
    LocalMux I__7516 (
            .O(N__37016),
            .I(\ADC_VDC.genclk.n27_adj_1409 ));
    InMux I__7515 (
            .O(N__37013),
            .I(N__37010));
    LocalMux I__7514 (
            .O(N__37010),
            .I(N__37007));
    Span12Mux_h I__7513 (
            .O(N__37007),
            .I(N__37004));
    Odrv12 I__7512 (
            .O(N__37004),
            .I(buf_data_vac_16));
    InMux I__7511 (
            .O(N__37001),
            .I(N__36998));
    LocalMux I__7510 (
            .O(N__36998),
            .I(N__36995));
    Span4Mux_v I__7509 (
            .O(N__36995),
            .I(N__36992));
    Span4Mux_h I__7508 (
            .O(N__36992),
            .I(N__36989));
    Odrv4 I__7507 (
            .O(N__36989),
            .I(buf_data_vac_20));
    InMux I__7506 (
            .O(N__36986),
            .I(N__36983));
    LocalMux I__7505 (
            .O(N__36983),
            .I(N__36980));
    Odrv12 I__7504 (
            .O(N__36980),
            .I(comm_buf_3_4));
    InMux I__7503 (
            .O(N__36977),
            .I(N__36974));
    LocalMux I__7502 (
            .O(N__36974),
            .I(n28_adj_1621));
    InMux I__7501 (
            .O(N__36971),
            .I(N__36968));
    LocalMux I__7500 (
            .O(N__36968),
            .I(n14_adj_1592));
    InMux I__7499 (
            .O(N__36965),
            .I(N__36961));
    CascadeMux I__7498 (
            .O(N__36964),
            .I(N__36958));
    LocalMux I__7497 (
            .O(N__36961),
            .I(N__36955));
    InMux I__7496 (
            .O(N__36958),
            .I(N__36951));
    Span4Mux_v I__7495 (
            .O(N__36955),
            .I(N__36948));
    CascadeMux I__7494 (
            .O(N__36954),
            .I(N__36945));
    LocalMux I__7493 (
            .O(N__36951),
            .I(N__36942));
    Span4Mux_v I__7492 (
            .O(N__36948),
            .I(N__36939));
    InMux I__7491 (
            .O(N__36945),
            .I(N__36936));
    Span4Mux_h I__7490 (
            .O(N__36942),
            .I(N__36931));
    Span4Mux_h I__7489 (
            .O(N__36939),
            .I(N__36931));
    LocalMux I__7488 (
            .O(N__36936),
            .I(buf_dds1_14));
    Odrv4 I__7487 (
            .O(N__36931),
            .I(buf_dds1_14));
    CascadeMux I__7486 (
            .O(N__36926),
            .I(N__36922));
    CascadeMux I__7485 (
            .O(N__36925),
            .I(N__36919));
    InMux I__7484 (
            .O(N__36922),
            .I(N__36916));
    InMux I__7483 (
            .O(N__36919),
            .I(N__36913));
    LocalMux I__7482 (
            .O(N__36916),
            .I(N__36910));
    LocalMux I__7481 (
            .O(N__36913),
            .I(N__36906));
    Span4Mux_h I__7480 (
            .O(N__36910),
            .I(N__36903));
    InMux I__7479 (
            .O(N__36909),
            .I(N__36900));
    Span4Mux_v I__7478 (
            .O(N__36906),
            .I(N__36897));
    Span4Mux_v I__7477 (
            .O(N__36903),
            .I(N__36894));
    LocalMux I__7476 (
            .O(N__36900),
            .I(buf_dds0_14));
    Odrv4 I__7475 (
            .O(N__36897),
            .I(buf_dds0_14));
    Odrv4 I__7474 (
            .O(N__36894),
            .I(buf_dds0_14));
    CascadeMux I__7473 (
            .O(N__36887),
            .I(n22115_cascade_));
    InMux I__7472 (
            .O(N__36884),
            .I(N__36881));
    LocalMux I__7471 (
            .O(N__36881),
            .I(N__36878));
    Span4Mux_h I__7470 (
            .O(N__36878),
            .I(N__36875));
    Span4Mux_v I__7469 (
            .O(N__36875),
            .I(N__36872));
    Odrv4 I__7468 (
            .O(N__36872),
            .I(n22163));
    IoInMux I__7467 (
            .O(N__36869),
            .I(N__36866));
    LocalMux I__7466 (
            .O(N__36866),
            .I(N__36862));
    InMux I__7465 (
            .O(N__36865),
            .I(N__36859));
    Span4Mux_s0_h I__7464 (
            .O(N__36862),
            .I(N__36856));
    LocalMux I__7463 (
            .O(N__36859),
            .I(N__36853));
    Sp12to4 I__7462 (
            .O(N__36856),
            .I(N__36850));
    Span4Mux_h I__7461 (
            .O(N__36853),
            .I(N__36847));
    Span12Mux_v I__7460 (
            .O(N__36850),
            .I(N__36844));
    Span4Mux_v I__7459 (
            .O(N__36847),
            .I(N__36840));
    Span12Mux_h I__7458 (
            .O(N__36844),
            .I(N__36837));
    InMux I__7457 (
            .O(N__36843),
            .I(N__36834));
    Span4Mux_h I__7456 (
            .O(N__36840),
            .I(N__36831));
    Odrv12 I__7455 (
            .O(N__36837),
            .I(VAC_FLT0));
    LocalMux I__7454 (
            .O(N__36834),
            .I(VAC_FLT0));
    Odrv4 I__7453 (
            .O(N__36831),
            .I(VAC_FLT0));
    CascadeMux I__7452 (
            .O(N__36824),
            .I(N__36821));
    InMux I__7451 (
            .O(N__36821),
            .I(N__36817));
    InMux I__7450 (
            .O(N__36820),
            .I(N__36814));
    LocalMux I__7449 (
            .O(N__36817),
            .I(N__36811));
    LocalMux I__7448 (
            .O(N__36814),
            .I(N__36808));
    Span4Mux_h I__7447 (
            .O(N__36811),
            .I(N__36805));
    Span4Mux_v I__7446 (
            .O(N__36808),
            .I(N__36802));
    Span4Mux_v I__7445 (
            .O(N__36805),
            .I(N__36799));
    Span4Mux_v I__7444 (
            .O(N__36802),
            .I(N__36796));
    Sp12to4 I__7443 (
            .O(N__36799),
            .I(N__36790));
    Sp12to4 I__7442 (
            .O(N__36796),
            .I(N__36790));
    InMux I__7441 (
            .O(N__36795),
            .I(N__36787));
    Span12Mux_h I__7440 (
            .O(N__36790),
            .I(N__36784));
    LocalMux I__7439 (
            .O(N__36787),
            .I(buf_adcdata_iac_22));
    Odrv12 I__7438 (
            .O(N__36784),
            .I(buf_adcdata_iac_22));
    InMux I__7437 (
            .O(N__36779),
            .I(N__36776));
    LocalMux I__7436 (
            .O(N__36776),
            .I(n22112));
    CascadeMux I__7435 (
            .O(N__36773),
            .I(N__36770));
    InMux I__7434 (
            .O(N__36770),
            .I(N__36767));
    LocalMux I__7433 (
            .O(N__36767),
            .I(N__36764));
    Span4Mux_v I__7432 (
            .O(N__36764),
            .I(N__36761));
    Span4Mux_v I__7431 (
            .O(N__36761),
            .I(N__36758));
    Span4Mux_v I__7430 (
            .O(N__36758),
            .I(N__36755));
    Odrv4 I__7429 (
            .O(N__36755),
            .I(n21037));
    InMux I__7428 (
            .O(N__36752),
            .I(N__36749));
    LocalMux I__7427 (
            .O(N__36749),
            .I(N__36746));
    Span4Mux_h I__7426 (
            .O(N__36746),
            .I(N__36743));
    Span4Mux_v I__7425 (
            .O(N__36743),
            .I(N__36740));
    Odrv4 I__7424 (
            .O(N__36740),
            .I(n23_adj_1534));
    CascadeMux I__7423 (
            .O(N__36737),
            .I(n22070_cascade_));
    InMux I__7422 (
            .O(N__36734),
            .I(N__36731));
    LocalMux I__7421 (
            .O(N__36731),
            .I(n20856));
    CascadeMux I__7420 (
            .O(N__36728),
            .I(n22073_cascade_));
    CascadeMux I__7419 (
            .O(N__36725),
            .I(N__36721));
    InMux I__7418 (
            .O(N__36724),
            .I(N__36710));
    InMux I__7417 (
            .O(N__36721),
            .I(N__36710));
    InMux I__7416 (
            .O(N__36720),
            .I(N__36702));
    InMux I__7415 (
            .O(N__36719),
            .I(N__36702));
    InMux I__7414 (
            .O(N__36718),
            .I(N__36693));
    InMux I__7413 (
            .O(N__36717),
            .I(N__36693));
    InMux I__7412 (
            .O(N__36716),
            .I(N__36693));
    InMux I__7411 (
            .O(N__36715),
            .I(N__36693));
    LocalMux I__7410 (
            .O(N__36710),
            .I(N__36690));
    InMux I__7409 (
            .O(N__36709),
            .I(N__36687));
    InMux I__7408 (
            .O(N__36708),
            .I(N__36680));
    InMux I__7407 (
            .O(N__36707),
            .I(N__36680));
    LocalMux I__7406 (
            .O(N__36702),
            .I(N__36677));
    LocalMux I__7405 (
            .O(N__36693),
            .I(N__36669));
    Span4Mux_v I__7404 (
            .O(N__36690),
            .I(N__36669));
    LocalMux I__7403 (
            .O(N__36687),
            .I(N__36666));
    InMux I__7402 (
            .O(N__36686),
            .I(N__36661));
    InMux I__7401 (
            .O(N__36685),
            .I(N__36661));
    LocalMux I__7400 (
            .O(N__36680),
            .I(N__36658));
    Span4Mux_v I__7399 (
            .O(N__36677),
            .I(N__36655));
    InMux I__7398 (
            .O(N__36676),
            .I(N__36648));
    InMux I__7397 (
            .O(N__36675),
            .I(N__36648));
    InMux I__7396 (
            .O(N__36674),
            .I(N__36648));
    Odrv4 I__7395 (
            .O(N__36669),
            .I(eis_end_N_725));
    Odrv12 I__7394 (
            .O(N__36666),
            .I(eis_end_N_725));
    LocalMux I__7393 (
            .O(N__36661),
            .I(eis_end_N_725));
    Odrv4 I__7392 (
            .O(N__36658),
            .I(eis_end_N_725));
    Odrv4 I__7391 (
            .O(N__36655),
            .I(eis_end_N_725));
    LocalMux I__7390 (
            .O(N__36648),
            .I(eis_end_N_725));
    CEMux I__7389 (
            .O(N__36635),
            .I(N__36631));
    CEMux I__7388 (
            .O(N__36634),
            .I(N__36628));
    LocalMux I__7387 (
            .O(N__36631),
            .I(N__36624));
    LocalMux I__7386 (
            .O(N__36628),
            .I(N__36621));
    CEMux I__7385 (
            .O(N__36627),
            .I(N__36618));
    Span4Mux_v I__7384 (
            .O(N__36624),
            .I(N__36614));
    Span4Mux_h I__7383 (
            .O(N__36621),
            .I(N__36609));
    LocalMux I__7382 (
            .O(N__36618),
            .I(N__36609));
    InMux I__7381 (
            .O(N__36617),
            .I(N__36606));
    Odrv4 I__7380 (
            .O(N__36614),
            .I(n11670));
    Odrv4 I__7379 (
            .O(N__36609),
            .I(n11670));
    LocalMux I__7378 (
            .O(N__36606),
            .I(n11670));
    SRMux I__7377 (
            .O(N__36599),
            .I(N__36595));
    SRMux I__7376 (
            .O(N__36598),
            .I(N__36592));
    LocalMux I__7375 (
            .O(N__36595),
            .I(n14687));
    LocalMux I__7374 (
            .O(N__36592),
            .I(n14687));
    InMux I__7373 (
            .O(N__36587),
            .I(N__36583));
    InMux I__7372 (
            .O(N__36586),
            .I(N__36579));
    LocalMux I__7371 (
            .O(N__36583),
            .I(N__36576));
    InMux I__7370 (
            .O(N__36582),
            .I(N__36573));
    LocalMux I__7369 (
            .O(N__36579),
            .I(N__36569));
    Span4Mux_v I__7368 (
            .O(N__36576),
            .I(N__36564));
    LocalMux I__7367 (
            .O(N__36573),
            .I(N__36564));
    InMux I__7366 (
            .O(N__36572),
            .I(N__36561));
    Span4Mux_v I__7365 (
            .O(N__36569),
            .I(N__36558));
    Span4Mux_h I__7364 (
            .O(N__36564),
            .I(N__36555));
    LocalMux I__7363 (
            .O(N__36561),
            .I(n10733));
    Odrv4 I__7362 (
            .O(N__36558),
            .I(n10733));
    Odrv4 I__7361 (
            .O(N__36555),
            .I(n10733));
    InMux I__7360 (
            .O(N__36548),
            .I(N__36544));
    InMux I__7359 (
            .O(N__36547),
            .I(N__36540));
    LocalMux I__7358 (
            .O(N__36544),
            .I(N__36537));
    InMux I__7357 (
            .O(N__36543),
            .I(N__36534));
    LocalMux I__7356 (
            .O(N__36540),
            .I(N__36531));
    Odrv12 I__7355 (
            .O(N__36537),
            .I(buf_dds0_5));
    LocalMux I__7354 (
            .O(N__36534),
            .I(buf_dds0_5));
    Odrv4 I__7353 (
            .O(N__36531),
            .I(buf_dds0_5));
    CascadeMux I__7352 (
            .O(N__36524),
            .I(n27_adj_1551_cascade_));
    InMux I__7351 (
            .O(N__36521),
            .I(N__36518));
    LocalMux I__7350 (
            .O(N__36518),
            .I(n25));
    CascadeMux I__7349 (
            .O(N__36515),
            .I(n19608_cascade_));
    InMux I__7348 (
            .O(N__36512),
            .I(N__36509));
    LocalMux I__7347 (
            .O(N__36509),
            .I(n10_adj_1594));
    InMux I__7346 (
            .O(N__36506),
            .I(N__36503));
    LocalMux I__7345 (
            .O(N__36503),
            .I(n26_adj_1543));
    InMux I__7344 (
            .O(N__36500),
            .I(N__36497));
    LocalMux I__7343 (
            .O(N__36497),
            .I(N__36493));
    InMux I__7342 (
            .O(N__36496),
            .I(N__36490));
    Span4Mux_h I__7341 (
            .O(N__36493),
            .I(N__36487));
    LocalMux I__7340 (
            .O(N__36490),
            .I(acadc_skipcnt_15));
    Odrv4 I__7339 (
            .O(N__36487),
            .I(acadc_skipcnt_15));
    InMux I__7338 (
            .O(N__36482),
            .I(N__36478));
    InMux I__7337 (
            .O(N__36481),
            .I(N__36475));
    LocalMux I__7336 (
            .O(N__36478),
            .I(N__36472));
    LocalMux I__7335 (
            .O(N__36475),
            .I(acadc_skipcnt_9));
    Odrv4 I__7334 (
            .O(N__36472),
            .I(acadc_skipcnt_9));
    InMux I__7333 (
            .O(N__36467),
            .I(N__36464));
    LocalMux I__7332 (
            .O(N__36464),
            .I(n21));
    CascadeMux I__7331 (
            .O(N__36461),
            .I(n24_adj_1537_cascade_));
    InMux I__7330 (
            .O(N__36458),
            .I(N__36455));
    LocalMux I__7329 (
            .O(N__36455),
            .I(n23_adj_1624));
    InMux I__7328 (
            .O(N__36452),
            .I(N__36449));
    LocalMux I__7327 (
            .O(N__36449),
            .I(n30));
    SRMux I__7326 (
            .O(N__36446),
            .I(N__36443));
    LocalMux I__7325 (
            .O(N__36443),
            .I(N__36440));
    Odrv4 I__7324 (
            .O(N__36440),
            .I(n20789));
    CascadeMux I__7323 (
            .O(N__36437),
            .I(N__36434));
    InMux I__7322 (
            .O(N__36434),
            .I(N__36428));
    InMux I__7321 (
            .O(N__36433),
            .I(N__36425));
    InMux I__7320 (
            .O(N__36432),
            .I(N__36422));
    CascadeMux I__7319 (
            .O(N__36431),
            .I(N__36411));
    LocalMux I__7318 (
            .O(N__36428),
            .I(N__36408));
    LocalMux I__7317 (
            .O(N__36425),
            .I(N__36405));
    LocalMux I__7316 (
            .O(N__36422),
            .I(N__36402));
    InMux I__7315 (
            .O(N__36421),
            .I(N__36399));
    InMux I__7314 (
            .O(N__36420),
            .I(N__36396));
    InMux I__7313 (
            .O(N__36419),
            .I(N__36391));
    InMux I__7312 (
            .O(N__36418),
            .I(N__36391));
    InMux I__7311 (
            .O(N__36417),
            .I(N__36382));
    InMux I__7310 (
            .O(N__36416),
            .I(N__36382));
    InMux I__7309 (
            .O(N__36415),
            .I(N__36382));
    InMux I__7308 (
            .O(N__36414),
            .I(N__36382));
    InMux I__7307 (
            .O(N__36411),
            .I(N__36379));
    Span4Mux_v I__7306 (
            .O(N__36408),
            .I(N__36370));
    Span4Mux_v I__7305 (
            .O(N__36405),
            .I(N__36370));
    Span4Mux_h I__7304 (
            .O(N__36402),
            .I(N__36370));
    LocalMux I__7303 (
            .O(N__36399),
            .I(N__36370));
    LocalMux I__7302 (
            .O(N__36396),
            .I(eis_state_0));
    LocalMux I__7301 (
            .O(N__36391),
            .I(eis_state_0));
    LocalMux I__7300 (
            .O(N__36382),
            .I(eis_state_0));
    LocalMux I__7299 (
            .O(N__36379),
            .I(eis_state_0));
    Odrv4 I__7298 (
            .O(N__36370),
            .I(eis_state_0));
    InMux I__7297 (
            .O(N__36359),
            .I(N__36356));
    LocalMux I__7296 (
            .O(N__36356),
            .I(N__36353));
    Span4Mux_v I__7295 (
            .O(N__36353),
            .I(N__36349));
    SRMux I__7294 (
            .O(N__36352),
            .I(N__36346));
    Span4Mux_v I__7293 (
            .O(N__36349),
            .I(N__36339));
    LocalMux I__7292 (
            .O(N__36346),
            .I(N__36339));
    InMux I__7291 (
            .O(N__36345),
            .I(N__36330));
    InMux I__7290 (
            .O(N__36344),
            .I(N__36330));
    Span4Mux_h I__7289 (
            .O(N__36339),
            .I(N__36327));
    SRMux I__7288 (
            .O(N__36338),
            .I(N__36324));
    InMux I__7287 (
            .O(N__36337),
            .I(N__36321));
    InMux I__7286 (
            .O(N__36336),
            .I(N__36316));
    InMux I__7285 (
            .O(N__36335),
            .I(N__36316));
    LocalMux I__7284 (
            .O(N__36330),
            .I(N__36313));
    Odrv4 I__7283 (
            .O(N__36327),
            .I(acadc_rst));
    LocalMux I__7282 (
            .O(N__36324),
            .I(acadc_rst));
    LocalMux I__7281 (
            .O(N__36321),
            .I(acadc_rst));
    LocalMux I__7280 (
            .O(N__36316),
            .I(acadc_rst));
    Odrv12 I__7279 (
            .O(N__36313),
            .I(acadc_rst));
    InMux I__7278 (
            .O(N__36302),
            .I(N__36299));
    LocalMux I__7277 (
            .O(N__36299),
            .I(N__36296));
    Sp12to4 I__7276 (
            .O(N__36296),
            .I(N__36292));
    InMux I__7275 (
            .O(N__36295),
            .I(N__36288));
    Span12Mux_v I__7274 (
            .O(N__36292),
            .I(N__36285));
    InMux I__7273 (
            .O(N__36291),
            .I(N__36282));
    LocalMux I__7272 (
            .O(N__36288),
            .I(buf_dds1_5));
    Odrv12 I__7271 (
            .O(N__36285),
            .I(buf_dds1_5));
    LocalMux I__7270 (
            .O(N__36282),
            .I(buf_dds1_5));
    InMux I__7269 (
            .O(N__36275),
            .I(N__36271));
    CascadeMux I__7268 (
            .O(N__36274),
            .I(N__36268));
    LocalMux I__7267 (
            .O(N__36271),
            .I(N__36265));
    InMux I__7266 (
            .O(N__36268),
            .I(N__36262));
    Span4Mux_v I__7265 (
            .O(N__36265),
            .I(N__36259));
    LocalMux I__7264 (
            .O(N__36262),
            .I(data_idxvec_14));
    Odrv4 I__7263 (
            .O(N__36259),
            .I(data_idxvec_14));
    InMux I__7262 (
            .O(N__36254),
            .I(N__36250));
    InMux I__7261 (
            .O(N__36253),
            .I(N__36247));
    LocalMux I__7260 (
            .O(N__36250),
            .I(N__36244));
    LocalMux I__7259 (
            .O(N__36247),
            .I(acadc_skipcnt_5));
    Odrv4 I__7258 (
            .O(N__36244),
            .I(acadc_skipcnt_5));
    InMux I__7257 (
            .O(N__36239),
            .I(N__36236));
    LocalMux I__7256 (
            .O(N__36236),
            .I(N__36232));
    InMux I__7255 (
            .O(N__36235),
            .I(N__36229));
    Span4Mux_h I__7254 (
            .O(N__36232),
            .I(N__36226));
    LocalMux I__7253 (
            .O(N__36229),
            .I(acadc_skipcnt_3));
    Odrv4 I__7252 (
            .O(N__36226),
            .I(acadc_skipcnt_3));
    InMux I__7251 (
            .O(N__36221),
            .I(N__36218));
    LocalMux I__7250 (
            .O(N__36218),
            .I(N__36214));
    InMux I__7249 (
            .O(N__36217),
            .I(N__36211));
    Span4Mux_h I__7248 (
            .O(N__36214),
            .I(N__36208));
    LocalMux I__7247 (
            .O(N__36211),
            .I(acadc_skipcnt_8));
    Odrv4 I__7246 (
            .O(N__36208),
            .I(acadc_skipcnt_8));
    CascadeMux I__7245 (
            .O(N__36203),
            .I(n20_adj_1617_cascade_));
    InMux I__7244 (
            .O(N__36200),
            .I(N__36197));
    LocalMux I__7243 (
            .O(N__36197),
            .I(n17_adj_1612));
    CascadeMux I__7242 (
            .O(N__36194),
            .I(n26_adj_1640_cascade_));
    InMux I__7241 (
            .O(N__36191),
            .I(N__36185));
    InMux I__7240 (
            .O(N__36190),
            .I(N__36185));
    LocalMux I__7239 (
            .O(N__36185),
            .I(n31));
    InMux I__7238 (
            .O(N__36182),
            .I(N__36177));
    InMux I__7237 (
            .O(N__36181),
            .I(N__36174));
    InMux I__7236 (
            .O(N__36180),
            .I(N__36171));
    LocalMux I__7235 (
            .O(N__36177),
            .I(N__36166));
    LocalMux I__7234 (
            .O(N__36174),
            .I(N__36166));
    LocalMux I__7233 (
            .O(N__36171),
            .I(N__36161));
    Span4Mux_v I__7232 (
            .O(N__36166),
            .I(N__36161));
    Odrv4 I__7231 (
            .O(N__36161),
            .I(data_index_2));
    CascadeMux I__7230 (
            .O(N__36158),
            .I(n11_cascade_));
    CascadeMux I__7229 (
            .O(N__36155),
            .I(n21099_cascade_));
    InMux I__7228 (
            .O(N__36152),
            .I(N__36149));
    LocalMux I__7227 (
            .O(N__36149),
            .I(n13));
    CEMux I__7226 (
            .O(N__36146),
            .I(N__36143));
    LocalMux I__7225 (
            .O(N__36143),
            .I(N__36139));
    CEMux I__7224 (
            .O(N__36142),
            .I(N__36136));
    Span4Mux_v I__7223 (
            .O(N__36139),
            .I(N__36131));
    LocalMux I__7222 (
            .O(N__36136),
            .I(N__36131));
    Odrv4 I__7221 (
            .O(N__36131),
            .I(n11760));
    InMux I__7220 (
            .O(N__36128),
            .I(N__36125));
    LocalMux I__7219 (
            .O(N__36125),
            .I(n17430));
    CascadeMux I__7218 (
            .O(N__36122),
            .I(N__36115));
    CascadeMux I__7217 (
            .O(N__36121),
            .I(N__36112));
    InMux I__7216 (
            .O(N__36120),
            .I(N__36106));
    InMux I__7215 (
            .O(N__36119),
            .I(N__36106));
    InMux I__7214 (
            .O(N__36118),
            .I(N__36103));
    InMux I__7213 (
            .O(N__36115),
            .I(N__36096));
    InMux I__7212 (
            .O(N__36112),
            .I(N__36096));
    InMux I__7211 (
            .O(N__36111),
            .I(N__36096));
    LocalMux I__7210 (
            .O(N__36106),
            .I(N__36093));
    LocalMux I__7209 (
            .O(N__36103),
            .I(acadc_dtrig_v));
    LocalMux I__7208 (
            .O(N__36096),
            .I(acadc_dtrig_v));
    Odrv4 I__7207 (
            .O(N__36093),
            .I(acadc_dtrig_v));
    InMux I__7206 (
            .O(N__36086),
            .I(N__36072));
    InMux I__7205 (
            .O(N__36085),
            .I(N__36072));
    InMux I__7204 (
            .O(N__36084),
            .I(N__36072));
    InMux I__7203 (
            .O(N__36083),
            .I(N__36072));
    InMux I__7202 (
            .O(N__36082),
            .I(N__36067));
    InMux I__7201 (
            .O(N__36081),
            .I(N__36067));
    LocalMux I__7200 (
            .O(N__36072),
            .I(acadc_dtrig_i));
    LocalMux I__7199 (
            .O(N__36067),
            .I(acadc_dtrig_i));
    CascadeMux I__7198 (
            .O(N__36062),
            .I(N__36059));
    InMux I__7197 (
            .O(N__36059),
            .I(N__36056));
    LocalMux I__7196 (
            .O(N__36056),
            .I(N__36053));
    Span4Mux_v I__7195 (
            .O(N__36053),
            .I(N__36050));
    Odrv4 I__7194 (
            .O(N__36050),
            .I(n4_adj_1569));
    InMux I__7193 (
            .O(N__36047),
            .I(N__36043));
    InMux I__7192 (
            .O(N__36046),
            .I(N__36040));
    LocalMux I__7191 (
            .O(N__36043),
            .I(N__36034));
    LocalMux I__7190 (
            .O(N__36040),
            .I(N__36034));
    InMux I__7189 (
            .O(N__36039),
            .I(N__36031));
    Span4Mux_h I__7188 (
            .O(N__36034),
            .I(N__36028));
    LocalMux I__7187 (
            .O(N__36031),
            .I(data_index_3));
    Odrv4 I__7186 (
            .O(N__36028),
            .I(data_index_3));
    InMux I__7185 (
            .O(N__36023),
            .I(N__36020));
    LocalMux I__7184 (
            .O(N__36020),
            .I(n8_adj_1563));
    CascadeMux I__7183 (
            .O(N__36017),
            .I(n8_adj_1563_cascade_));
    InMux I__7182 (
            .O(N__36014),
            .I(N__36008));
    InMux I__7181 (
            .O(N__36013),
            .I(N__36008));
    LocalMux I__7180 (
            .O(N__36008),
            .I(N__36005));
    Odrv4 I__7179 (
            .O(N__36005),
            .I(n7_adj_1562));
    CascadeMux I__7178 (
            .O(N__36002),
            .I(N__35999));
    CascadeBuf I__7177 (
            .O(N__35999),
            .I(N__35996));
    CascadeMux I__7176 (
            .O(N__35996),
            .I(N__35993));
    CascadeBuf I__7175 (
            .O(N__35993),
            .I(N__35990));
    CascadeMux I__7174 (
            .O(N__35990),
            .I(N__35987));
    CascadeBuf I__7173 (
            .O(N__35987),
            .I(N__35984));
    CascadeMux I__7172 (
            .O(N__35984),
            .I(N__35981));
    CascadeBuf I__7171 (
            .O(N__35981),
            .I(N__35978));
    CascadeMux I__7170 (
            .O(N__35978),
            .I(N__35975));
    CascadeBuf I__7169 (
            .O(N__35975),
            .I(N__35972));
    CascadeMux I__7168 (
            .O(N__35972),
            .I(N__35969));
    CascadeBuf I__7167 (
            .O(N__35969),
            .I(N__35966));
    CascadeMux I__7166 (
            .O(N__35966),
            .I(N__35963));
    CascadeBuf I__7165 (
            .O(N__35963),
            .I(N__35960));
    CascadeMux I__7164 (
            .O(N__35960),
            .I(N__35956));
    CascadeMux I__7163 (
            .O(N__35959),
            .I(N__35953));
    CascadeBuf I__7162 (
            .O(N__35956),
            .I(N__35950));
    CascadeBuf I__7161 (
            .O(N__35953),
            .I(N__35947));
    CascadeMux I__7160 (
            .O(N__35950),
            .I(N__35944));
    CascadeMux I__7159 (
            .O(N__35947),
            .I(N__35941));
    CascadeBuf I__7158 (
            .O(N__35944),
            .I(N__35938));
    InMux I__7157 (
            .O(N__35941),
            .I(N__35935));
    CascadeMux I__7156 (
            .O(N__35938),
            .I(N__35932));
    LocalMux I__7155 (
            .O(N__35935),
            .I(N__35929));
    InMux I__7154 (
            .O(N__35932),
            .I(N__35926));
    Span4Mux_v I__7153 (
            .O(N__35929),
            .I(N__35923));
    LocalMux I__7152 (
            .O(N__35926),
            .I(N__35920));
    Span4Mux_v I__7151 (
            .O(N__35923),
            .I(N__35917));
    Span4Mux_v I__7150 (
            .O(N__35920),
            .I(N__35914));
    Span4Mux_h I__7149 (
            .O(N__35917),
            .I(N__35911));
    Span4Mux_h I__7148 (
            .O(N__35914),
            .I(N__35908));
    Span4Mux_h I__7147 (
            .O(N__35911),
            .I(N__35905));
    Span4Mux_h I__7146 (
            .O(N__35908),
            .I(N__35902));
    Odrv4 I__7145 (
            .O(N__35905),
            .I(data_index_9_N_216_3));
    Odrv4 I__7144 (
            .O(N__35902),
            .I(data_index_9_N_216_3));
    CascadeMux I__7143 (
            .O(N__35897),
            .I(N__35894));
    InMux I__7142 (
            .O(N__35894),
            .I(N__35891));
    LocalMux I__7141 (
            .O(N__35891),
            .I(N__35888));
    Odrv4 I__7140 (
            .O(N__35888),
            .I(n16598));
    InMux I__7139 (
            .O(N__35885),
            .I(N__35882));
    LocalMux I__7138 (
            .O(N__35882),
            .I(N__35879));
    Odrv4 I__7137 (
            .O(N__35879),
            .I(n20957));
    InMux I__7136 (
            .O(N__35876),
            .I(N__35873));
    LocalMux I__7135 (
            .O(N__35873),
            .I(N__35870));
    Span4Mux_h I__7134 (
            .O(N__35870),
            .I(N__35864));
    InMux I__7133 (
            .O(N__35869),
            .I(N__35861));
    CascadeMux I__7132 (
            .O(N__35868),
            .I(N__35852));
    CascadeMux I__7131 (
            .O(N__35867),
            .I(N__35848));
    Span4Mux_h I__7130 (
            .O(N__35864),
            .I(N__35844));
    LocalMux I__7129 (
            .O(N__35861),
            .I(N__35841));
    InMux I__7128 (
            .O(N__35860),
            .I(N__35836));
    InMux I__7127 (
            .O(N__35859),
            .I(N__35836));
    InMux I__7126 (
            .O(N__35858),
            .I(N__35831));
    InMux I__7125 (
            .O(N__35857),
            .I(N__35831));
    InMux I__7124 (
            .O(N__35856),
            .I(N__35828));
    InMux I__7123 (
            .O(N__35855),
            .I(N__35817));
    InMux I__7122 (
            .O(N__35852),
            .I(N__35817));
    InMux I__7121 (
            .O(N__35851),
            .I(N__35817));
    InMux I__7120 (
            .O(N__35848),
            .I(N__35817));
    InMux I__7119 (
            .O(N__35847),
            .I(N__35817));
    Odrv4 I__7118 (
            .O(N__35844),
            .I(DTRIG_N_919_adj_1451));
    Odrv4 I__7117 (
            .O(N__35841),
            .I(DTRIG_N_919_adj_1451));
    LocalMux I__7116 (
            .O(N__35836),
            .I(DTRIG_N_919_adj_1451));
    LocalMux I__7115 (
            .O(N__35831),
            .I(DTRIG_N_919_adj_1451));
    LocalMux I__7114 (
            .O(N__35828),
            .I(DTRIG_N_919_adj_1451));
    LocalMux I__7113 (
            .O(N__35817),
            .I(DTRIG_N_919_adj_1451));
    InMux I__7112 (
            .O(N__35804),
            .I(N__35800));
    InMux I__7111 (
            .O(N__35803),
            .I(N__35796));
    LocalMux I__7110 (
            .O(N__35800),
            .I(N__35793));
    InMux I__7109 (
            .O(N__35799),
            .I(N__35781));
    LocalMux I__7108 (
            .O(N__35796),
            .I(N__35776));
    Span12Mux_h I__7107 (
            .O(N__35793),
            .I(N__35776));
    InMux I__7106 (
            .O(N__35792),
            .I(N__35769));
    InMux I__7105 (
            .O(N__35791),
            .I(N__35769));
    InMux I__7104 (
            .O(N__35790),
            .I(N__35769));
    InMux I__7103 (
            .O(N__35789),
            .I(N__35766));
    InMux I__7102 (
            .O(N__35788),
            .I(N__35761));
    InMux I__7101 (
            .O(N__35787),
            .I(N__35761));
    InMux I__7100 (
            .O(N__35786),
            .I(N__35754));
    InMux I__7099 (
            .O(N__35785),
            .I(N__35754));
    InMux I__7098 (
            .O(N__35784),
            .I(N__35754));
    LocalMux I__7097 (
            .O(N__35781),
            .I(adc_state_1_adj_1417));
    Odrv12 I__7096 (
            .O(N__35776),
            .I(adc_state_1_adj_1417));
    LocalMux I__7095 (
            .O(N__35769),
            .I(adc_state_1_adj_1417));
    LocalMux I__7094 (
            .O(N__35766),
            .I(adc_state_1_adj_1417));
    LocalMux I__7093 (
            .O(N__35761),
            .I(adc_state_1_adj_1417));
    LocalMux I__7092 (
            .O(N__35754),
            .I(adc_state_1_adj_1417));
    InMux I__7091 (
            .O(N__35741),
            .I(N__35738));
    LocalMux I__7090 (
            .O(N__35738),
            .I(N__35735));
    Span4Mux_v I__7089 (
            .O(N__35735),
            .I(N__35732));
    Sp12to4 I__7088 (
            .O(N__35732),
            .I(N__35729));
    Span12Mux_h I__7087 (
            .O(N__35729),
            .I(N__35726));
    Span12Mux_v I__7086 (
            .O(N__35726),
            .I(N__35723));
    Odrv12 I__7085 (
            .O(N__35723),
            .I(ICE_GPMO_0));
    InMux I__7084 (
            .O(N__35720),
            .I(N__35717));
    LocalMux I__7083 (
            .O(N__35717),
            .I(N__35713));
    InMux I__7082 (
            .O(N__35716),
            .I(N__35710));
    Span4Mux_v I__7081 (
            .O(N__35713),
            .I(N__35707));
    LocalMux I__7080 (
            .O(N__35710),
            .I(N__35704));
    Span4Mux_h I__7079 (
            .O(N__35707),
            .I(N__35699));
    Span4Mux_v I__7078 (
            .O(N__35704),
            .I(N__35699));
    Span4Mux_v I__7077 (
            .O(N__35699),
            .I(N__35694));
    InMux I__7076 (
            .O(N__35698),
            .I(N__35691));
    InMux I__7075 (
            .O(N__35697),
            .I(N__35688));
    Odrv4 I__7074 (
            .O(N__35694),
            .I(auxmode));
    LocalMux I__7073 (
            .O(N__35691),
            .I(auxmode));
    LocalMux I__7072 (
            .O(N__35688),
            .I(auxmode));
    CascadeMux I__7071 (
            .O(N__35681),
            .I(acadc_rst_cascade_));
    InMux I__7070 (
            .O(N__35678),
            .I(N__35675));
    LocalMux I__7069 (
            .O(N__35675),
            .I(N__35670));
    InMux I__7068 (
            .O(N__35674),
            .I(N__35665));
    InMux I__7067 (
            .O(N__35673),
            .I(N__35665));
    Odrv4 I__7066 (
            .O(N__35670),
            .I(tacadc_rst));
    LocalMux I__7065 (
            .O(N__35665),
            .I(tacadc_rst));
    InMux I__7064 (
            .O(N__35660),
            .I(N__35657));
    LocalMux I__7063 (
            .O(N__35657),
            .I(N__35654));
    Span4Mux_h I__7062 (
            .O(N__35654),
            .I(N__35650));
    InMux I__7061 (
            .O(N__35653),
            .I(N__35647));
    Odrv4 I__7060 (
            .O(N__35650),
            .I(buf_readRTD_7));
    LocalMux I__7059 (
            .O(N__35647),
            .I(buf_readRTD_7));
    InMux I__7058 (
            .O(N__35642),
            .I(N__35639));
    LocalMux I__7057 (
            .O(N__35639),
            .I(N__35636));
    Span4Mux_v I__7056 (
            .O(N__35636),
            .I(N__35633));
    Odrv4 I__7055 (
            .O(N__35633),
            .I(n19_adj_1502));
    CascadeMux I__7054 (
            .O(N__35630),
            .I(n24_adj_1622_cascade_));
    InMux I__7053 (
            .O(N__35627),
            .I(N__35624));
    LocalMux I__7052 (
            .O(N__35624),
            .I(N__35621));
    Span4Mux_v I__7051 (
            .O(N__35621),
            .I(N__35618));
    Span4Mux_v I__7050 (
            .O(N__35618),
            .I(N__35615));
    Span4Mux_h I__7049 (
            .O(N__35615),
            .I(N__35611));
    InMux I__7048 (
            .O(N__35614),
            .I(N__35608));
    Odrv4 I__7047 (
            .O(N__35611),
            .I(buf_adcdata_vdc_12));
    LocalMux I__7046 (
            .O(N__35608),
            .I(buf_adcdata_vdc_12));
    InMux I__7045 (
            .O(N__35603),
            .I(N__35600));
    LocalMux I__7044 (
            .O(N__35600),
            .I(N__35597));
    Span4Mux_v I__7043 (
            .O(N__35597),
            .I(N__35594));
    Span4Mux_h I__7042 (
            .O(N__35594),
            .I(N__35590));
    InMux I__7041 (
            .O(N__35593),
            .I(N__35586));
    Span4Mux_h I__7040 (
            .O(N__35590),
            .I(N__35583));
    InMux I__7039 (
            .O(N__35589),
            .I(N__35580));
    LocalMux I__7038 (
            .O(N__35586),
            .I(buf_adcdata_vac_12));
    Odrv4 I__7037 (
            .O(N__35583),
            .I(buf_adcdata_vac_12));
    LocalMux I__7036 (
            .O(N__35580),
            .I(buf_adcdata_vac_12));
    CascadeMux I__7035 (
            .O(N__35573),
            .I(n35_cascade_));
    SRMux I__7034 (
            .O(N__35570),
            .I(N__35563));
    SRMux I__7033 (
            .O(N__35569),
            .I(N__35559));
    SRMux I__7032 (
            .O(N__35568),
            .I(N__35555));
    SRMux I__7031 (
            .O(N__35567),
            .I(N__35551));
    SRMux I__7030 (
            .O(N__35566),
            .I(N__35547));
    LocalMux I__7029 (
            .O(N__35563),
            .I(N__35543));
    SRMux I__7028 (
            .O(N__35562),
            .I(N__35540));
    LocalMux I__7027 (
            .O(N__35559),
            .I(N__35536));
    SRMux I__7026 (
            .O(N__35558),
            .I(N__35533));
    LocalMux I__7025 (
            .O(N__35555),
            .I(N__35530));
    SRMux I__7024 (
            .O(N__35554),
            .I(N__35527));
    LocalMux I__7023 (
            .O(N__35551),
            .I(N__35524));
    SRMux I__7022 (
            .O(N__35550),
            .I(N__35521));
    LocalMux I__7021 (
            .O(N__35547),
            .I(N__35518));
    SRMux I__7020 (
            .O(N__35546),
            .I(N__35515));
    Span4Mux_v I__7019 (
            .O(N__35543),
            .I(N__35510));
    LocalMux I__7018 (
            .O(N__35540),
            .I(N__35510));
    SRMux I__7017 (
            .O(N__35539),
            .I(N__35507));
    Span4Mux_v I__7016 (
            .O(N__35536),
            .I(N__35501));
    LocalMux I__7015 (
            .O(N__35533),
            .I(N__35501));
    Span4Mux_h I__7014 (
            .O(N__35530),
            .I(N__35498));
    LocalMux I__7013 (
            .O(N__35527),
            .I(N__35495));
    Span4Mux_h I__7012 (
            .O(N__35524),
            .I(N__35492));
    LocalMux I__7011 (
            .O(N__35521),
            .I(N__35489));
    Span4Mux_v I__7010 (
            .O(N__35518),
            .I(N__35484));
    LocalMux I__7009 (
            .O(N__35515),
            .I(N__35484));
    Span4Mux_v I__7008 (
            .O(N__35510),
            .I(N__35479));
    LocalMux I__7007 (
            .O(N__35507),
            .I(N__35479));
    SRMux I__7006 (
            .O(N__35506),
            .I(N__35476));
    Span4Mux_v I__7005 (
            .O(N__35501),
            .I(N__35473));
    Span4Mux_v I__7004 (
            .O(N__35498),
            .I(N__35468));
    Span4Mux_h I__7003 (
            .O(N__35495),
            .I(N__35468));
    Span4Mux_v I__7002 (
            .O(N__35492),
            .I(N__35463));
    Span4Mux_h I__7001 (
            .O(N__35489),
            .I(N__35463));
    Span4Mux_v I__7000 (
            .O(N__35484),
            .I(N__35458));
    Span4Mux_v I__6999 (
            .O(N__35479),
            .I(N__35458));
    LocalMux I__6998 (
            .O(N__35476),
            .I(N__35455));
    Span4Mux_h I__6997 (
            .O(N__35473),
            .I(N__35452));
    Span4Mux_v I__6996 (
            .O(N__35468),
            .I(N__35443));
    Span4Mux_v I__6995 (
            .O(N__35463),
            .I(N__35443));
    Span4Mux_h I__6994 (
            .O(N__35458),
            .I(N__35443));
    Span4Mux_h I__6993 (
            .O(N__35455),
            .I(N__35443));
    Span4Mux_h I__6992 (
            .O(N__35452),
            .I(N__35440));
    Span4Mux_h I__6991 (
            .O(N__35443),
            .I(N__35437));
    Odrv4 I__6990 (
            .O(N__35440),
            .I(iac_raw_buf_N_735));
    Odrv4 I__6989 (
            .O(N__35437),
            .I(iac_raw_buf_N_735));
    InMux I__6988 (
            .O(N__35432),
            .I(N__35429));
    LocalMux I__6987 (
            .O(N__35429),
            .I(N__35426));
    Odrv4 I__6986 (
            .O(N__35426),
            .I(n17_adj_1645));
    CascadeMux I__6985 (
            .O(N__35423),
            .I(N__35413));
    CascadeMux I__6984 (
            .O(N__35422),
            .I(N__35397));
    InMux I__6983 (
            .O(N__35421),
            .I(N__35387));
    InMux I__6982 (
            .O(N__35420),
            .I(N__35382));
    InMux I__6981 (
            .O(N__35419),
            .I(N__35382));
    InMux I__6980 (
            .O(N__35418),
            .I(N__35377));
    InMux I__6979 (
            .O(N__35417),
            .I(N__35377));
    InMux I__6978 (
            .O(N__35416),
            .I(N__35373));
    InMux I__6977 (
            .O(N__35413),
            .I(N__35358));
    InMux I__6976 (
            .O(N__35412),
            .I(N__35353));
    InMux I__6975 (
            .O(N__35411),
            .I(N__35353));
    InMux I__6974 (
            .O(N__35410),
            .I(N__35348));
    InMux I__6973 (
            .O(N__35409),
            .I(N__35348));
    InMux I__6972 (
            .O(N__35408),
            .I(N__35332));
    InMux I__6971 (
            .O(N__35407),
            .I(N__35332));
    InMux I__6970 (
            .O(N__35406),
            .I(N__35332));
    InMux I__6969 (
            .O(N__35405),
            .I(N__35332));
    InMux I__6968 (
            .O(N__35404),
            .I(N__35321));
    InMux I__6967 (
            .O(N__35403),
            .I(N__35321));
    InMux I__6966 (
            .O(N__35402),
            .I(N__35321));
    InMux I__6965 (
            .O(N__35401),
            .I(N__35321));
    InMux I__6964 (
            .O(N__35400),
            .I(N__35321));
    InMux I__6963 (
            .O(N__35397),
            .I(N__35316));
    InMux I__6962 (
            .O(N__35396),
            .I(N__35307));
    InMux I__6961 (
            .O(N__35395),
            .I(N__35307));
    InMux I__6960 (
            .O(N__35394),
            .I(N__35307));
    InMux I__6959 (
            .O(N__35393),
            .I(N__35307));
    InMux I__6958 (
            .O(N__35392),
            .I(N__35298));
    InMux I__6957 (
            .O(N__35391),
            .I(N__35298));
    InMux I__6956 (
            .O(N__35390),
            .I(N__35298));
    LocalMux I__6955 (
            .O(N__35387),
            .I(N__35291));
    LocalMux I__6954 (
            .O(N__35382),
            .I(N__35291));
    LocalMux I__6953 (
            .O(N__35377),
            .I(N__35291));
    InMux I__6952 (
            .O(N__35376),
            .I(N__35288));
    LocalMux I__6951 (
            .O(N__35373),
            .I(N__35285));
    InMux I__6950 (
            .O(N__35372),
            .I(N__35270));
    InMux I__6949 (
            .O(N__35371),
            .I(N__35270));
    InMux I__6948 (
            .O(N__35370),
            .I(N__35270));
    InMux I__6947 (
            .O(N__35369),
            .I(N__35270));
    InMux I__6946 (
            .O(N__35368),
            .I(N__35270));
    InMux I__6945 (
            .O(N__35367),
            .I(N__35270));
    InMux I__6944 (
            .O(N__35366),
            .I(N__35270));
    InMux I__6943 (
            .O(N__35365),
            .I(N__35259));
    InMux I__6942 (
            .O(N__35364),
            .I(N__35259));
    InMux I__6941 (
            .O(N__35363),
            .I(N__35259));
    InMux I__6940 (
            .O(N__35362),
            .I(N__35259));
    InMux I__6939 (
            .O(N__35361),
            .I(N__35259));
    LocalMux I__6938 (
            .O(N__35358),
            .I(N__35256));
    LocalMux I__6937 (
            .O(N__35353),
            .I(N__35253));
    LocalMux I__6936 (
            .O(N__35348),
            .I(N__35250));
    InMux I__6935 (
            .O(N__35347),
            .I(N__35243));
    InMux I__6934 (
            .O(N__35346),
            .I(N__35243));
    InMux I__6933 (
            .O(N__35345),
            .I(N__35243));
    InMux I__6932 (
            .O(N__35344),
            .I(N__35234));
    InMux I__6931 (
            .O(N__35343),
            .I(N__35234));
    InMux I__6930 (
            .O(N__35342),
            .I(N__35234));
    InMux I__6929 (
            .O(N__35341),
            .I(N__35234));
    LocalMux I__6928 (
            .O(N__35332),
            .I(N__35229));
    LocalMux I__6927 (
            .O(N__35321),
            .I(N__35229));
    InMux I__6926 (
            .O(N__35320),
            .I(N__35224));
    InMux I__6925 (
            .O(N__35319),
            .I(N__35224));
    LocalMux I__6924 (
            .O(N__35316),
            .I(N__35219));
    LocalMux I__6923 (
            .O(N__35307),
            .I(N__35219));
    InMux I__6922 (
            .O(N__35306),
            .I(N__35211));
    InMux I__6921 (
            .O(N__35305),
            .I(N__35208));
    LocalMux I__6920 (
            .O(N__35298),
            .I(N__35205));
    Span4Mux_v I__6919 (
            .O(N__35291),
            .I(N__35202));
    LocalMux I__6918 (
            .O(N__35288),
            .I(N__35197));
    Span4Mux_v I__6917 (
            .O(N__35285),
            .I(N__35197));
    LocalMux I__6916 (
            .O(N__35270),
            .I(N__35192));
    LocalMux I__6915 (
            .O(N__35259),
            .I(N__35192));
    Span4Mux_v I__6914 (
            .O(N__35256),
            .I(N__35185));
    Span4Mux_v I__6913 (
            .O(N__35253),
            .I(N__35185));
    Span4Mux_v I__6912 (
            .O(N__35250),
            .I(N__35185));
    LocalMux I__6911 (
            .O(N__35243),
            .I(N__35178));
    LocalMux I__6910 (
            .O(N__35234),
            .I(N__35178));
    Span4Mux_h I__6909 (
            .O(N__35229),
            .I(N__35178));
    LocalMux I__6908 (
            .O(N__35224),
            .I(N__35175));
    Span4Mux_v I__6907 (
            .O(N__35219),
            .I(N__35172));
    InMux I__6906 (
            .O(N__35218),
            .I(N__35158));
    InMux I__6905 (
            .O(N__35217),
            .I(N__35158));
    InMux I__6904 (
            .O(N__35216),
            .I(N__35158));
    InMux I__6903 (
            .O(N__35215),
            .I(N__35153));
    InMux I__6902 (
            .O(N__35214),
            .I(N__35153));
    LocalMux I__6901 (
            .O(N__35211),
            .I(N__35150));
    LocalMux I__6900 (
            .O(N__35208),
            .I(N__35147));
    Span4Mux_h I__6899 (
            .O(N__35205),
            .I(N__35140));
    Span4Mux_v I__6898 (
            .O(N__35202),
            .I(N__35140));
    Span4Mux_h I__6897 (
            .O(N__35197),
            .I(N__35140));
    Span4Mux_v I__6896 (
            .O(N__35192),
            .I(N__35134));
    Span4Mux_h I__6895 (
            .O(N__35185),
            .I(N__35134));
    Span4Mux_h I__6894 (
            .O(N__35178),
            .I(N__35131));
    Span4Mux_h I__6893 (
            .O(N__35175),
            .I(N__35125));
    Span4Mux_h I__6892 (
            .O(N__35172),
            .I(N__35122));
    InMux I__6891 (
            .O(N__35171),
            .I(N__35115));
    InMux I__6890 (
            .O(N__35170),
            .I(N__35115));
    InMux I__6889 (
            .O(N__35169),
            .I(N__35115));
    InMux I__6888 (
            .O(N__35168),
            .I(N__35112));
    InMux I__6887 (
            .O(N__35167),
            .I(N__35109));
    InMux I__6886 (
            .O(N__35166),
            .I(N__35106));
    InMux I__6885 (
            .O(N__35165),
            .I(N__35103));
    LocalMux I__6884 (
            .O(N__35158),
            .I(N__35096));
    LocalMux I__6883 (
            .O(N__35153),
            .I(N__35096));
    Span4Mux_h I__6882 (
            .O(N__35150),
            .I(N__35096));
    Span12Mux_v I__6881 (
            .O(N__35147),
            .I(N__35091));
    Sp12to4 I__6880 (
            .O(N__35140),
            .I(N__35091));
    InMux I__6879 (
            .O(N__35139),
            .I(N__35088));
    Span4Mux_h I__6878 (
            .O(N__35134),
            .I(N__35083));
    Span4Mux_h I__6877 (
            .O(N__35131),
            .I(N__35083));
    InMux I__6876 (
            .O(N__35130),
            .I(N__35076));
    InMux I__6875 (
            .O(N__35129),
            .I(N__35076));
    InMux I__6874 (
            .O(N__35128),
            .I(N__35076));
    Span4Mux_v I__6873 (
            .O(N__35125),
            .I(N__35069));
    Span4Mux_h I__6872 (
            .O(N__35122),
            .I(N__35069));
    LocalMux I__6871 (
            .O(N__35115),
            .I(N__35069));
    LocalMux I__6870 (
            .O(N__35112),
            .I(adc_state_0));
    LocalMux I__6869 (
            .O(N__35109),
            .I(adc_state_0));
    LocalMux I__6868 (
            .O(N__35106),
            .I(adc_state_0));
    LocalMux I__6867 (
            .O(N__35103),
            .I(adc_state_0));
    Odrv4 I__6866 (
            .O(N__35096),
            .I(adc_state_0));
    Odrv12 I__6865 (
            .O(N__35091),
            .I(adc_state_0));
    LocalMux I__6864 (
            .O(N__35088),
            .I(adc_state_0));
    Odrv4 I__6863 (
            .O(N__35083),
            .I(adc_state_0));
    LocalMux I__6862 (
            .O(N__35076),
            .I(adc_state_0));
    Odrv4 I__6861 (
            .O(N__35069),
            .I(adc_state_0));
    InMux I__6860 (
            .O(N__35048),
            .I(N__35045));
    LocalMux I__6859 (
            .O(N__35045),
            .I(N__35041));
    InMux I__6858 (
            .O(N__35044),
            .I(N__35038));
    Span4Mux_v I__6857 (
            .O(N__35041),
            .I(N__35035));
    LocalMux I__6856 (
            .O(N__35038),
            .I(N__35032));
    Span4Mux_h I__6855 (
            .O(N__35035),
            .I(N__35026));
    Span4Mux_h I__6854 (
            .O(N__35032),
            .I(N__35021));
    InMux I__6853 (
            .O(N__35031),
            .I(N__35014));
    InMux I__6852 (
            .O(N__35030),
            .I(N__35009));
    InMux I__6851 (
            .O(N__35029),
            .I(N__35009));
    Span4Mux_h I__6850 (
            .O(N__35026),
            .I(N__35005));
    InMux I__6849 (
            .O(N__35025),
            .I(N__35000));
    InMux I__6848 (
            .O(N__35024),
            .I(N__35000));
    Span4Mux_h I__6847 (
            .O(N__35021),
            .I(N__34997));
    InMux I__6846 (
            .O(N__35020),
            .I(N__34988));
    InMux I__6845 (
            .O(N__35019),
            .I(N__34988));
    InMux I__6844 (
            .O(N__35018),
            .I(N__34988));
    InMux I__6843 (
            .O(N__35017),
            .I(N__34988));
    LocalMux I__6842 (
            .O(N__35014),
            .I(N__34983));
    LocalMux I__6841 (
            .O(N__35009),
            .I(N__34983));
    InMux I__6840 (
            .O(N__35008),
            .I(N__34980));
    Odrv4 I__6839 (
            .O(N__35005),
            .I(adc_state_1));
    LocalMux I__6838 (
            .O(N__35000),
            .I(adc_state_1));
    Odrv4 I__6837 (
            .O(N__34997),
            .I(adc_state_1));
    LocalMux I__6836 (
            .O(N__34988),
            .I(adc_state_1));
    Odrv12 I__6835 (
            .O(N__34983),
            .I(adc_state_1));
    LocalMux I__6834 (
            .O(N__34980),
            .I(adc_state_1));
    CascadeMux I__6833 (
            .O(N__34967),
            .I(N__34964));
    InMux I__6832 (
            .O(N__34964),
            .I(N__34961));
    LocalMux I__6831 (
            .O(N__34961),
            .I(N__34956));
    InMux I__6830 (
            .O(N__34960),
            .I(N__34953));
    CascadeMux I__6829 (
            .O(N__34959),
            .I(N__34950));
    Span4Mux_v I__6828 (
            .O(N__34956),
            .I(N__34946));
    LocalMux I__6827 (
            .O(N__34953),
            .I(N__34942));
    InMux I__6826 (
            .O(N__34950),
            .I(N__34933));
    InMux I__6825 (
            .O(N__34949),
            .I(N__34933));
    Span4Mux_h I__6824 (
            .O(N__34946),
            .I(N__34930));
    CascadeMux I__6823 (
            .O(N__34945),
            .I(N__34927));
    Span4Mux_v I__6822 (
            .O(N__34942),
            .I(N__34921));
    InMux I__6821 (
            .O(N__34941),
            .I(N__34918));
    InMux I__6820 (
            .O(N__34940),
            .I(N__34913));
    InMux I__6819 (
            .O(N__34939),
            .I(N__34913));
    InMux I__6818 (
            .O(N__34938),
            .I(N__34910));
    LocalMux I__6817 (
            .O(N__34933),
            .I(N__34905));
    Span4Mux_h I__6816 (
            .O(N__34930),
            .I(N__34905));
    InMux I__6815 (
            .O(N__34927),
            .I(N__34896));
    InMux I__6814 (
            .O(N__34926),
            .I(N__34896));
    InMux I__6813 (
            .O(N__34925),
            .I(N__34896));
    InMux I__6812 (
            .O(N__34924),
            .I(N__34896));
    Span4Mux_h I__6811 (
            .O(N__34921),
            .I(N__34893));
    LocalMux I__6810 (
            .O(N__34918),
            .I(N__34888));
    LocalMux I__6809 (
            .O(N__34913),
            .I(N__34888));
    LocalMux I__6808 (
            .O(N__34910),
            .I(DTRIG_N_919));
    Odrv4 I__6807 (
            .O(N__34905),
            .I(DTRIG_N_919));
    LocalMux I__6806 (
            .O(N__34896),
            .I(DTRIG_N_919));
    Odrv4 I__6805 (
            .O(N__34893),
            .I(DTRIG_N_919));
    Odrv12 I__6804 (
            .O(N__34888),
            .I(DTRIG_N_919));
    CascadeMux I__6803 (
            .O(N__34877),
            .I(N__34874));
    InMux I__6802 (
            .O(N__34874),
            .I(N__34871));
    LocalMux I__6801 (
            .O(N__34871),
            .I(N__34868));
    Odrv12 I__6800 (
            .O(N__34868),
            .I(n8));
    InMux I__6799 (
            .O(N__34865),
            .I(N__34861));
    CascadeMux I__6798 (
            .O(N__34864),
            .I(N__34858));
    LocalMux I__6797 (
            .O(N__34861),
            .I(N__34855));
    InMux I__6796 (
            .O(N__34858),
            .I(N__34852));
    Span4Mux_h I__6795 (
            .O(N__34855),
            .I(N__34849));
    LocalMux I__6794 (
            .O(N__34852),
            .I(N__34846));
    Odrv4 I__6793 (
            .O(N__34849),
            .I(n11354));
    Odrv4 I__6792 (
            .O(N__34846),
            .I(n11354));
    CascadeMux I__6791 (
            .O(N__34841),
            .I(n10534_cascade_));
    CascadeMux I__6790 (
            .O(N__34838),
            .I(N__34835));
    InMux I__6789 (
            .O(N__34835),
            .I(N__34831));
    CascadeMux I__6788 (
            .O(N__34834),
            .I(N__34826));
    LocalMux I__6787 (
            .O(N__34831),
            .I(N__34823));
    InMux I__6786 (
            .O(N__34830),
            .I(N__34820));
    InMux I__6785 (
            .O(N__34829),
            .I(N__34815));
    InMux I__6784 (
            .O(N__34826),
            .I(N__34815));
    Span4Mux_h I__6783 (
            .O(N__34823),
            .I(N__34812));
    LocalMux I__6782 (
            .O(N__34820),
            .I(N__34809));
    LocalMux I__6781 (
            .O(N__34815),
            .I(N__34806));
    Span4Mux_h I__6780 (
            .O(N__34812),
            .I(N__34803));
    Odrv4 I__6779 (
            .O(N__34809),
            .I(n20670));
    Odrv12 I__6778 (
            .O(N__34806),
            .I(n20670));
    Odrv4 I__6777 (
            .O(N__34803),
            .I(n20670));
    InMux I__6776 (
            .O(N__34796),
            .I(N__34792));
    InMux I__6775 (
            .O(N__34795),
            .I(N__34789));
    LocalMux I__6774 (
            .O(N__34792),
            .I(N__34786));
    LocalMux I__6773 (
            .O(N__34789),
            .I(N__34783));
    Span12Mux_h I__6772 (
            .O(N__34786),
            .I(N__34780));
    Span12Mux_v I__6771 (
            .O(N__34783),
            .I(N__34777));
    Odrv12 I__6770 (
            .O(N__34780),
            .I(n20672));
    Odrv12 I__6769 (
            .O(N__34777),
            .I(n20672));
    CascadeMux I__6768 (
            .O(N__34772),
            .I(N__34769));
    InMux I__6767 (
            .O(N__34769),
            .I(N__34766));
    LocalMux I__6766 (
            .O(N__34766),
            .I(N__34762));
    CascadeMux I__6765 (
            .O(N__34765),
            .I(N__34758));
    Span4Mux_h I__6764 (
            .O(N__34762),
            .I(N__34755));
    InMux I__6763 (
            .O(N__34761),
            .I(N__34750));
    InMux I__6762 (
            .O(N__34758),
            .I(N__34750));
    Odrv4 I__6761 (
            .O(N__34755),
            .I(cmd_rdadctmp_9));
    LocalMux I__6760 (
            .O(N__34750),
            .I(cmd_rdadctmp_9));
    InMux I__6759 (
            .O(N__34745),
            .I(N__34742));
    LocalMux I__6758 (
            .O(N__34742),
            .I(N__34738));
    InMux I__6757 (
            .O(N__34741),
            .I(N__34735));
    Span4Mux_h I__6756 (
            .O(N__34738),
            .I(N__34731));
    LocalMux I__6755 (
            .O(N__34735),
            .I(N__34728));
    InMux I__6754 (
            .O(N__34734),
            .I(N__34725));
    Span4Mux_h I__6753 (
            .O(N__34731),
            .I(N__34720));
    Span4Mux_h I__6752 (
            .O(N__34728),
            .I(N__34720));
    LocalMux I__6751 (
            .O(N__34725),
            .I(buf_adcdata_vac_1));
    Odrv4 I__6750 (
            .O(N__34720),
            .I(buf_adcdata_vac_1));
    InMux I__6749 (
            .O(N__34715),
            .I(N__34712));
    LocalMux I__6748 (
            .O(N__34712),
            .I(N__34709));
    Odrv4 I__6747 (
            .O(N__34709),
            .I(n20840));
    CascadeMux I__6746 (
            .O(N__34706),
            .I(N__34703));
    InMux I__6745 (
            .O(N__34703),
            .I(N__34698));
    InMux I__6744 (
            .O(N__34702),
            .I(N__34693));
    InMux I__6743 (
            .O(N__34701),
            .I(N__34693));
    LocalMux I__6742 (
            .O(N__34698),
            .I(cmd_rdadctmp_21));
    LocalMux I__6741 (
            .O(N__34693),
            .I(cmd_rdadctmp_21));
    CascadeMux I__6740 (
            .O(N__34688),
            .I(N__34683));
    CascadeMux I__6739 (
            .O(N__34687),
            .I(N__34680));
    CascadeMux I__6738 (
            .O(N__34686),
            .I(N__34677));
    InMux I__6737 (
            .O(N__34683),
            .I(N__34674));
    InMux I__6736 (
            .O(N__34680),
            .I(N__34671));
    InMux I__6735 (
            .O(N__34677),
            .I(N__34668));
    LocalMux I__6734 (
            .O(N__34674),
            .I(cmd_rdadctmp_20));
    LocalMux I__6733 (
            .O(N__34671),
            .I(cmd_rdadctmp_20));
    LocalMux I__6732 (
            .O(N__34668),
            .I(cmd_rdadctmp_20));
    InMux I__6731 (
            .O(N__34661),
            .I(N__34641));
    InMux I__6730 (
            .O(N__34660),
            .I(N__34641));
    InMux I__6729 (
            .O(N__34659),
            .I(N__34641));
    InMux I__6728 (
            .O(N__34658),
            .I(N__34638));
    InMux I__6727 (
            .O(N__34657),
            .I(N__34631));
    InMux I__6726 (
            .O(N__34656),
            .I(N__34631));
    InMux I__6725 (
            .O(N__34655),
            .I(N__34631));
    InMux I__6724 (
            .O(N__34654),
            .I(N__34628));
    InMux I__6723 (
            .O(N__34653),
            .I(N__34625));
    InMux I__6722 (
            .O(N__34652),
            .I(N__34618));
    InMux I__6721 (
            .O(N__34651),
            .I(N__34609));
    InMux I__6720 (
            .O(N__34650),
            .I(N__34609));
    InMux I__6719 (
            .O(N__34649),
            .I(N__34609));
    InMux I__6718 (
            .O(N__34648),
            .I(N__34609));
    LocalMux I__6717 (
            .O(N__34641),
            .I(N__34606));
    LocalMux I__6716 (
            .O(N__34638),
            .I(N__34599));
    LocalMux I__6715 (
            .O(N__34631),
            .I(N__34599));
    LocalMux I__6714 (
            .O(N__34628),
            .I(N__34599));
    LocalMux I__6713 (
            .O(N__34625),
            .I(N__34596));
    InMux I__6712 (
            .O(N__34624),
            .I(N__34588));
    InMux I__6711 (
            .O(N__34623),
            .I(N__34588));
    InMux I__6710 (
            .O(N__34622),
            .I(N__34585));
    InMux I__6709 (
            .O(N__34621),
            .I(N__34580));
    LocalMux I__6708 (
            .O(N__34618),
            .I(N__34577));
    LocalMux I__6707 (
            .O(N__34609),
            .I(N__34574));
    Span4Mux_v I__6706 (
            .O(N__34606),
            .I(N__34569));
    Span4Mux_v I__6705 (
            .O(N__34599),
            .I(N__34569));
    Span4Mux_v I__6704 (
            .O(N__34596),
            .I(N__34566));
    InMux I__6703 (
            .O(N__34595),
            .I(N__34563));
    InMux I__6702 (
            .O(N__34594),
            .I(N__34558));
    InMux I__6701 (
            .O(N__34593),
            .I(N__34558));
    LocalMux I__6700 (
            .O(N__34588),
            .I(N__34553));
    LocalMux I__6699 (
            .O(N__34585),
            .I(N__34553));
    InMux I__6698 (
            .O(N__34584),
            .I(N__34548));
    InMux I__6697 (
            .O(N__34583),
            .I(N__34548));
    LocalMux I__6696 (
            .O(N__34580),
            .I(N__34543));
    Span12Mux_s9_v I__6695 (
            .O(N__34577),
            .I(N__34543));
    Span4Mux_h I__6694 (
            .O(N__34574),
            .I(N__34538));
    Span4Mux_v I__6693 (
            .O(N__34569),
            .I(N__34538));
    Span4Mux_h I__6692 (
            .O(N__34566),
            .I(N__34535));
    LocalMux I__6691 (
            .O(N__34563),
            .I(n20590));
    LocalMux I__6690 (
            .O(N__34558),
            .I(n20590));
    Odrv4 I__6689 (
            .O(N__34553),
            .I(n20590));
    LocalMux I__6688 (
            .O(N__34548),
            .I(n20590));
    Odrv12 I__6687 (
            .O(N__34543),
            .I(n20590));
    Odrv4 I__6686 (
            .O(N__34538),
            .I(n20590));
    Odrv4 I__6685 (
            .O(N__34535),
            .I(n20590));
    InMux I__6684 (
            .O(N__34520),
            .I(N__34515));
    InMux I__6683 (
            .O(N__34519),
            .I(N__34512));
    CascadeMux I__6682 (
            .O(N__34518),
            .I(N__34509));
    LocalMux I__6681 (
            .O(N__34515),
            .I(N__34506));
    LocalMux I__6680 (
            .O(N__34512),
            .I(N__34503));
    InMux I__6679 (
            .O(N__34509),
            .I(N__34500));
    Span4Mux_v I__6678 (
            .O(N__34506),
            .I(N__34497));
    Span4Mux_v I__6677 (
            .O(N__34503),
            .I(N__34494));
    LocalMux I__6676 (
            .O(N__34500),
            .I(cmd_rdadctmp_19));
    Odrv4 I__6675 (
            .O(N__34497),
            .I(cmd_rdadctmp_19));
    Odrv4 I__6674 (
            .O(N__34494),
            .I(cmd_rdadctmp_19));
    CascadeMux I__6673 (
            .O(N__34487),
            .I(N__34484));
    InMux I__6672 (
            .O(N__34484),
            .I(N__34479));
    InMux I__6671 (
            .O(N__34483),
            .I(N__34476));
    CascadeMux I__6670 (
            .O(N__34482),
            .I(N__34473));
    LocalMux I__6669 (
            .O(N__34479),
            .I(N__34468));
    LocalMux I__6668 (
            .O(N__34476),
            .I(N__34468));
    InMux I__6667 (
            .O(N__34473),
            .I(N__34465));
    Odrv12 I__6666 (
            .O(N__34468),
            .I(cmd_rdadctmp_25));
    LocalMux I__6665 (
            .O(N__34465),
            .I(cmd_rdadctmp_25));
    CascadeMux I__6664 (
            .O(N__34460),
            .I(N__34457));
    InMux I__6663 (
            .O(N__34457),
            .I(N__34447));
    InMux I__6662 (
            .O(N__34456),
            .I(N__34447));
    InMux I__6661 (
            .O(N__34455),
            .I(N__34444));
    InMux I__6660 (
            .O(N__34454),
            .I(N__34441));
    InMux I__6659 (
            .O(N__34453),
            .I(N__34436));
    InMux I__6658 (
            .O(N__34452),
            .I(N__34433));
    LocalMux I__6657 (
            .O(N__34447),
            .I(N__34419));
    LocalMux I__6656 (
            .O(N__34444),
            .I(N__34419));
    LocalMux I__6655 (
            .O(N__34441),
            .I(N__34416));
    InMux I__6654 (
            .O(N__34440),
            .I(N__34411));
    InMux I__6653 (
            .O(N__34439),
            .I(N__34411));
    LocalMux I__6652 (
            .O(N__34436),
            .I(N__34405));
    LocalMux I__6651 (
            .O(N__34433),
            .I(N__34405));
    InMux I__6650 (
            .O(N__34432),
            .I(N__34402));
    InMux I__6649 (
            .O(N__34431),
            .I(N__34399));
    InMux I__6648 (
            .O(N__34430),
            .I(N__34396));
    InMux I__6647 (
            .O(N__34429),
            .I(N__34393));
    InMux I__6646 (
            .O(N__34428),
            .I(N__34388));
    InMux I__6645 (
            .O(N__34427),
            .I(N__34388));
    InMux I__6644 (
            .O(N__34426),
            .I(N__34383));
    InMux I__6643 (
            .O(N__34425),
            .I(N__34383));
    InMux I__6642 (
            .O(N__34424),
            .I(N__34377));
    Span4Mux_h I__6641 (
            .O(N__34419),
            .I(N__34370));
    Span4Mux_v I__6640 (
            .O(N__34416),
            .I(N__34370));
    LocalMux I__6639 (
            .O(N__34411),
            .I(N__34370));
    InMux I__6638 (
            .O(N__34410),
            .I(N__34367));
    Span4Mux_v I__6637 (
            .O(N__34405),
            .I(N__34362));
    LocalMux I__6636 (
            .O(N__34402),
            .I(N__34362));
    LocalMux I__6635 (
            .O(N__34399),
            .I(N__34357));
    LocalMux I__6634 (
            .O(N__34396),
            .I(N__34357));
    LocalMux I__6633 (
            .O(N__34393),
            .I(N__34350));
    LocalMux I__6632 (
            .O(N__34388),
            .I(N__34350));
    LocalMux I__6631 (
            .O(N__34383),
            .I(N__34350));
    InMux I__6630 (
            .O(N__34382),
            .I(N__34343));
    InMux I__6629 (
            .O(N__34381),
            .I(N__34343));
    InMux I__6628 (
            .O(N__34380),
            .I(N__34343));
    LocalMux I__6627 (
            .O(N__34377),
            .I(N__34340));
    Span4Mux_v I__6626 (
            .O(N__34370),
            .I(N__34329));
    LocalMux I__6625 (
            .O(N__34367),
            .I(N__34326));
    Span4Mux_v I__6624 (
            .O(N__34362),
            .I(N__34317));
    Span4Mux_v I__6623 (
            .O(N__34357),
            .I(N__34317));
    Span4Mux_h I__6622 (
            .O(N__34350),
            .I(N__34317));
    LocalMux I__6621 (
            .O(N__34343),
            .I(N__34317));
    Span4Mux_v I__6620 (
            .O(N__34340),
            .I(N__34314));
    InMux I__6619 (
            .O(N__34339),
            .I(N__34305));
    InMux I__6618 (
            .O(N__34338),
            .I(N__34305));
    InMux I__6617 (
            .O(N__34337),
            .I(N__34305));
    InMux I__6616 (
            .O(N__34336),
            .I(N__34305));
    InMux I__6615 (
            .O(N__34335),
            .I(N__34300));
    InMux I__6614 (
            .O(N__34334),
            .I(N__34300));
    CascadeMux I__6613 (
            .O(N__34333),
            .I(N__34297));
    CascadeMux I__6612 (
            .O(N__34332),
            .I(N__34293));
    Span4Mux_v I__6611 (
            .O(N__34329),
            .I(N__34286));
    Span4Mux_v I__6610 (
            .O(N__34326),
            .I(N__34286));
    Span4Mux_h I__6609 (
            .O(N__34317),
            .I(N__34283));
    Sp12to4 I__6608 (
            .O(N__34314),
            .I(N__34276));
    LocalMux I__6607 (
            .O(N__34305),
            .I(N__34276));
    LocalMux I__6606 (
            .O(N__34300),
            .I(N__34276));
    InMux I__6605 (
            .O(N__34297),
            .I(N__34271));
    InMux I__6604 (
            .O(N__34296),
            .I(N__34271));
    InMux I__6603 (
            .O(N__34293),
            .I(N__34264));
    InMux I__6602 (
            .O(N__34292),
            .I(N__34264));
    InMux I__6601 (
            .O(N__34291),
            .I(N__34264));
    Sp12to4 I__6600 (
            .O(N__34286),
            .I(N__34261));
    Span4Mux_h I__6599 (
            .O(N__34283),
            .I(N__34258));
    Span12Mux_h I__6598 (
            .O(N__34276),
            .I(N__34251));
    LocalMux I__6597 (
            .O(N__34271),
            .I(N__34251));
    LocalMux I__6596 (
            .O(N__34264),
            .I(N__34251));
    Odrv12 I__6595 (
            .O(N__34261),
            .I(n12534));
    Odrv4 I__6594 (
            .O(N__34258),
            .I(n12534));
    Odrv12 I__6593 (
            .O(N__34251),
            .I(n12534));
    CascadeMux I__6592 (
            .O(N__34244),
            .I(N__34241));
    InMux I__6591 (
            .O(N__34241),
            .I(N__34235));
    InMux I__6590 (
            .O(N__34240),
            .I(N__34235));
    LocalMux I__6589 (
            .O(N__34235),
            .I(N__34231));
    CascadeMux I__6588 (
            .O(N__34234),
            .I(N__34228));
    Span4Mux_v I__6587 (
            .O(N__34231),
            .I(N__34225));
    InMux I__6586 (
            .O(N__34228),
            .I(N__34222));
    Odrv4 I__6585 (
            .O(N__34225),
            .I(cmd_rdadctmp_26));
    LocalMux I__6584 (
            .O(N__34222),
            .I(cmd_rdadctmp_26));
    CEMux I__6583 (
            .O(N__34217),
            .I(N__34213));
    CEMux I__6582 (
            .O(N__34216),
            .I(N__34210));
    LocalMux I__6581 (
            .O(N__34213),
            .I(N__34207));
    LocalMux I__6580 (
            .O(N__34210),
            .I(N__34204));
    Span4Mux_h I__6579 (
            .O(N__34207),
            .I(N__34201));
    Span4Mux_v I__6578 (
            .O(N__34204),
            .I(N__34198));
    Odrv4 I__6577 (
            .O(N__34201),
            .I(n12110));
    Odrv4 I__6576 (
            .O(N__34198),
            .I(n12110));
    CascadeMux I__6575 (
            .O(N__34193),
            .I(n12110_cascade_));
    SRMux I__6574 (
            .O(N__34190),
            .I(N__34186));
    SRMux I__6573 (
            .O(N__34189),
            .I(N__34183));
    LocalMux I__6572 (
            .O(N__34186),
            .I(N__34180));
    LocalMux I__6571 (
            .O(N__34183),
            .I(N__34177));
    Span4Mux_h I__6570 (
            .O(N__34180),
            .I(N__34174));
    Span4Mux_v I__6569 (
            .O(N__34177),
            .I(N__34171));
    Odrv4 I__6568 (
            .O(N__34174),
            .I(n14780));
    Odrv4 I__6567 (
            .O(N__34171),
            .I(n14780));
    InMux I__6566 (
            .O(N__34166),
            .I(N__34162));
    CascadeMux I__6565 (
            .O(N__34165),
            .I(N__34159));
    LocalMux I__6564 (
            .O(N__34162),
            .I(N__34156));
    InMux I__6563 (
            .O(N__34159),
            .I(N__34153));
    Span4Mux_h I__6562 (
            .O(N__34156),
            .I(N__34150));
    LocalMux I__6561 (
            .O(N__34153),
            .I(data_idxvec_10));
    Odrv4 I__6560 (
            .O(N__34150),
            .I(data_idxvec_10));
    CascadeMux I__6559 (
            .O(N__34145),
            .I(n20905_cascade_));
    InMux I__6558 (
            .O(N__34142),
            .I(N__34139));
    LocalMux I__6557 (
            .O(N__34139),
            .I(N__34136));
    Span4Mux_v I__6556 (
            .O(N__34136),
            .I(N__34133));
    Span4Mux_h I__6555 (
            .O(N__34133),
            .I(N__34130));
    Odrv4 I__6554 (
            .O(N__34130),
            .I(n20839));
    CascadeMux I__6553 (
            .O(N__34127),
            .I(n22148_cascade_));
    InMux I__6552 (
            .O(N__34124),
            .I(N__34121));
    LocalMux I__6551 (
            .O(N__34121),
            .I(N__34118));
    Span4Mux_h I__6550 (
            .O(N__34118),
            .I(N__34115));
    Odrv4 I__6549 (
            .O(N__34115),
            .I(n22121));
    CascadeMux I__6548 (
            .O(N__34112),
            .I(n22151_cascade_));
    CascadeMux I__6547 (
            .O(N__34109),
            .I(n20889_cascade_));
    InMux I__6546 (
            .O(N__34106),
            .I(N__34103));
    LocalMux I__6545 (
            .O(N__34103),
            .I(N__34100));
    Span4Mux_h I__6544 (
            .O(N__34100),
            .I(N__34097));
    Span4Mux_h I__6543 (
            .O(N__34097),
            .I(N__34094));
    Odrv4 I__6542 (
            .O(N__34094),
            .I(buf_data_iac_18));
    InMux I__6541 (
            .O(N__34091),
            .I(N__34088));
    LocalMux I__6540 (
            .O(N__34088),
            .I(n20906));
    CascadeMux I__6539 (
            .O(N__34085),
            .I(n12152_cascade_));
    CascadeMux I__6538 (
            .O(N__34082),
            .I(N__34079));
    InMux I__6537 (
            .O(N__34079),
            .I(N__34076));
    LocalMux I__6536 (
            .O(N__34076),
            .I(n12_adj_1639));
    CascadeMux I__6535 (
            .O(N__34073),
            .I(n12194_cascade_));
    InMux I__6534 (
            .O(N__34070),
            .I(N__34067));
    LocalMux I__6533 (
            .O(N__34067),
            .I(N__34064));
    Span4Mux_h I__6532 (
            .O(N__34064),
            .I(N__34060));
    InMux I__6531 (
            .O(N__34063),
            .I(N__34057));
    Span4Mux_h I__6530 (
            .O(N__34060),
            .I(N__34052));
    LocalMux I__6529 (
            .O(N__34057),
            .I(N__34052));
    Span4Mux_h I__6528 (
            .O(N__34052),
            .I(N__34048));
    InMux I__6527 (
            .O(N__34051),
            .I(N__34045));
    Span4Mux_v I__6526 (
            .O(N__34048),
            .I(N__34042));
    LocalMux I__6525 (
            .O(N__34045),
            .I(buf_adcdata_iac_0));
    Odrv4 I__6524 (
            .O(N__34042),
            .I(buf_adcdata_iac_0));
    CascadeMux I__6523 (
            .O(N__34037),
            .I(n22_cascade_));
    InMux I__6522 (
            .O(N__34034),
            .I(N__34031));
    LocalMux I__6521 (
            .O(N__34031),
            .I(N__34028));
    Span12Mux_h I__6520 (
            .O(N__34028),
            .I(N__34025));
    Odrv12 I__6519 (
            .O(N__34025),
            .I(buf_data_iac_0));
    CascadeMux I__6518 (
            .O(N__34022),
            .I(n30_adj_1484_cascade_));
    CascadeMux I__6517 (
            .O(N__34019),
            .I(N__34016));
    InMux I__6516 (
            .O(N__34016),
            .I(N__34013));
    LocalMux I__6515 (
            .O(N__34013),
            .I(N__34010));
    Span4Mux_v I__6514 (
            .O(N__34010),
            .I(N__34007));
    Odrv4 I__6513 (
            .O(N__34007),
            .I(n22_adj_1489));
    InMux I__6512 (
            .O(N__34004),
            .I(N__34001));
    LocalMux I__6511 (
            .O(N__34001),
            .I(N__33998));
    Span4Mux_h I__6510 (
            .O(N__33998),
            .I(N__33995));
    Span4Mux_h I__6509 (
            .O(N__33995),
            .I(N__33992));
    Odrv4 I__6508 (
            .O(N__33992),
            .I(buf_data_iac_1));
    CascadeMux I__6507 (
            .O(N__33989),
            .I(n30_adj_1504_cascade_));
    InMux I__6506 (
            .O(N__33986),
            .I(N__33983));
    LocalMux I__6505 (
            .O(N__33983),
            .I(N__33979));
    CascadeMux I__6504 (
            .O(N__33982),
            .I(N__33976));
    Span4Mux_v I__6503 (
            .O(N__33979),
            .I(N__33973));
    InMux I__6502 (
            .O(N__33976),
            .I(N__33970));
    Odrv4 I__6501 (
            .O(N__33973),
            .I(buf_adcdata_vdc_0));
    LocalMux I__6500 (
            .O(N__33970),
            .I(buf_adcdata_vdc_0));
    InMux I__6499 (
            .O(N__33965),
            .I(N__33961));
    InMux I__6498 (
            .O(N__33964),
            .I(N__33958));
    LocalMux I__6497 (
            .O(N__33961),
            .I(N__33954));
    LocalMux I__6496 (
            .O(N__33958),
            .I(N__33951));
    CascadeMux I__6495 (
            .O(N__33957),
            .I(N__33948));
    Span4Mux_v I__6494 (
            .O(N__33954),
            .I(N__33945));
    Span12Mux_v I__6493 (
            .O(N__33951),
            .I(N__33942));
    InMux I__6492 (
            .O(N__33948),
            .I(N__33939));
    Span4Mux_h I__6491 (
            .O(N__33945),
            .I(N__33936));
    Span12Mux_h I__6490 (
            .O(N__33942),
            .I(N__33933));
    LocalMux I__6489 (
            .O(N__33939),
            .I(buf_adcdata_vac_0));
    Odrv4 I__6488 (
            .O(N__33936),
            .I(buf_adcdata_vac_0));
    Odrv12 I__6487 (
            .O(N__33933),
            .I(buf_adcdata_vac_0));
    InMux I__6486 (
            .O(N__33926),
            .I(N__33923));
    LocalMux I__6485 (
            .O(N__33923),
            .I(n19_adj_1485));
    InMux I__6484 (
            .O(N__33920),
            .I(\ADC_VDC.genclk.n19494 ));
    InMux I__6483 (
            .O(N__33917),
            .I(\ADC_VDC.genclk.n19495 ));
    InMux I__6482 (
            .O(N__33914),
            .I(\ADC_VDC.genclk.n19496 ));
    InMux I__6481 (
            .O(N__33911),
            .I(\ADC_VDC.genclk.n19497 ));
    CEMux I__6480 (
            .O(N__33908),
            .I(N__33904));
    CEMux I__6479 (
            .O(N__33907),
            .I(N__33901));
    LocalMux I__6478 (
            .O(N__33904),
            .I(N__33898));
    LocalMux I__6477 (
            .O(N__33901),
            .I(N__33895));
    Span4Mux_v I__6476 (
            .O(N__33898),
            .I(N__33892));
    Span4Mux_v I__6475 (
            .O(N__33895),
            .I(N__33889));
    Span4Mux_h I__6474 (
            .O(N__33892),
            .I(N__33886));
    Odrv4 I__6473 (
            .O(N__33889),
            .I(\ADC_VDC.genclk.div_state_1__N_1275 ));
    Odrv4 I__6472 (
            .O(N__33886),
            .I(\ADC_VDC.genclk.div_state_1__N_1275 ));
    SRMux I__6471 (
            .O(N__33881),
            .I(N__33877));
    SRMux I__6470 (
            .O(N__33880),
            .I(N__33874));
    LocalMux I__6469 (
            .O(N__33877),
            .I(N__33869));
    LocalMux I__6468 (
            .O(N__33874),
            .I(N__33866));
    SRMux I__6467 (
            .O(N__33873),
            .I(N__33863));
    SRMux I__6466 (
            .O(N__33872),
            .I(N__33860));
    Span4Mux_h I__6465 (
            .O(N__33869),
            .I(N__33857));
    Span4Mux_h I__6464 (
            .O(N__33866),
            .I(N__33850));
    LocalMux I__6463 (
            .O(N__33863),
            .I(N__33850));
    LocalMux I__6462 (
            .O(N__33860),
            .I(N__33850));
    Odrv4 I__6461 (
            .O(N__33857),
            .I(\ADC_VDC.genclk.n15067 ));
    Odrv4 I__6460 (
            .O(N__33850),
            .I(\ADC_VDC.genclk.n15067 ));
    InMux I__6459 (
            .O(N__33845),
            .I(N__33841));
    InMux I__6458 (
            .O(N__33844),
            .I(N__33837));
    LocalMux I__6457 (
            .O(N__33841),
            .I(N__33834));
    InMux I__6456 (
            .O(N__33840),
            .I(N__33831));
    LocalMux I__6455 (
            .O(N__33837),
            .I(N__33824));
    Span4Mux_v I__6454 (
            .O(N__33834),
            .I(N__33824));
    LocalMux I__6453 (
            .O(N__33831),
            .I(N__33824));
    Span4Mux_h I__6452 (
            .O(N__33824),
            .I(N__33820));
    InMux I__6451 (
            .O(N__33823),
            .I(N__33817));
    Span4Mux_v I__6450 (
            .O(N__33820),
            .I(N__33814));
    LocalMux I__6449 (
            .O(N__33817),
            .I(\RTD.bit_cnt_3 ));
    Odrv4 I__6448 (
            .O(N__33814),
            .I(\RTD.bit_cnt_3 ));
    InMux I__6447 (
            .O(N__33809),
            .I(N__33799));
    InMux I__6446 (
            .O(N__33808),
            .I(N__33799));
    InMux I__6445 (
            .O(N__33807),
            .I(N__33799));
    InMux I__6444 (
            .O(N__33806),
            .I(N__33796));
    LocalMux I__6443 (
            .O(N__33799),
            .I(\RTD.bit_cnt_1 ));
    LocalMux I__6442 (
            .O(N__33796),
            .I(\RTD.bit_cnt_1 ));
    InMux I__6441 (
            .O(N__33791),
            .I(N__33784));
    InMux I__6440 (
            .O(N__33790),
            .I(N__33784));
    InMux I__6439 (
            .O(N__33789),
            .I(N__33781));
    LocalMux I__6438 (
            .O(N__33784),
            .I(\RTD.bit_cnt_2 ));
    LocalMux I__6437 (
            .O(N__33781),
            .I(\RTD.bit_cnt_2 ));
    CascadeMux I__6436 (
            .O(N__33776),
            .I(N__33772));
    CascadeMux I__6435 (
            .O(N__33775),
            .I(N__33769));
    InMux I__6434 (
            .O(N__33772),
            .I(N__33757));
    InMux I__6433 (
            .O(N__33769),
            .I(N__33757));
    InMux I__6432 (
            .O(N__33768),
            .I(N__33757));
    InMux I__6431 (
            .O(N__33767),
            .I(N__33757));
    InMux I__6430 (
            .O(N__33766),
            .I(N__33754));
    LocalMux I__6429 (
            .O(N__33757),
            .I(\RTD.bit_cnt_0 ));
    LocalMux I__6428 (
            .O(N__33754),
            .I(\RTD.bit_cnt_0 ));
    CEMux I__6427 (
            .O(N__33749),
            .I(N__33746));
    LocalMux I__6426 (
            .O(N__33746),
            .I(N__33743));
    Span4Mux_h I__6425 (
            .O(N__33743),
            .I(N__33740));
    Span4Mux_h I__6424 (
            .O(N__33740),
            .I(N__33737));
    Span4Mux_h I__6423 (
            .O(N__33737),
            .I(N__33734));
    Odrv4 I__6422 (
            .O(N__33734),
            .I(\RTD.n11756 ));
    SRMux I__6421 (
            .O(N__33731),
            .I(N__33728));
    LocalMux I__6420 (
            .O(N__33728),
            .I(N__33725));
    Span4Mux_h I__6419 (
            .O(N__33725),
            .I(N__33722));
    Span4Mux_h I__6418 (
            .O(N__33722),
            .I(N__33719));
    Span4Mux_h I__6417 (
            .O(N__33719),
            .I(N__33716));
    Odrv4 I__6416 (
            .O(N__33716),
            .I(\RTD.n15081 ));
    InMux I__6415 (
            .O(N__33713),
            .I(\ADC_VDC.genclk.n19485 ));
    InMux I__6414 (
            .O(N__33710),
            .I(\ADC_VDC.genclk.n19486 ));
    InMux I__6413 (
            .O(N__33707),
            .I(\ADC_VDC.genclk.n19487 ));
    InMux I__6412 (
            .O(N__33704),
            .I(\ADC_VDC.genclk.n19488 ));
    InMux I__6411 (
            .O(N__33701),
            .I(\ADC_VDC.genclk.n19489 ));
    InMux I__6410 (
            .O(N__33698),
            .I(bfn_13_6_0_));
    InMux I__6409 (
            .O(N__33695),
            .I(\ADC_VDC.genclk.n19491 ));
    InMux I__6408 (
            .O(N__33692),
            .I(\ADC_VDC.genclk.n19492 ));
    InMux I__6407 (
            .O(N__33689),
            .I(\ADC_VDC.genclk.n19493 ));
    CEMux I__6406 (
            .O(N__33686),
            .I(N__33683));
    LocalMux I__6405 (
            .O(N__33683),
            .I(N__33680));
    Odrv4 I__6404 (
            .O(N__33680),
            .I(\ADC_VDC.genclk.n6 ));
    InMux I__6403 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__6402 (
            .O(N__33674),
            .I(N__33670));
    InMux I__6401 (
            .O(N__33673),
            .I(N__33664));
    Span4Mux_h I__6400 (
            .O(N__33670),
            .I(N__33661));
    InMux I__6399 (
            .O(N__33669),
            .I(N__33654));
    InMux I__6398 (
            .O(N__33668),
            .I(N__33654));
    InMux I__6397 (
            .O(N__33667),
            .I(N__33654));
    LocalMux I__6396 (
            .O(N__33664),
            .I(\ADC_VDC.genclk.div_state_0 ));
    Odrv4 I__6395 (
            .O(N__33661),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__6394 (
            .O(N__33654),
            .I(\ADC_VDC.genclk.div_state_0 ));
    CEMux I__6393 (
            .O(N__33647),
            .I(N__33644));
    LocalMux I__6392 (
            .O(N__33644),
            .I(N__33641));
    Span4Mux_h I__6391 (
            .O(N__33641),
            .I(N__33638));
    Span4Mux_h I__6390 (
            .O(N__33638),
            .I(N__33635));
    Odrv4 I__6389 (
            .O(N__33635),
            .I(\ADC_VDC.n11766 ));
    CascadeMux I__6388 (
            .O(N__33632),
            .I(N__33625));
    CascadeMux I__6387 (
            .O(N__33631),
            .I(N__33622));
    InMux I__6386 (
            .O(N__33630),
            .I(N__33618));
    CascadeMux I__6385 (
            .O(N__33629),
            .I(N__33615));
    InMux I__6384 (
            .O(N__33628),
            .I(N__33603));
    InMux I__6383 (
            .O(N__33625),
            .I(N__33603));
    InMux I__6382 (
            .O(N__33622),
            .I(N__33603));
    InMux I__6381 (
            .O(N__33621),
            .I(N__33603));
    LocalMux I__6380 (
            .O(N__33618),
            .I(N__33600));
    InMux I__6379 (
            .O(N__33615),
            .I(N__33597));
    CascadeMux I__6378 (
            .O(N__33614),
            .I(N__33594));
    InMux I__6377 (
            .O(N__33613),
            .I(N__33589));
    InMux I__6376 (
            .O(N__33612),
            .I(N__33589));
    LocalMux I__6375 (
            .O(N__33603),
            .I(N__33585));
    Span4Mux_v I__6374 (
            .O(N__33600),
            .I(N__33582));
    LocalMux I__6373 (
            .O(N__33597),
            .I(N__33579));
    InMux I__6372 (
            .O(N__33594),
            .I(N__33576));
    LocalMux I__6371 (
            .O(N__33589),
            .I(N__33573));
    InMux I__6370 (
            .O(N__33588),
            .I(N__33570));
    Span4Mux_v I__6369 (
            .O(N__33585),
            .I(N__33567));
    Span4Mux_h I__6368 (
            .O(N__33582),
            .I(N__33560));
    Span4Mux_v I__6367 (
            .O(N__33579),
            .I(N__33560));
    LocalMux I__6366 (
            .O(N__33576),
            .I(N__33560));
    Span4Mux_v I__6365 (
            .O(N__33573),
            .I(N__33555));
    LocalMux I__6364 (
            .O(N__33570),
            .I(N__33555));
    Span4Mux_v I__6363 (
            .O(N__33567),
            .I(N__33552));
    Span4Mux_v I__6362 (
            .O(N__33560),
            .I(N__33549));
    Span4Mux_v I__6361 (
            .O(N__33555),
            .I(N__33546));
    Span4Mux_h I__6360 (
            .O(N__33552),
            .I(N__33543));
    Span4Mux_h I__6359 (
            .O(N__33549),
            .I(N__33540));
    Span4Mux_h I__6358 (
            .O(N__33546),
            .I(N__33537));
    Sp12to4 I__6357 (
            .O(N__33543),
            .I(N__33532));
    Sp12to4 I__6356 (
            .O(N__33540),
            .I(N__33532));
    Span4Mux_h I__6355 (
            .O(N__33537),
            .I(N__33529));
    Odrv12 I__6354 (
            .O(N__33532),
            .I(VDC_SDO));
    Odrv4 I__6353 (
            .O(N__33529),
            .I(VDC_SDO));
    InMux I__6352 (
            .O(N__33524),
            .I(N__33511));
    InMux I__6351 (
            .O(N__33523),
            .I(N__33508));
    InMux I__6350 (
            .O(N__33522),
            .I(N__33505));
    InMux I__6349 (
            .O(N__33521),
            .I(N__33502));
    CascadeMux I__6348 (
            .O(N__33520),
            .I(N__33499));
    InMux I__6347 (
            .O(N__33519),
            .I(N__33494));
    InMux I__6346 (
            .O(N__33518),
            .I(N__33494));
    InMux I__6345 (
            .O(N__33517),
            .I(N__33488));
    InMux I__6344 (
            .O(N__33516),
            .I(N__33481));
    InMux I__6343 (
            .O(N__33515),
            .I(N__33481));
    InMux I__6342 (
            .O(N__33514),
            .I(N__33481));
    LocalMux I__6341 (
            .O(N__33511),
            .I(N__33478));
    LocalMux I__6340 (
            .O(N__33508),
            .I(N__33468));
    LocalMux I__6339 (
            .O(N__33505),
            .I(N__33465));
    LocalMux I__6338 (
            .O(N__33502),
            .I(N__33462));
    InMux I__6337 (
            .O(N__33499),
            .I(N__33459));
    LocalMux I__6336 (
            .O(N__33494),
            .I(N__33456));
    InMux I__6335 (
            .O(N__33493),
            .I(N__33451));
    InMux I__6334 (
            .O(N__33492),
            .I(N__33451));
    InMux I__6333 (
            .O(N__33491),
            .I(N__33448));
    LocalMux I__6332 (
            .O(N__33488),
            .I(N__33443));
    LocalMux I__6331 (
            .O(N__33481),
            .I(N__33443));
    Span4Mux_h I__6330 (
            .O(N__33478),
            .I(N__33440));
    InMux I__6329 (
            .O(N__33477),
            .I(N__33437));
    InMux I__6328 (
            .O(N__33476),
            .I(N__33432));
    InMux I__6327 (
            .O(N__33475),
            .I(N__33432));
    InMux I__6326 (
            .O(N__33474),
            .I(N__33429));
    InMux I__6325 (
            .O(N__33473),
            .I(N__33426));
    InMux I__6324 (
            .O(N__33472),
            .I(N__33421));
    InMux I__6323 (
            .O(N__33471),
            .I(N__33421));
    Span4Mux_v I__6322 (
            .O(N__33468),
            .I(N__33412));
    Span4Mux_v I__6321 (
            .O(N__33465),
            .I(N__33412));
    Span4Mux_h I__6320 (
            .O(N__33462),
            .I(N__33412));
    LocalMux I__6319 (
            .O(N__33459),
            .I(N__33412));
    Span4Mux_h I__6318 (
            .O(N__33456),
            .I(N__33409));
    LocalMux I__6317 (
            .O(N__33451),
            .I(N__33400));
    LocalMux I__6316 (
            .O(N__33448),
            .I(N__33400));
    Span4Mux_h I__6315 (
            .O(N__33443),
            .I(N__33400));
    Span4Mux_h I__6314 (
            .O(N__33440),
            .I(N__33400));
    LocalMux I__6313 (
            .O(N__33437),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6312 (
            .O(N__33432),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6311 (
            .O(N__33429),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6310 (
            .O(N__33426),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6309 (
            .O(N__33421),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__6308 (
            .O(N__33412),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__6307 (
            .O(N__33409),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__6306 (
            .O(N__33400),
            .I(\ADC_VDC.adc_state_0 ));
    CascadeMux I__6305 (
            .O(N__33383),
            .I(N__33380));
    InMux I__6304 (
            .O(N__33380),
            .I(N__33377));
    LocalMux I__6303 (
            .O(N__33377),
            .I(\ADC_VDC.n62 ));
    CascadeMux I__6302 (
            .O(N__33374),
            .I(N__33368));
    CascadeMux I__6301 (
            .O(N__33373),
            .I(N__33359));
    InMux I__6300 (
            .O(N__33372),
            .I(N__33355));
    CascadeMux I__6299 (
            .O(N__33371),
            .I(N__33351));
    InMux I__6298 (
            .O(N__33368),
            .I(N__33341));
    InMux I__6297 (
            .O(N__33367),
            .I(N__33322));
    InMux I__6296 (
            .O(N__33366),
            .I(N__33322));
    InMux I__6295 (
            .O(N__33365),
            .I(N__33322));
    InMux I__6294 (
            .O(N__33364),
            .I(N__33322));
    InMux I__6293 (
            .O(N__33363),
            .I(N__33322));
    InMux I__6292 (
            .O(N__33362),
            .I(N__33322));
    InMux I__6291 (
            .O(N__33359),
            .I(N__33322));
    CascadeMux I__6290 (
            .O(N__33358),
            .I(N__33319));
    LocalMux I__6289 (
            .O(N__33355),
            .I(N__33316));
    InMux I__6288 (
            .O(N__33354),
            .I(N__33311));
    InMux I__6287 (
            .O(N__33351),
            .I(N__33311));
    InMux I__6286 (
            .O(N__33350),
            .I(N__33302));
    InMux I__6285 (
            .O(N__33349),
            .I(N__33302));
    InMux I__6284 (
            .O(N__33348),
            .I(N__33302));
    InMux I__6283 (
            .O(N__33347),
            .I(N__33302));
    InMux I__6282 (
            .O(N__33346),
            .I(N__33286));
    InMux I__6281 (
            .O(N__33345),
            .I(N__33286));
    InMux I__6280 (
            .O(N__33344),
            .I(N__33280));
    LocalMux I__6279 (
            .O(N__33341),
            .I(N__33277));
    CascadeMux I__6278 (
            .O(N__33340),
            .I(N__33274));
    InMux I__6277 (
            .O(N__33339),
            .I(N__33267));
    InMux I__6276 (
            .O(N__33338),
            .I(N__33262));
    InMux I__6275 (
            .O(N__33337),
            .I(N__33262));
    LocalMux I__6274 (
            .O(N__33322),
            .I(N__33259));
    InMux I__6273 (
            .O(N__33319),
            .I(N__33256));
    Span4Mux_h I__6272 (
            .O(N__33316),
            .I(N__33249));
    LocalMux I__6271 (
            .O(N__33311),
            .I(N__33249));
    LocalMux I__6270 (
            .O(N__33302),
            .I(N__33249));
    InMux I__6269 (
            .O(N__33301),
            .I(N__33246));
    InMux I__6268 (
            .O(N__33300),
            .I(N__33241));
    InMux I__6267 (
            .O(N__33299),
            .I(N__33241));
    InMux I__6266 (
            .O(N__33298),
            .I(N__33217));
    InMux I__6265 (
            .O(N__33297),
            .I(N__33217));
    InMux I__6264 (
            .O(N__33296),
            .I(N__33217));
    InMux I__6263 (
            .O(N__33295),
            .I(N__33217));
    InMux I__6262 (
            .O(N__33294),
            .I(N__33217));
    InMux I__6261 (
            .O(N__33293),
            .I(N__33217));
    InMux I__6260 (
            .O(N__33292),
            .I(N__33217));
    InMux I__6259 (
            .O(N__33291),
            .I(N__33217));
    LocalMux I__6258 (
            .O(N__33286),
            .I(N__33214));
    InMux I__6257 (
            .O(N__33285),
            .I(N__33207));
    InMux I__6256 (
            .O(N__33284),
            .I(N__33207));
    InMux I__6255 (
            .O(N__33283),
            .I(N__33207));
    LocalMux I__6254 (
            .O(N__33280),
            .I(N__33202));
    Span4Mux_v I__6253 (
            .O(N__33277),
            .I(N__33202));
    InMux I__6252 (
            .O(N__33274),
            .I(N__33191));
    InMux I__6251 (
            .O(N__33273),
            .I(N__33191));
    InMux I__6250 (
            .O(N__33272),
            .I(N__33191));
    InMux I__6249 (
            .O(N__33271),
            .I(N__33191));
    InMux I__6248 (
            .O(N__33270),
            .I(N__33191));
    LocalMux I__6247 (
            .O(N__33267),
            .I(N__33180));
    LocalMux I__6246 (
            .O(N__33262),
            .I(N__33180));
    Span4Mux_h I__6245 (
            .O(N__33259),
            .I(N__33180));
    LocalMux I__6244 (
            .O(N__33256),
            .I(N__33180));
    Span4Mux_h I__6243 (
            .O(N__33249),
            .I(N__33180));
    LocalMux I__6242 (
            .O(N__33246),
            .I(N__33175));
    LocalMux I__6241 (
            .O(N__33241),
            .I(N__33175));
    InMux I__6240 (
            .O(N__33240),
            .I(N__33172));
    InMux I__6239 (
            .O(N__33239),
            .I(N__33167));
    InMux I__6238 (
            .O(N__33238),
            .I(N__33167));
    InMux I__6237 (
            .O(N__33237),
            .I(N__33164));
    InMux I__6236 (
            .O(N__33236),
            .I(N__33157));
    InMux I__6235 (
            .O(N__33235),
            .I(N__33157));
    InMux I__6234 (
            .O(N__33234),
            .I(N__33157));
    LocalMux I__6233 (
            .O(N__33217),
            .I(N__33146));
    Span4Mux_h I__6232 (
            .O(N__33214),
            .I(N__33146));
    LocalMux I__6231 (
            .O(N__33207),
            .I(N__33146));
    Span4Mux_h I__6230 (
            .O(N__33202),
            .I(N__33146));
    LocalMux I__6229 (
            .O(N__33191),
            .I(N__33146));
    Span4Mux_v I__6228 (
            .O(N__33180),
            .I(N__33141));
    Span4Mux_h I__6227 (
            .O(N__33175),
            .I(N__33141));
    LocalMux I__6226 (
            .O(N__33172),
            .I(adc_state_2));
    LocalMux I__6225 (
            .O(N__33167),
            .I(adc_state_2));
    LocalMux I__6224 (
            .O(N__33164),
            .I(adc_state_2));
    LocalMux I__6223 (
            .O(N__33157),
            .I(adc_state_2));
    Odrv4 I__6222 (
            .O(N__33146),
            .I(adc_state_2));
    Odrv4 I__6221 (
            .O(N__33141),
            .I(adc_state_2));
    CascadeMux I__6220 (
            .O(N__33128),
            .I(N__33105));
    CascadeMux I__6219 (
            .O(N__33127),
            .I(N__33102));
    CascadeMux I__6218 (
            .O(N__33126),
            .I(N__33093));
    InMux I__6217 (
            .O(N__33125),
            .I(N__33090));
    CascadeMux I__6216 (
            .O(N__33124),
            .I(N__33087));
    InMux I__6215 (
            .O(N__33123),
            .I(N__33076));
    InMux I__6214 (
            .O(N__33122),
            .I(N__33076));
    InMux I__6213 (
            .O(N__33121),
            .I(N__33063));
    InMux I__6212 (
            .O(N__33120),
            .I(N__33063));
    InMux I__6211 (
            .O(N__33119),
            .I(N__33063));
    InMux I__6210 (
            .O(N__33118),
            .I(N__33063));
    InMux I__6209 (
            .O(N__33117),
            .I(N__33063));
    InMux I__6208 (
            .O(N__33116),
            .I(N__33063));
    InMux I__6207 (
            .O(N__33115),
            .I(N__33046));
    InMux I__6206 (
            .O(N__33114),
            .I(N__33046));
    InMux I__6205 (
            .O(N__33113),
            .I(N__33046));
    InMux I__6204 (
            .O(N__33112),
            .I(N__33046));
    InMux I__6203 (
            .O(N__33111),
            .I(N__33046));
    InMux I__6202 (
            .O(N__33110),
            .I(N__33046));
    InMux I__6201 (
            .O(N__33109),
            .I(N__33046));
    InMux I__6200 (
            .O(N__33108),
            .I(N__33046));
    InMux I__6199 (
            .O(N__33105),
            .I(N__33035));
    InMux I__6198 (
            .O(N__33102),
            .I(N__33035));
    InMux I__6197 (
            .O(N__33101),
            .I(N__33035));
    InMux I__6196 (
            .O(N__33100),
            .I(N__33028));
    InMux I__6195 (
            .O(N__33099),
            .I(N__33028));
    InMux I__6194 (
            .O(N__33098),
            .I(N__33028));
    InMux I__6193 (
            .O(N__33097),
            .I(N__33023));
    InMux I__6192 (
            .O(N__33096),
            .I(N__33023));
    InMux I__6191 (
            .O(N__33093),
            .I(N__33019));
    LocalMux I__6190 (
            .O(N__33090),
            .I(N__33016));
    InMux I__6189 (
            .O(N__33087),
            .I(N__33013));
    InMux I__6188 (
            .O(N__33086),
            .I(N__33008));
    InMux I__6187 (
            .O(N__33085),
            .I(N__32997));
    InMux I__6186 (
            .O(N__33084),
            .I(N__32997));
    InMux I__6185 (
            .O(N__33083),
            .I(N__32997));
    InMux I__6184 (
            .O(N__33082),
            .I(N__32997));
    InMux I__6183 (
            .O(N__33081),
            .I(N__32997));
    LocalMux I__6182 (
            .O(N__33076),
            .I(N__32994));
    LocalMux I__6181 (
            .O(N__33063),
            .I(N__32989));
    LocalMux I__6180 (
            .O(N__33046),
            .I(N__32989));
    InMux I__6179 (
            .O(N__33045),
            .I(N__32974));
    InMux I__6178 (
            .O(N__33044),
            .I(N__32974));
    InMux I__6177 (
            .O(N__33043),
            .I(N__32974));
    InMux I__6176 (
            .O(N__33042),
            .I(N__32974));
    LocalMux I__6175 (
            .O(N__33035),
            .I(N__32967));
    LocalMux I__6174 (
            .O(N__33028),
            .I(N__32967));
    LocalMux I__6173 (
            .O(N__33023),
            .I(N__32967));
    InMux I__6172 (
            .O(N__33022),
            .I(N__32964));
    LocalMux I__6171 (
            .O(N__33019),
            .I(N__32961));
    Span4Mux_h I__6170 (
            .O(N__33016),
            .I(N__32956));
    LocalMux I__6169 (
            .O(N__33013),
            .I(N__32956));
    InMux I__6168 (
            .O(N__33012),
            .I(N__32951));
    InMux I__6167 (
            .O(N__33011),
            .I(N__32951));
    LocalMux I__6166 (
            .O(N__33008),
            .I(N__32942));
    LocalMux I__6165 (
            .O(N__32997),
            .I(N__32942));
    Span4Mux_v I__6164 (
            .O(N__32994),
            .I(N__32942));
    Span4Mux_v I__6163 (
            .O(N__32989),
            .I(N__32942));
    InMux I__6162 (
            .O(N__32988),
            .I(N__32929));
    InMux I__6161 (
            .O(N__32987),
            .I(N__32929));
    InMux I__6160 (
            .O(N__32986),
            .I(N__32929));
    InMux I__6159 (
            .O(N__32985),
            .I(N__32929));
    InMux I__6158 (
            .O(N__32984),
            .I(N__32929));
    InMux I__6157 (
            .O(N__32983),
            .I(N__32929));
    LocalMux I__6156 (
            .O(N__32974),
            .I(N__32924));
    Span12Mux_h I__6155 (
            .O(N__32967),
            .I(N__32924));
    LocalMux I__6154 (
            .O(N__32964),
            .I(adc_state_3));
    Odrv4 I__6153 (
            .O(N__32961),
            .I(adc_state_3));
    Odrv4 I__6152 (
            .O(N__32956),
            .I(adc_state_3));
    LocalMux I__6151 (
            .O(N__32951),
            .I(adc_state_3));
    Odrv4 I__6150 (
            .O(N__32942),
            .I(adc_state_3));
    LocalMux I__6149 (
            .O(N__32929),
            .I(adc_state_3));
    Odrv12 I__6148 (
            .O(N__32924),
            .I(adc_state_3));
    CascadeMux I__6147 (
            .O(N__32909),
            .I(\ADC_VDC.n62_cascade_ ));
    CascadeMux I__6146 (
            .O(N__32906),
            .I(N__32899));
    InMux I__6145 (
            .O(N__32905),
            .I(N__32887));
    InMux I__6144 (
            .O(N__32904),
            .I(N__32887));
    InMux I__6143 (
            .O(N__32903),
            .I(N__32887));
    InMux I__6142 (
            .O(N__32902),
            .I(N__32884));
    InMux I__6141 (
            .O(N__32899),
            .I(N__32879));
    InMux I__6140 (
            .O(N__32898),
            .I(N__32879));
    InMux I__6139 (
            .O(N__32897),
            .I(N__32876));
    InMux I__6138 (
            .O(N__32896),
            .I(N__32873));
    InMux I__6137 (
            .O(N__32895),
            .I(N__32861));
    InMux I__6136 (
            .O(N__32894),
            .I(N__32861));
    LocalMux I__6135 (
            .O(N__32887),
            .I(N__32852));
    LocalMux I__6134 (
            .O(N__32884),
            .I(N__32852));
    LocalMux I__6133 (
            .O(N__32879),
            .I(N__32847));
    LocalMux I__6132 (
            .O(N__32876),
            .I(N__32847));
    LocalMux I__6131 (
            .O(N__32873),
            .I(N__32842));
    InMux I__6130 (
            .O(N__32872),
            .I(N__32835));
    InMux I__6129 (
            .O(N__32871),
            .I(N__32835));
    InMux I__6128 (
            .O(N__32870),
            .I(N__32835));
    InMux I__6127 (
            .O(N__32869),
            .I(N__32832));
    InMux I__6126 (
            .O(N__32868),
            .I(N__32829));
    InMux I__6125 (
            .O(N__32867),
            .I(N__32824));
    InMux I__6124 (
            .O(N__32866),
            .I(N__32824));
    LocalMux I__6123 (
            .O(N__32861),
            .I(N__32821));
    InMux I__6122 (
            .O(N__32860),
            .I(N__32818));
    InMux I__6121 (
            .O(N__32859),
            .I(N__32815));
    InMux I__6120 (
            .O(N__32858),
            .I(N__32810));
    InMux I__6119 (
            .O(N__32857),
            .I(N__32810));
    Span4Mux_h I__6118 (
            .O(N__32852),
            .I(N__32807));
    Span4Mux_h I__6117 (
            .O(N__32847),
            .I(N__32804));
    InMux I__6116 (
            .O(N__32846),
            .I(N__32799));
    InMux I__6115 (
            .O(N__32845),
            .I(N__32799));
    Span4Mux_h I__6114 (
            .O(N__32842),
            .I(N__32794));
    LocalMux I__6113 (
            .O(N__32835),
            .I(N__32794));
    LocalMux I__6112 (
            .O(N__32832),
            .I(N__32785));
    LocalMux I__6111 (
            .O(N__32829),
            .I(N__32785));
    LocalMux I__6110 (
            .O(N__32824),
            .I(N__32785));
    Span12Mux_v I__6109 (
            .O(N__32821),
            .I(N__32785));
    LocalMux I__6108 (
            .O(N__32818),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6107 (
            .O(N__32815),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6106 (
            .O(N__32810),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6105 (
            .O(N__32807),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6104 (
            .O(N__32804),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6103 (
            .O(N__32799),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6102 (
            .O(N__32794),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv12 I__6101 (
            .O(N__32785),
            .I(\ADC_VDC.adc_state_1 ));
    InMux I__6100 (
            .O(N__32768),
            .I(N__32765));
    LocalMux I__6099 (
            .O(N__32765),
            .I(N__32762));
    Span4Mux_h I__6098 (
            .O(N__32762),
            .I(N__32759));
    Span4Mux_h I__6097 (
            .O(N__32759),
            .I(N__32756));
    Odrv4 I__6096 (
            .O(N__32756),
            .I(\ADC_VDC.n11 ));
    InMux I__6095 (
            .O(N__32753),
            .I(bfn_13_5_0_));
    InMux I__6094 (
            .O(N__32750),
            .I(\ADC_VDC.genclk.n19483 ));
    InMux I__6093 (
            .O(N__32747),
            .I(\ADC_VDC.genclk.n19484 ));
    InMux I__6092 (
            .O(N__32744),
            .I(n19383));
    IoInMux I__6091 (
            .O(N__32741),
            .I(N__32738));
    LocalMux I__6090 (
            .O(N__32738),
            .I(N__32735));
    Span12Mux_s7_v I__6089 (
            .O(N__32735),
            .I(N__32730));
    ClkMux I__6088 (
            .O(N__32734),
            .I(N__32727));
    ClkMux I__6087 (
            .O(N__32733),
            .I(N__32724));
    Span12Mux_v I__6086 (
            .O(N__32730),
            .I(N__32721));
    LocalMux I__6085 (
            .O(N__32727),
            .I(N__32718));
    LocalMux I__6084 (
            .O(N__32724),
            .I(N__32715));
    Span12Mux_h I__6083 (
            .O(N__32721),
            .I(N__32711));
    Span4Mux_v I__6082 (
            .O(N__32718),
            .I(N__32708));
    Span4Mux_h I__6081 (
            .O(N__32715),
            .I(N__32705));
    InMux I__6080 (
            .O(N__32714),
            .I(N__32702));
    Odrv12 I__6079 (
            .O(N__32711),
            .I(TEST_LED));
    Odrv4 I__6078 (
            .O(N__32708),
            .I(TEST_LED));
    Odrv4 I__6077 (
            .O(N__32705),
            .I(TEST_LED));
    LocalMux I__6076 (
            .O(N__32702),
            .I(TEST_LED));
    CascadeMux I__6075 (
            .O(N__32693),
            .I(N__32690));
    InMux I__6074 (
            .O(N__32690),
            .I(N__32686));
    InMux I__6073 (
            .O(N__32689),
            .I(N__32683));
    LocalMux I__6072 (
            .O(N__32686),
            .I(\ADC_VDC.genclk.t0off_13 ));
    LocalMux I__6071 (
            .O(N__32683),
            .I(\ADC_VDC.genclk.t0off_13 ));
    InMux I__6070 (
            .O(N__32678),
            .I(N__32674));
    InMux I__6069 (
            .O(N__32677),
            .I(N__32671));
    LocalMux I__6068 (
            .O(N__32674),
            .I(\ADC_VDC.genclk.t0off_3 ));
    LocalMux I__6067 (
            .O(N__32671),
            .I(\ADC_VDC.genclk.t0off_3 ));
    CascadeMux I__6066 (
            .O(N__32666),
            .I(N__32662));
    InMux I__6065 (
            .O(N__32665),
            .I(N__32659));
    InMux I__6064 (
            .O(N__32662),
            .I(N__32656));
    LocalMux I__6063 (
            .O(N__32659),
            .I(\ADC_VDC.genclk.t0off_5 ));
    LocalMux I__6062 (
            .O(N__32656),
            .I(\ADC_VDC.genclk.t0off_5 ));
    InMux I__6061 (
            .O(N__32651),
            .I(N__32647));
    InMux I__6060 (
            .O(N__32650),
            .I(N__32644));
    LocalMux I__6059 (
            .O(N__32647),
            .I(\ADC_VDC.genclk.t0off_8 ));
    LocalMux I__6058 (
            .O(N__32644),
            .I(\ADC_VDC.genclk.t0off_8 ));
    InMux I__6057 (
            .O(N__32639),
            .I(N__32636));
    LocalMux I__6056 (
            .O(N__32636),
            .I(N__32633));
    Odrv4 I__6055 (
            .O(N__32633),
            .I(\ADC_VDC.genclk.n27 ));
    CascadeMux I__6054 (
            .O(N__32630),
            .I(\ADC_VDC.genclk.n26_cascade_ ));
    CascadeMux I__6053 (
            .O(N__32627),
            .I(\ADC_VDC.genclk.n21206_cascade_ ));
    CascadeMux I__6052 (
            .O(N__32624),
            .I(N__32621));
    InMux I__6051 (
            .O(N__32621),
            .I(N__32617));
    InMux I__6050 (
            .O(N__32620),
            .I(N__32614));
    LocalMux I__6049 (
            .O(N__32617),
            .I(\ADC_VDC.genclk.t0off_6 ));
    LocalMux I__6048 (
            .O(N__32614),
            .I(\ADC_VDC.genclk.t0off_6 ));
    InMux I__6047 (
            .O(N__32609),
            .I(N__32605));
    InMux I__6046 (
            .O(N__32608),
            .I(N__32602));
    LocalMux I__6045 (
            .O(N__32605),
            .I(\ADC_VDC.genclk.t0off_0 ));
    LocalMux I__6044 (
            .O(N__32602),
            .I(\ADC_VDC.genclk.t0off_0 ));
    CascadeMux I__6043 (
            .O(N__32597),
            .I(N__32593));
    CascadeMux I__6042 (
            .O(N__32596),
            .I(N__32590));
    InMux I__6041 (
            .O(N__32593),
            .I(N__32587));
    InMux I__6040 (
            .O(N__32590),
            .I(N__32584));
    LocalMux I__6039 (
            .O(N__32587),
            .I(\ADC_VDC.genclk.t0off_4 ));
    LocalMux I__6038 (
            .O(N__32584),
            .I(\ADC_VDC.genclk.t0off_4 ));
    InMux I__6037 (
            .O(N__32579),
            .I(N__32575));
    InMux I__6036 (
            .O(N__32578),
            .I(N__32572));
    LocalMux I__6035 (
            .O(N__32575),
            .I(\ADC_VDC.genclk.t0off_1 ));
    LocalMux I__6034 (
            .O(N__32572),
            .I(\ADC_VDC.genclk.t0off_1 ));
    InMux I__6033 (
            .O(N__32567),
            .I(N__32564));
    LocalMux I__6032 (
            .O(N__32564),
            .I(\ADC_VDC.genclk.n21208 ));
    InMux I__6031 (
            .O(N__32561),
            .I(N__32557));
    InMux I__6030 (
            .O(N__32560),
            .I(N__32554));
    LocalMux I__6029 (
            .O(N__32557),
            .I(\ADC_VDC.genclk.t0off_14 ));
    LocalMux I__6028 (
            .O(N__32554),
            .I(\ADC_VDC.genclk.t0off_14 ));
    CascadeMux I__6027 (
            .O(N__32549),
            .I(N__32546));
    InMux I__6026 (
            .O(N__32546),
            .I(N__32542));
    InMux I__6025 (
            .O(N__32545),
            .I(N__32539));
    LocalMux I__6024 (
            .O(N__32542),
            .I(\ADC_VDC.genclk.t0off_9 ));
    LocalMux I__6023 (
            .O(N__32539),
            .I(\ADC_VDC.genclk.t0off_9 ));
    CascadeMux I__6022 (
            .O(N__32534),
            .I(N__32530));
    InMux I__6021 (
            .O(N__32533),
            .I(N__32527));
    InMux I__6020 (
            .O(N__32530),
            .I(N__32524));
    LocalMux I__6019 (
            .O(N__32527),
            .I(\ADC_VDC.genclk.t0off_15 ));
    LocalMux I__6018 (
            .O(N__32524),
            .I(\ADC_VDC.genclk.t0off_15 ));
    CascadeMux I__6017 (
            .O(N__32519),
            .I(N__32516));
    InMux I__6016 (
            .O(N__32516),
            .I(N__32512));
    InMux I__6015 (
            .O(N__32515),
            .I(N__32509));
    LocalMux I__6014 (
            .O(N__32512),
            .I(\ADC_VDC.genclk.t0off_11 ));
    LocalMux I__6013 (
            .O(N__32509),
            .I(\ADC_VDC.genclk.t0off_11 ));
    InMux I__6012 (
            .O(N__32504),
            .I(N__32501));
    LocalMux I__6011 (
            .O(N__32501),
            .I(\ADC_VDC.genclk.n28 ));
    InMux I__6010 (
            .O(N__32498),
            .I(N__32495));
    LocalMux I__6009 (
            .O(N__32495),
            .I(\ADC_VDC.genclk.n21206 ));
    InMux I__6008 (
            .O(N__32492),
            .I(n19375));
    InMux I__6007 (
            .O(N__32489),
            .I(n19376));
    InMux I__6006 (
            .O(N__32486),
            .I(bfn_12_18_0_));
    InMux I__6005 (
            .O(N__32483),
            .I(N__32479));
    InMux I__6004 (
            .O(N__32482),
            .I(N__32476));
    LocalMux I__6003 (
            .O(N__32479),
            .I(N__32473));
    LocalMux I__6002 (
            .O(N__32476),
            .I(acadc_skipcnt_10));
    Odrv4 I__6001 (
            .O(N__32473),
            .I(acadc_skipcnt_10));
    InMux I__6000 (
            .O(N__32468),
            .I(n19378));
    InMux I__5999 (
            .O(N__32465),
            .I(N__32461));
    InMux I__5998 (
            .O(N__32464),
            .I(N__32458));
    LocalMux I__5997 (
            .O(N__32461),
            .I(N__32455));
    LocalMux I__5996 (
            .O(N__32458),
            .I(acadc_skipcnt_11));
    Odrv4 I__5995 (
            .O(N__32455),
            .I(acadc_skipcnt_11));
    InMux I__5994 (
            .O(N__32450),
            .I(n19379));
    InMux I__5993 (
            .O(N__32447),
            .I(N__32443));
    InMux I__5992 (
            .O(N__32446),
            .I(N__32440));
    LocalMux I__5991 (
            .O(N__32443),
            .I(N__32437));
    LocalMux I__5990 (
            .O(N__32440),
            .I(acadc_skipcnt_12));
    Odrv4 I__5989 (
            .O(N__32437),
            .I(acadc_skipcnt_12));
    InMux I__5988 (
            .O(N__32432),
            .I(n19380));
    InMux I__5987 (
            .O(N__32429),
            .I(n19381));
    InMux I__5986 (
            .O(N__32426),
            .I(N__32422));
    InMux I__5985 (
            .O(N__32425),
            .I(N__32419));
    LocalMux I__5984 (
            .O(N__32422),
            .I(N__32416));
    LocalMux I__5983 (
            .O(N__32419),
            .I(acadc_skipcnt_14));
    Odrv4 I__5982 (
            .O(N__32416),
            .I(acadc_skipcnt_14));
    InMux I__5981 (
            .O(N__32411),
            .I(n19382));
    InMux I__5980 (
            .O(N__32408),
            .I(bfn_12_17_0_));
    InMux I__5979 (
            .O(N__32405),
            .I(n19370));
    InMux I__5978 (
            .O(N__32402),
            .I(n19371));
    InMux I__5977 (
            .O(N__32399),
            .I(n19372));
    InMux I__5976 (
            .O(N__32396),
            .I(n19373));
    CascadeMux I__5975 (
            .O(N__32393),
            .I(N__32390));
    InMux I__5974 (
            .O(N__32390),
            .I(N__32386));
    InMux I__5973 (
            .O(N__32389),
            .I(N__32383));
    LocalMux I__5972 (
            .O(N__32386),
            .I(N__32380));
    LocalMux I__5971 (
            .O(N__32383),
            .I(acadc_skipcnt_6));
    Odrv4 I__5970 (
            .O(N__32380),
            .I(acadc_skipcnt_6));
    InMux I__5969 (
            .O(N__32375),
            .I(n19374));
    InMux I__5968 (
            .O(N__32372),
            .I(N__32368));
    CascadeMux I__5967 (
            .O(N__32371),
            .I(N__32365));
    LocalMux I__5966 (
            .O(N__32368),
            .I(N__32362));
    InMux I__5965 (
            .O(N__32365),
            .I(N__32358));
    Span12Mux_v I__5964 (
            .O(N__32362),
            .I(N__32355));
    InMux I__5963 (
            .O(N__32361),
            .I(N__32352));
    LocalMux I__5962 (
            .O(N__32358),
            .I(acadc_skipCount_14));
    Odrv12 I__5961 (
            .O(N__32355),
            .I(acadc_skipCount_14));
    LocalMux I__5960 (
            .O(N__32352),
            .I(acadc_skipCount_14));
    InMux I__5959 (
            .O(N__32345),
            .I(N__32342));
    LocalMux I__5958 (
            .O(N__32342),
            .I(N__32339));
    Span4Mux_v I__5957 (
            .O(N__32339),
            .I(N__32334));
    InMux I__5956 (
            .O(N__32338),
            .I(N__32329));
    InMux I__5955 (
            .O(N__32337),
            .I(N__32329));
    Odrv4 I__5954 (
            .O(N__32334),
            .I(acadc_skipCount_10));
    LocalMux I__5953 (
            .O(N__32329),
            .I(acadc_skipCount_10));
    CascadeMux I__5952 (
            .O(N__32324),
            .I(N__32321));
    InMux I__5951 (
            .O(N__32321),
            .I(N__32317));
    InMux I__5950 (
            .O(N__32320),
            .I(N__32314));
    LocalMux I__5949 (
            .O(N__32317),
            .I(acadc_skipcnt_0));
    LocalMux I__5948 (
            .O(N__32314),
            .I(acadc_skipcnt_0));
    CascadeMux I__5947 (
            .O(N__32309),
            .I(n16594_cascade_));
    InMux I__5946 (
            .O(N__32306),
            .I(N__32303));
    LocalMux I__5945 (
            .O(N__32303),
            .I(n22196));
    CascadeMux I__5944 (
            .O(N__32300),
            .I(n16602_cascade_));
    InMux I__5943 (
            .O(N__32297),
            .I(N__32294));
    LocalMux I__5942 (
            .O(N__32294),
            .I(n16602));
    InMux I__5941 (
            .O(N__32291),
            .I(n19407));
    CascadeMux I__5940 (
            .O(N__32288),
            .I(n22169_cascade_));
    InMux I__5939 (
            .O(N__32285),
            .I(N__32282));
    LocalMux I__5938 (
            .O(N__32282),
            .I(N__32279));
    Span4Mux_h I__5937 (
            .O(N__32279),
            .I(N__32276));
    Span4Mux_v I__5936 (
            .O(N__32276),
            .I(N__32273));
    Odrv4 I__5935 (
            .O(N__32273),
            .I(n22079));
    CascadeMux I__5934 (
            .O(N__32270),
            .I(n20568_cascade_));
    InMux I__5933 (
            .O(N__32267),
            .I(N__32263));
    InMux I__5932 (
            .O(N__32266),
            .I(N__32260));
    LocalMux I__5931 (
            .O(N__32263),
            .I(data_idxvec_15));
    LocalMux I__5930 (
            .O(N__32260),
            .I(data_idxvec_15));
    InMux I__5929 (
            .O(N__32255),
            .I(N__32251));
    InMux I__5928 (
            .O(N__32254),
            .I(N__32248));
    LocalMux I__5927 (
            .O(N__32251),
            .I(eis_end));
    LocalMux I__5926 (
            .O(N__32248),
            .I(eis_end));
    CascadeMux I__5925 (
            .O(N__32243),
            .I(n26_adj_1528_cascade_));
    InMux I__5924 (
            .O(N__32240),
            .I(N__32237));
    LocalMux I__5923 (
            .O(N__32237),
            .I(n22166));
    InMux I__5922 (
            .O(N__32234),
            .I(N__32231));
    LocalMux I__5921 (
            .O(N__32231),
            .I(n20742));
    InMux I__5920 (
            .O(N__32228),
            .I(N__32221));
    InMux I__5919 (
            .O(N__32227),
            .I(N__32221));
    InMux I__5918 (
            .O(N__32226),
            .I(N__32218));
    LocalMux I__5917 (
            .O(N__32221),
            .I(N__32214));
    LocalMux I__5916 (
            .O(N__32218),
            .I(N__32210));
    CascadeMux I__5915 (
            .O(N__32217),
            .I(N__32207));
    Span4Mux_v I__5914 (
            .O(N__32214),
            .I(N__32204));
    InMux I__5913 (
            .O(N__32213),
            .I(N__32201));
    Span4Mux_h I__5912 (
            .O(N__32210),
            .I(N__32198));
    InMux I__5911 (
            .O(N__32207),
            .I(N__32195));
    Span4Mux_h I__5910 (
            .O(N__32204),
            .I(N__32192));
    LocalMux I__5909 (
            .O(N__32201),
            .I(N__32189));
    Span4Mux_h I__5908 (
            .O(N__32198),
            .I(N__32186));
    LocalMux I__5907 (
            .O(N__32195),
            .I(N__32181));
    Span4Mux_h I__5906 (
            .O(N__32192),
            .I(N__32181));
    Odrv12 I__5905 (
            .O(N__32189),
            .I(acadc_trig));
    Odrv4 I__5904 (
            .O(N__32186),
            .I(acadc_trig));
    Odrv4 I__5903 (
            .O(N__32181),
            .I(acadc_trig));
    InMux I__5902 (
            .O(N__32174),
            .I(n19398));
    InMux I__5901 (
            .O(N__32171),
            .I(n19399));
    InMux I__5900 (
            .O(N__32168),
            .I(bfn_12_12_0_));
    InMux I__5899 (
            .O(N__32165),
            .I(n19401));
    InMux I__5898 (
            .O(N__32162),
            .I(n19402));
    InMux I__5897 (
            .O(N__32159),
            .I(n19403));
    InMux I__5896 (
            .O(N__32156),
            .I(n19404));
    CascadeMux I__5895 (
            .O(N__32153),
            .I(N__32150));
    InMux I__5894 (
            .O(N__32150),
            .I(N__32146));
    CascadeMux I__5893 (
            .O(N__32149),
            .I(N__32143));
    LocalMux I__5892 (
            .O(N__32146),
            .I(N__32140));
    InMux I__5891 (
            .O(N__32143),
            .I(N__32137));
    Span4Mux_h I__5890 (
            .O(N__32140),
            .I(N__32134));
    LocalMux I__5889 (
            .O(N__32137),
            .I(data_idxvec_13));
    Odrv4 I__5888 (
            .O(N__32134),
            .I(data_idxvec_13));
    InMux I__5887 (
            .O(N__32129),
            .I(n19405));
    InMux I__5886 (
            .O(N__32126),
            .I(n19406));
    CascadeMux I__5885 (
            .O(N__32123),
            .I(N__32117));
    InMux I__5884 (
            .O(N__32122),
            .I(N__32113));
    InMux I__5883 (
            .O(N__32121),
            .I(N__32110));
    InMux I__5882 (
            .O(N__32120),
            .I(N__32105));
    InMux I__5881 (
            .O(N__32117),
            .I(N__32105));
    CascadeMux I__5880 (
            .O(N__32116),
            .I(N__32102));
    LocalMux I__5879 (
            .O(N__32113),
            .I(N__32096));
    LocalMux I__5878 (
            .O(N__32110),
            .I(N__32091));
    LocalMux I__5877 (
            .O(N__32105),
            .I(N__32091));
    InMux I__5876 (
            .O(N__32102),
            .I(N__32086));
    InMux I__5875 (
            .O(N__32101),
            .I(N__32086));
    InMux I__5874 (
            .O(N__32100),
            .I(N__32083));
    InMux I__5873 (
            .O(N__32099),
            .I(N__32080));
    Span4Mux_v I__5872 (
            .O(N__32096),
            .I(N__32077));
    Span4Mux_h I__5871 (
            .O(N__32091),
            .I(N__32074));
    LocalMux I__5870 (
            .O(N__32086),
            .I(N__32071));
    LocalMux I__5869 (
            .O(N__32083),
            .I(N__32068));
    LocalMux I__5868 (
            .O(N__32080),
            .I(N__32065));
    Odrv4 I__5867 (
            .O(N__32077),
            .I(n14522));
    Odrv4 I__5866 (
            .O(N__32074),
            .I(n14522));
    Odrv4 I__5865 (
            .O(N__32071),
            .I(n14522));
    Odrv4 I__5864 (
            .O(N__32068),
            .I(n14522));
    Odrv12 I__5863 (
            .O(N__32065),
            .I(n14522));
    InMux I__5862 (
            .O(N__32054),
            .I(N__32050));
    InMux I__5861 (
            .O(N__32053),
            .I(N__32047));
    LocalMux I__5860 (
            .O(N__32050),
            .I(N__32041));
    LocalMux I__5859 (
            .O(N__32047),
            .I(N__32038));
    InMux I__5858 (
            .O(N__32046),
            .I(N__32033));
    InMux I__5857 (
            .O(N__32045),
            .I(N__32033));
    CascadeMux I__5856 (
            .O(N__32044),
            .I(N__32029));
    Span4Mux_v I__5855 (
            .O(N__32041),
            .I(N__32020));
    Span4Mux_h I__5854 (
            .O(N__32038),
            .I(N__32020));
    LocalMux I__5853 (
            .O(N__32033),
            .I(N__32020));
    InMux I__5852 (
            .O(N__32032),
            .I(N__32013));
    InMux I__5851 (
            .O(N__32029),
            .I(N__32013));
    InMux I__5850 (
            .O(N__32028),
            .I(N__32013));
    InMux I__5849 (
            .O(N__32027),
            .I(N__32010));
    Odrv4 I__5848 (
            .O(N__32020),
            .I(n11918));
    LocalMux I__5847 (
            .O(N__32013),
            .I(n11918));
    LocalMux I__5846 (
            .O(N__32010),
            .I(n11918));
    CascadeMux I__5845 (
            .O(N__32003),
            .I(N__31998));
    InMux I__5844 (
            .O(N__32002),
            .I(N__31995));
    InMux I__5843 (
            .O(N__32001),
            .I(N__31990));
    InMux I__5842 (
            .O(N__31998),
            .I(N__31990));
    LocalMux I__5841 (
            .O(N__31995),
            .I(cmd_rdadctmp_22));
    LocalMux I__5840 (
            .O(N__31990),
            .I(cmd_rdadctmp_22));
    InMux I__5839 (
            .O(N__31985),
            .I(bfn_12_11_0_));
    InMux I__5838 (
            .O(N__31982),
            .I(n19393));
    InMux I__5837 (
            .O(N__31979),
            .I(n19394));
    InMux I__5836 (
            .O(N__31976),
            .I(n19395));
    InMux I__5835 (
            .O(N__31973),
            .I(n19396));
    InMux I__5834 (
            .O(N__31970),
            .I(n19397));
    InMux I__5833 (
            .O(N__31967),
            .I(N__31962));
    InMux I__5832 (
            .O(N__31966),
            .I(N__31959));
    CascadeMux I__5831 (
            .O(N__31965),
            .I(N__31956));
    LocalMux I__5830 (
            .O(N__31962),
            .I(N__31953));
    LocalMux I__5829 (
            .O(N__31959),
            .I(N__31950));
    InMux I__5828 (
            .O(N__31956),
            .I(N__31947));
    Span4Mux_v I__5827 (
            .O(N__31953),
            .I(N__31944));
    Span4Mux_v I__5826 (
            .O(N__31950),
            .I(N__31941));
    LocalMux I__5825 (
            .O(N__31947),
            .I(N__31936));
    Sp12to4 I__5824 (
            .O(N__31944),
            .I(N__31936));
    Span4Mux_h I__5823 (
            .O(N__31941),
            .I(N__31933));
    Odrv12 I__5822 (
            .O(N__31936),
            .I(buf_adcdata_vac_22));
    Odrv4 I__5821 (
            .O(N__31933),
            .I(buf_adcdata_vac_22));
    CascadeMux I__5820 (
            .O(N__31928),
            .I(N__31925));
    InMux I__5819 (
            .O(N__31925),
            .I(N__31921));
    InMux I__5818 (
            .O(N__31924),
            .I(N__31918));
    LocalMux I__5817 (
            .O(N__31921),
            .I(buf_adcdata_vdc_22));
    LocalMux I__5816 (
            .O(N__31918),
            .I(buf_adcdata_vdc_22));
    InMux I__5815 (
            .O(N__31913),
            .I(N__31910));
    LocalMux I__5814 (
            .O(N__31910),
            .I(N__31907));
    Odrv4 I__5813 (
            .O(N__31907),
            .I(n22160));
    InMux I__5812 (
            .O(N__31904),
            .I(N__31900));
    InMux I__5811 (
            .O(N__31903),
            .I(N__31897));
    LocalMux I__5810 (
            .O(N__31900),
            .I(N__31894));
    LocalMux I__5809 (
            .O(N__31897),
            .I(comm_buf_6_4));
    Odrv4 I__5808 (
            .O(N__31894),
            .I(comm_buf_6_4));
    InMux I__5807 (
            .O(N__31889),
            .I(N__31886));
    LocalMux I__5806 (
            .O(N__31886),
            .I(N__31883));
    Span4Mux_h I__5805 (
            .O(N__31883),
            .I(N__31877));
    InMux I__5804 (
            .O(N__31882),
            .I(N__31874));
    InMux I__5803 (
            .O(N__31881),
            .I(N__31869));
    InMux I__5802 (
            .O(N__31880),
            .I(N__31869));
    Odrv4 I__5801 (
            .O(N__31877),
            .I(n20646));
    LocalMux I__5800 (
            .O(N__31874),
            .I(n20646));
    LocalMux I__5799 (
            .O(N__31869),
            .I(n20646));
    InMux I__5798 (
            .O(N__31862),
            .I(N__31859));
    LocalMux I__5797 (
            .O(N__31859),
            .I(N__31856));
    Span4Mux_h I__5796 (
            .O(N__31856),
            .I(N__31853));
    Odrv4 I__5795 (
            .O(N__31853),
            .I(n30_adj_1630));
    InMux I__5794 (
            .O(N__31850),
            .I(N__31847));
    LocalMux I__5793 (
            .O(N__31847),
            .I(N__31844));
    Span4Mux_v I__5792 (
            .O(N__31844),
            .I(N__31841));
    Odrv4 I__5791 (
            .O(N__31841),
            .I(n30_adj_1634));
    InMux I__5790 (
            .O(N__31838),
            .I(N__31835));
    LocalMux I__5789 (
            .O(N__31835),
            .I(N__31832));
    Span4Mux_h I__5788 (
            .O(N__31832),
            .I(N__31829));
    Span4Mux_v I__5787 (
            .O(N__31829),
            .I(N__31826));
    Odrv4 I__5786 (
            .O(N__31826),
            .I(n30_adj_1638));
    InMux I__5785 (
            .O(N__31823),
            .I(N__31820));
    LocalMux I__5784 (
            .O(N__31820),
            .I(comm_buf_2_4));
    InMux I__5783 (
            .O(N__31817),
            .I(N__31814));
    LocalMux I__5782 (
            .O(N__31814),
            .I(N__31811));
    Span4Mux_v I__5781 (
            .O(N__31811),
            .I(N__31808));
    Odrv4 I__5780 (
            .O(N__31808),
            .I(n30_adj_1644));
    InMux I__5779 (
            .O(N__31805),
            .I(N__31802));
    LocalMux I__5778 (
            .O(N__31802),
            .I(N__31799));
    Span4Mux_v I__5777 (
            .O(N__31799),
            .I(N__31796));
    Odrv4 I__5776 (
            .O(N__31796),
            .I(n30_adj_1648));
    InMux I__5775 (
            .O(N__31793),
            .I(N__31790));
    LocalMux I__5774 (
            .O(N__31790),
            .I(N__31786));
    CascadeMux I__5773 (
            .O(N__31789),
            .I(N__31783));
    Span4Mux_h I__5772 (
            .O(N__31786),
            .I(N__31779));
    InMux I__5771 (
            .O(N__31783),
            .I(N__31776));
    InMux I__5770 (
            .O(N__31782),
            .I(N__31773));
    Sp12to4 I__5769 (
            .O(N__31779),
            .I(N__31768));
    LocalMux I__5768 (
            .O(N__31776),
            .I(N__31768));
    LocalMux I__5767 (
            .O(N__31773),
            .I(cmd_rdadctmp_22_adj_1457));
    Odrv12 I__5766 (
            .O(N__31768),
            .I(cmd_rdadctmp_22_adj_1457));
    InMux I__5765 (
            .O(N__31763),
            .I(N__31760));
    LocalMux I__5764 (
            .O(N__31760),
            .I(N__31757));
    Span4Mux_h I__5763 (
            .O(N__31757),
            .I(N__31754));
    Odrv4 I__5762 (
            .O(N__31754),
            .I(\ADC_VDC.n10552 ));
    CascadeMux I__5761 (
            .O(N__31751),
            .I(N__31748));
    InMux I__5760 (
            .O(N__31748),
            .I(N__31745));
    LocalMux I__5759 (
            .O(N__31745),
            .I(N__31741));
    CascadeMux I__5758 (
            .O(N__31744),
            .I(N__31738));
    Span4Mux_v I__5757 (
            .O(N__31741),
            .I(N__31735));
    InMux I__5756 (
            .O(N__31738),
            .I(N__31732));
    Span4Mux_h I__5755 (
            .O(N__31735),
            .I(N__31729));
    LocalMux I__5754 (
            .O(N__31732),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    Odrv4 I__5753 (
            .O(N__31729),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    CEMux I__5752 (
            .O(N__31724),
            .I(N__31721));
    LocalMux I__5751 (
            .O(N__31721),
            .I(\ADC_VDC.n12915 ));
    SRMux I__5750 (
            .O(N__31718),
            .I(N__31715));
    LocalMux I__5749 (
            .O(N__31715),
            .I(N__31712));
    Span4Mux_v I__5748 (
            .O(N__31712),
            .I(N__31709));
    Span4Mux_h I__5747 (
            .O(N__31709),
            .I(N__31706));
    Odrv4 I__5746 (
            .O(N__31706),
            .I(\ADC_VDC.n20392 ));
    InMux I__5745 (
            .O(N__31703),
            .I(N__31698));
    InMux I__5744 (
            .O(N__31702),
            .I(N__31695));
    InMux I__5743 (
            .O(N__31701),
            .I(N__31692));
    LocalMux I__5742 (
            .O(N__31698),
            .I(N__31689));
    LocalMux I__5741 (
            .O(N__31695),
            .I(N__31684));
    LocalMux I__5740 (
            .O(N__31692),
            .I(N__31684));
    Span4Mux_h I__5739 (
            .O(N__31689),
            .I(N__31679));
    Span4Mux_v I__5738 (
            .O(N__31684),
            .I(N__31679));
    Span4Mux_h I__5737 (
            .O(N__31679),
            .I(N__31676));
    Odrv4 I__5736 (
            .O(N__31676),
            .I(\RTD.n17720 ));
    SRMux I__5735 (
            .O(N__31673),
            .I(N__31670));
    LocalMux I__5734 (
            .O(N__31670),
            .I(N__31666));
    SRMux I__5733 (
            .O(N__31669),
            .I(N__31663));
    Span4Mux_v I__5732 (
            .O(N__31666),
            .I(N__31658));
    LocalMux I__5731 (
            .O(N__31663),
            .I(N__31658));
    Odrv4 I__5730 (
            .O(N__31658),
            .I(n14801));
    CascadeMux I__5729 (
            .O(N__31655),
            .I(n2_adj_1587_cascade_));
    InMux I__5728 (
            .O(N__31652),
            .I(N__31649));
    LocalMux I__5727 (
            .O(N__31649),
            .I(comm_buf_5_4));
    InMux I__5726 (
            .O(N__31646),
            .I(N__31643));
    LocalMux I__5725 (
            .O(N__31643),
            .I(n21324));
    CascadeMux I__5724 (
            .O(N__31640),
            .I(n4_adj_1588_cascade_));
    InMux I__5723 (
            .O(N__31637),
            .I(N__31634));
    LocalMux I__5722 (
            .O(N__31634),
            .I(n22136));
    InMux I__5721 (
            .O(N__31631),
            .I(N__31628));
    LocalMux I__5720 (
            .O(N__31628),
            .I(n1_adj_1586));
    InMux I__5719 (
            .O(N__31625),
            .I(N__31622));
    LocalMux I__5718 (
            .O(N__31622),
            .I(n19006));
    CascadeMux I__5717 (
            .O(N__31619),
            .I(n19006_cascade_));
    InMux I__5716 (
            .O(N__31616),
            .I(N__31613));
    LocalMux I__5715 (
            .O(N__31613),
            .I(N__31610));
    Span12Mux_h I__5714 (
            .O(N__31610),
            .I(N__31607));
    Odrv12 I__5713 (
            .O(N__31607),
            .I(n30_adj_1627));
    InMux I__5712 (
            .O(N__31604),
            .I(\ADC_VDC.genclk.n19482 ));
    CEMux I__5711 (
            .O(N__31601),
            .I(N__31598));
    LocalMux I__5710 (
            .O(N__31598),
            .I(N__31594));
    CEMux I__5709 (
            .O(N__31597),
            .I(N__31591));
    Span4Mux_v I__5708 (
            .O(N__31594),
            .I(N__31588));
    LocalMux I__5707 (
            .O(N__31591),
            .I(N__31585));
    Span4Mux_h I__5706 (
            .O(N__31588),
            .I(N__31580));
    Span4Mux_v I__5705 (
            .O(N__31585),
            .I(N__31580));
    Odrv4 I__5704 (
            .O(N__31580),
            .I(\ADC_VDC.genclk.n11751 ));
    CascadeMux I__5703 (
            .O(N__31577),
            .I(n12_adj_1615_cascade_));
    CascadeMux I__5702 (
            .O(N__31574),
            .I(n12236_cascade_));
    InMux I__5701 (
            .O(N__31571),
            .I(N__31568));
    LocalMux I__5700 (
            .O(N__31568),
            .I(N__31565));
    Span4Mux_v I__5699 (
            .O(N__31565),
            .I(N__31562));
    Sp12to4 I__5698 (
            .O(N__31562),
            .I(N__31559));
    Odrv12 I__5697 (
            .O(N__31559),
            .I(buf_data_vac_0));
    InMux I__5696 (
            .O(N__31556),
            .I(N__31553));
    LocalMux I__5695 (
            .O(N__31553),
            .I(N__31550));
    Span4Mux_h I__5694 (
            .O(N__31550),
            .I(N__31547));
    Span4Mux_h I__5693 (
            .O(N__31547),
            .I(N__31544));
    Span4Mux_h I__5692 (
            .O(N__31544),
            .I(N__31541));
    Odrv4 I__5691 (
            .O(N__31541),
            .I(buf_data_vac_1));
    InMux I__5690 (
            .O(N__31538),
            .I(N__31535));
    LocalMux I__5689 (
            .O(N__31535),
            .I(N__31532));
    Span4Mux_v I__5688 (
            .O(N__31532),
            .I(N__31529));
    Sp12to4 I__5687 (
            .O(N__31529),
            .I(N__31526));
    Odrv12 I__5686 (
            .O(N__31526),
            .I(buf_data_vac_2));
    InMux I__5685 (
            .O(N__31523),
            .I(N__31520));
    LocalMux I__5684 (
            .O(N__31520),
            .I(N__31517));
    Span4Mux_h I__5683 (
            .O(N__31517),
            .I(N__31514));
    Span4Mux_h I__5682 (
            .O(N__31514),
            .I(N__31511));
    Odrv4 I__5681 (
            .O(N__31511),
            .I(buf_data_vac_3));
    InMux I__5680 (
            .O(N__31508),
            .I(N__31505));
    LocalMux I__5679 (
            .O(N__31505),
            .I(N__31502));
    Span4Mux_h I__5678 (
            .O(N__31502),
            .I(N__31499));
    Span4Mux_h I__5677 (
            .O(N__31499),
            .I(N__31496));
    Odrv4 I__5676 (
            .O(N__31496),
            .I(buf_data_vac_4));
    CEMux I__5675 (
            .O(N__31493),
            .I(N__31490));
    LocalMux I__5674 (
            .O(N__31490),
            .I(N__31486));
    CEMux I__5673 (
            .O(N__31489),
            .I(N__31483));
    Span4Mux_v I__5672 (
            .O(N__31486),
            .I(N__31478));
    LocalMux I__5671 (
            .O(N__31483),
            .I(N__31478));
    Odrv4 I__5670 (
            .O(N__31478),
            .I(n12236));
    InMux I__5669 (
            .O(N__31475),
            .I(\ADC_VDC.genclk.n19473 ));
    CascadeMux I__5668 (
            .O(N__31472),
            .I(N__31468));
    InMux I__5667 (
            .O(N__31471),
            .I(N__31465));
    InMux I__5666 (
            .O(N__31468),
            .I(N__31462));
    LocalMux I__5665 (
            .O(N__31465),
            .I(\ADC_VDC.genclk.t0off_7 ));
    LocalMux I__5664 (
            .O(N__31462),
            .I(\ADC_VDC.genclk.t0off_7 ));
    InMux I__5663 (
            .O(N__31457),
            .I(\ADC_VDC.genclk.n19474 ));
    InMux I__5662 (
            .O(N__31454),
            .I(bfn_12_4_0_));
    InMux I__5661 (
            .O(N__31451),
            .I(\ADC_VDC.genclk.n19476 ));
    InMux I__5660 (
            .O(N__31448),
            .I(N__31444));
    InMux I__5659 (
            .O(N__31447),
            .I(N__31441));
    LocalMux I__5658 (
            .O(N__31444),
            .I(\ADC_VDC.genclk.t0off_10 ));
    LocalMux I__5657 (
            .O(N__31441),
            .I(\ADC_VDC.genclk.t0off_10 ));
    InMux I__5656 (
            .O(N__31436),
            .I(\ADC_VDC.genclk.n19477 ));
    InMux I__5655 (
            .O(N__31433),
            .I(\ADC_VDC.genclk.n19478 ));
    InMux I__5654 (
            .O(N__31430),
            .I(N__31426));
    InMux I__5653 (
            .O(N__31429),
            .I(N__31423));
    LocalMux I__5652 (
            .O(N__31426),
            .I(\ADC_VDC.genclk.t0off_12 ));
    LocalMux I__5651 (
            .O(N__31423),
            .I(\ADC_VDC.genclk.t0off_12 ));
    InMux I__5650 (
            .O(N__31418),
            .I(\ADC_VDC.genclk.n19479 ));
    InMux I__5649 (
            .O(N__31415),
            .I(\ADC_VDC.genclk.n19480 ));
    InMux I__5648 (
            .O(N__31412),
            .I(\ADC_VDC.genclk.n19481 ));
    CascadeMux I__5647 (
            .O(N__31409),
            .I(N__31406));
    InMux I__5646 (
            .O(N__31406),
            .I(N__31403));
    LocalMux I__5645 (
            .O(N__31403),
            .I(\SIG_DDS.tmp_buf_0 ));
    CEMux I__5644 (
            .O(N__31400),
            .I(N__31397));
    LocalMux I__5643 (
            .O(N__31397),
            .I(N__31394));
    Span4Mux_v I__5642 (
            .O(N__31394),
            .I(N__31391));
    Span4Mux_h I__5641 (
            .O(N__31391),
            .I(N__31386));
    CEMux I__5640 (
            .O(N__31390),
            .I(N__31383));
    CEMux I__5639 (
            .O(N__31389),
            .I(N__31380));
    Odrv4 I__5638 (
            .O(N__31386),
            .I(\SIG_DDS.n12738 ));
    LocalMux I__5637 (
            .O(N__31383),
            .I(\SIG_DDS.n12738 ));
    LocalMux I__5636 (
            .O(N__31380),
            .I(\SIG_DDS.n12738 ));
    InMux I__5635 (
            .O(N__31373),
            .I(N__31370));
    LocalMux I__5634 (
            .O(N__31370),
            .I(N__31366));
    InMux I__5633 (
            .O(N__31369),
            .I(N__31363));
    Span4Mux_h I__5632 (
            .O(N__31366),
            .I(N__31360));
    LocalMux I__5631 (
            .O(N__31363),
            .I(N__31357));
    Span4Mux_v I__5630 (
            .O(N__31360),
            .I(N__31354));
    Span12Mux_h I__5629 (
            .O(N__31357),
            .I(N__31351));
    Odrv4 I__5628 (
            .O(N__31354),
            .I(EIS_SYNCCLK));
    Odrv12 I__5627 (
            .O(N__31351),
            .I(EIS_SYNCCLK));
    IoInMux I__5626 (
            .O(N__31346),
            .I(N__31343));
    LocalMux I__5625 (
            .O(N__31343),
            .I(N__31340));
    Span4Mux_s3_v I__5624 (
            .O(N__31340),
            .I(N__31337));
    Odrv4 I__5623 (
            .O(N__31337),
            .I(OUT_SYNCCLK));
    InMux I__5622 (
            .O(N__31334),
            .I(bfn_12_3_0_));
    InMux I__5621 (
            .O(N__31331),
            .I(\ADC_VDC.genclk.n19468 ));
    CascadeMux I__5620 (
            .O(N__31328),
            .I(N__31325));
    InMux I__5619 (
            .O(N__31325),
            .I(N__31321));
    InMux I__5618 (
            .O(N__31324),
            .I(N__31318));
    LocalMux I__5617 (
            .O(N__31321),
            .I(\ADC_VDC.genclk.t0off_2 ));
    LocalMux I__5616 (
            .O(N__31318),
            .I(\ADC_VDC.genclk.t0off_2 ));
    InMux I__5615 (
            .O(N__31313),
            .I(\ADC_VDC.genclk.n19469 ));
    InMux I__5614 (
            .O(N__31310),
            .I(\ADC_VDC.genclk.n19470 ));
    InMux I__5613 (
            .O(N__31307),
            .I(\ADC_VDC.genclk.n19471 ));
    InMux I__5612 (
            .O(N__31304),
            .I(\ADC_VDC.genclk.n19472 ));
    InMux I__5611 (
            .O(N__31301),
            .I(N__31296));
    InMux I__5610 (
            .O(N__31300),
            .I(N__31291));
    InMux I__5609 (
            .O(N__31299),
            .I(N__31291));
    LocalMux I__5608 (
            .O(N__31296),
            .I(buf_dds0_6));
    LocalMux I__5607 (
            .O(N__31291),
            .I(buf_dds0_6));
    CascadeMux I__5606 (
            .O(N__31286),
            .I(N__31283));
    InMux I__5605 (
            .O(N__31283),
            .I(N__31280));
    LocalMux I__5604 (
            .O(N__31280),
            .I(N__31277));
    Span4Mux_h I__5603 (
            .O(N__31277),
            .I(N__31272));
    InMux I__5602 (
            .O(N__31276),
            .I(N__31267));
    InMux I__5601 (
            .O(N__31275),
            .I(N__31267));
    Odrv4 I__5600 (
            .O(N__31272),
            .I(buf_dds1_6));
    LocalMux I__5599 (
            .O(N__31267),
            .I(buf_dds1_6));
    CEMux I__5598 (
            .O(N__31262),
            .I(N__31259));
    LocalMux I__5597 (
            .O(N__31259),
            .I(N__31256));
    Span4Mux_h I__5596 (
            .O(N__31256),
            .I(N__31253));
    Odrv4 I__5595 (
            .O(N__31253),
            .I(n11757));
    CascadeMux I__5594 (
            .O(N__31250),
            .I(N__31246));
    InMux I__5593 (
            .O(N__31249),
            .I(N__31241));
    InMux I__5592 (
            .O(N__31246),
            .I(N__31234));
    InMux I__5591 (
            .O(N__31245),
            .I(N__31234));
    InMux I__5590 (
            .O(N__31244),
            .I(N__31234));
    LocalMux I__5589 (
            .O(N__31241),
            .I(wdtick_cnt_0));
    LocalMux I__5588 (
            .O(N__31234),
            .I(wdtick_cnt_0));
    InMux I__5587 (
            .O(N__31229),
            .I(N__31223));
    InMux I__5586 (
            .O(N__31228),
            .I(N__31216));
    InMux I__5585 (
            .O(N__31227),
            .I(N__31216));
    InMux I__5584 (
            .O(N__31226),
            .I(N__31216));
    LocalMux I__5583 (
            .O(N__31223),
            .I(wdtick_cnt_1));
    LocalMux I__5582 (
            .O(N__31216),
            .I(wdtick_cnt_1));
    CascadeMux I__5581 (
            .O(N__31211),
            .I(N__31208));
    InMux I__5580 (
            .O(N__31208),
            .I(N__31203));
    InMux I__5579 (
            .O(N__31207),
            .I(N__31198));
    InMux I__5578 (
            .O(N__31206),
            .I(N__31198));
    LocalMux I__5577 (
            .O(N__31203),
            .I(wdtick_cnt_2));
    LocalMux I__5576 (
            .O(N__31198),
            .I(wdtick_cnt_2));
    InMux I__5575 (
            .O(N__31193),
            .I(N__31190));
    LocalMux I__5574 (
            .O(N__31190),
            .I(N__31185));
    InMux I__5573 (
            .O(N__31189),
            .I(N__31182));
    InMux I__5572 (
            .O(N__31188),
            .I(N__31179));
    Span12Mux_h I__5571 (
            .O(N__31185),
            .I(N__31174));
    LocalMux I__5570 (
            .O(N__31182),
            .I(N__31174));
    LocalMux I__5569 (
            .O(N__31179),
            .I(buf_dds0_0));
    Odrv12 I__5568 (
            .O(N__31174),
            .I(buf_dds0_0));
    CascadeMux I__5567 (
            .O(N__31169),
            .I(n17411_cascade_));
    CascadeMux I__5566 (
            .O(N__31166),
            .I(N__31163));
    CascadeBuf I__5565 (
            .O(N__31163),
            .I(N__31160));
    CascadeMux I__5564 (
            .O(N__31160),
            .I(N__31157));
    CascadeBuf I__5563 (
            .O(N__31157),
            .I(N__31154));
    CascadeMux I__5562 (
            .O(N__31154),
            .I(N__31151));
    CascadeBuf I__5561 (
            .O(N__31151),
            .I(N__31148));
    CascadeMux I__5560 (
            .O(N__31148),
            .I(N__31145));
    CascadeBuf I__5559 (
            .O(N__31145),
            .I(N__31142));
    CascadeMux I__5558 (
            .O(N__31142),
            .I(N__31139));
    CascadeBuf I__5557 (
            .O(N__31139),
            .I(N__31136));
    CascadeMux I__5556 (
            .O(N__31136),
            .I(N__31133));
    CascadeBuf I__5555 (
            .O(N__31133),
            .I(N__31130));
    CascadeMux I__5554 (
            .O(N__31130),
            .I(N__31127));
    CascadeBuf I__5553 (
            .O(N__31127),
            .I(N__31124));
    CascadeMux I__5552 (
            .O(N__31124),
            .I(N__31121));
    CascadeBuf I__5551 (
            .O(N__31121),
            .I(N__31118));
    CascadeMux I__5550 (
            .O(N__31118),
            .I(N__31114));
    CascadeMux I__5549 (
            .O(N__31117),
            .I(N__31111));
    CascadeBuf I__5548 (
            .O(N__31114),
            .I(N__31108));
    CascadeBuf I__5547 (
            .O(N__31111),
            .I(N__31105));
    CascadeMux I__5546 (
            .O(N__31108),
            .I(N__31102));
    CascadeMux I__5545 (
            .O(N__31105),
            .I(N__31099));
    InMux I__5544 (
            .O(N__31102),
            .I(N__31096));
    InMux I__5543 (
            .O(N__31099),
            .I(N__31093));
    LocalMux I__5542 (
            .O(N__31096),
            .I(N__31090));
    LocalMux I__5541 (
            .O(N__31093),
            .I(N__31087));
    Span4Mux_h I__5540 (
            .O(N__31090),
            .I(N__31084));
    Span12Mux_s9_h I__5539 (
            .O(N__31087),
            .I(N__31081));
    Span4Mux_h I__5538 (
            .O(N__31084),
            .I(N__31078));
    Span12Mux_v I__5537 (
            .O(N__31081),
            .I(N__31075));
    Span4Mux_v I__5536 (
            .O(N__31078),
            .I(N__31072));
    Odrv12 I__5535 (
            .O(N__31075),
            .I(data_index_9_N_216_5));
    Odrv4 I__5534 (
            .O(N__31072),
            .I(data_index_9_N_216_5));
    InMux I__5533 (
            .O(N__31067),
            .I(N__31061));
    InMux I__5532 (
            .O(N__31066),
            .I(N__31061));
    LocalMux I__5531 (
            .O(N__31061),
            .I(n17409));
    InMux I__5530 (
            .O(N__31058),
            .I(N__31055));
    LocalMux I__5529 (
            .O(N__31055),
            .I(n17411));
    InMux I__5528 (
            .O(N__31052),
            .I(N__31047));
    InMux I__5527 (
            .O(N__31051),
            .I(N__31044));
    InMux I__5526 (
            .O(N__31050),
            .I(N__31041));
    LocalMux I__5525 (
            .O(N__31047),
            .I(data_index_5));
    LocalMux I__5524 (
            .O(N__31044),
            .I(data_index_5));
    LocalMux I__5523 (
            .O(N__31041),
            .I(data_index_5));
    CascadeMux I__5522 (
            .O(N__31034),
            .I(n8828_cascade_));
    InMux I__5521 (
            .O(N__31031),
            .I(N__31026));
    InMux I__5520 (
            .O(N__31030),
            .I(N__31023));
    InMux I__5519 (
            .O(N__31029),
            .I(N__31020));
    LocalMux I__5518 (
            .O(N__31026),
            .I(data_index_0));
    LocalMux I__5517 (
            .O(N__31023),
            .I(data_index_0));
    LocalMux I__5516 (
            .O(N__31020),
            .I(data_index_0));
    InMux I__5515 (
            .O(N__31013),
            .I(N__31010));
    LocalMux I__5514 (
            .O(N__31010),
            .I(N__31006));
    InMux I__5513 (
            .O(N__31009),
            .I(N__31003));
    Span4Mux_h I__5512 (
            .O(N__31006),
            .I(N__31000));
    LocalMux I__5511 (
            .O(N__31003),
            .I(n8_adj_1532));
    Odrv4 I__5510 (
            .O(N__31000),
            .I(n8_adj_1532));
    InMux I__5509 (
            .O(N__30995),
            .I(N__30990));
    InMux I__5508 (
            .O(N__30994),
            .I(N__30987));
    InMux I__5507 (
            .O(N__30993),
            .I(N__30984));
    LocalMux I__5506 (
            .O(N__30990),
            .I(N__30979));
    LocalMux I__5505 (
            .O(N__30987),
            .I(N__30979));
    LocalMux I__5504 (
            .O(N__30984),
            .I(N__30974));
    Span4Mux_v I__5503 (
            .O(N__30979),
            .I(N__30974));
    Odrv4 I__5502 (
            .O(N__30974),
            .I(buf_dds1_13));
    CascadeMux I__5501 (
            .O(N__30971),
            .I(N__30968));
    InMux I__5500 (
            .O(N__30968),
            .I(N__30959));
    InMux I__5499 (
            .O(N__30967),
            .I(N__30959));
    InMux I__5498 (
            .O(N__30966),
            .I(N__30959));
    LocalMux I__5497 (
            .O(N__30959),
            .I(cmd_rdadctmp_18));
    IoInMux I__5496 (
            .O(N__30956),
            .I(N__30953));
    LocalMux I__5495 (
            .O(N__30953),
            .I(N__30950));
    Span4Mux_s3_h I__5494 (
            .O(N__30950),
            .I(N__30947));
    Sp12to4 I__5493 (
            .O(N__30947),
            .I(N__30943));
    InMux I__5492 (
            .O(N__30946),
            .I(N__30939));
    Span12Mux_v I__5491 (
            .O(N__30943),
            .I(N__30936));
    InMux I__5490 (
            .O(N__30942),
            .I(N__30933));
    LocalMux I__5489 (
            .O(N__30939),
            .I(N__30930));
    Odrv12 I__5488 (
            .O(N__30936),
            .I(AMPV_POW));
    LocalMux I__5487 (
            .O(N__30933),
            .I(AMPV_POW));
    Odrv4 I__5486 (
            .O(N__30930),
            .I(AMPV_POW));
    CascadeMux I__5485 (
            .O(N__30923),
            .I(N__30920));
    InMux I__5484 (
            .O(N__30920),
            .I(N__30917));
    LocalMux I__5483 (
            .O(N__30917),
            .I(N__30914));
    Odrv12 I__5482 (
            .O(N__30914),
            .I(n23_adj_1536));
    InMux I__5481 (
            .O(N__30911),
            .I(N__30904));
    InMux I__5480 (
            .O(N__30910),
            .I(N__30904));
    InMux I__5479 (
            .O(N__30909),
            .I(N__30901));
    LocalMux I__5478 (
            .O(N__30904),
            .I(cmd_rdadctmp_21_adj_1429));
    LocalMux I__5477 (
            .O(N__30901),
            .I(cmd_rdadctmp_21_adj_1429));
    InMux I__5476 (
            .O(N__30896),
            .I(N__30892));
    InMux I__5475 (
            .O(N__30895),
            .I(N__30889));
    LocalMux I__5474 (
            .O(N__30892),
            .I(N__30886));
    LocalMux I__5473 (
            .O(N__30889),
            .I(n7_adj_1531));
    Odrv4 I__5472 (
            .O(N__30886),
            .I(n7_adj_1531));
    CascadeMux I__5471 (
            .O(N__30881),
            .I(N__30878));
    InMux I__5470 (
            .O(N__30878),
            .I(N__30873));
    CascadeMux I__5469 (
            .O(N__30877),
            .I(N__30870));
    CascadeMux I__5468 (
            .O(N__30876),
            .I(N__30867));
    LocalMux I__5467 (
            .O(N__30873),
            .I(N__30864));
    InMux I__5466 (
            .O(N__30870),
            .I(N__30859));
    InMux I__5465 (
            .O(N__30867),
            .I(N__30859));
    Odrv12 I__5464 (
            .O(N__30864),
            .I(cmd_rdadctmp_22_adj_1428));
    LocalMux I__5463 (
            .O(N__30859),
            .I(cmd_rdadctmp_22_adj_1428));
    InMux I__5462 (
            .O(N__30854),
            .I(N__30851));
    LocalMux I__5461 (
            .O(N__30851),
            .I(N__30847));
    CascadeMux I__5460 (
            .O(N__30850),
            .I(N__30844));
    Span4Mux_v I__5459 (
            .O(N__30847),
            .I(N__30841));
    InMux I__5458 (
            .O(N__30844),
            .I(N__30838));
    Odrv4 I__5457 (
            .O(N__30841),
            .I(buf_adcdata_vdc_9));
    LocalMux I__5456 (
            .O(N__30838),
            .I(buf_adcdata_vdc_9));
    InMux I__5455 (
            .O(N__30833),
            .I(N__30830));
    LocalMux I__5454 (
            .O(N__30830),
            .I(N__30827));
    Span4Mux_v I__5453 (
            .O(N__30827),
            .I(N__30824));
    Span4Mux_h I__5452 (
            .O(N__30824),
            .I(N__30820));
    InMux I__5451 (
            .O(N__30823),
            .I(N__30817));
    Span4Mux_h I__5450 (
            .O(N__30820),
            .I(N__30814));
    LocalMux I__5449 (
            .O(N__30817),
            .I(N__30808));
    Span4Mux_v I__5448 (
            .O(N__30814),
            .I(N__30808));
    InMux I__5447 (
            .O(N__30813),
            .I(N__30805));
    Odrv4 I__5446 (
            .O(N__30808),
            .I(buf_adcdata_vac_9));
    LocalMux I__5445 (
            .O(N__30805),
            .I(buf_adcdata_vac_9));
    CascadeMux I__5444 (
            .O(N__30800),
            .I(N__30797));
    CascadeBuf I__5443 (
            .O(N__30797),
            .I(N__30794));
    CascadeMux I__5442 (
            .O(N__30794),
            .I(N__30791));
    CascadeBuf I__5441 (
            .O(N__30791),
            .I(N__30788));
    CascadeMux I__5440 (
            .O(N__30788),
            .I(N__30785));
    CascadeBuf I__5439 (
            .O(N__30785),
            .I(N__30782));
    CascadeMux I__5438 (
            .O(N__30782),
            .I(N__30779));
    CascadeBuf I__5437 (
            .O(N__30779),
            .I(N__30776));
    CascadeMux I__5436 (
            .O(N__30776),
            .I(N__30773));
    CascadeBuf I__5435 (
            .O(N__30773),
            .I(N__30770));
    CascadeMux I__5434 (
            .O(N__30770),
            .I(N__30767));
    CascadeBuf I__5433 (
            .O(N__30767),
            .I(N__30764));
    CascadeMux I__5432 (
            .O(N__30764),
            .I(N__30761));
    CascadeBuf I__5431 (
            .O(N__30761),
            .I(N__30757));
    CascadeMux I__5430 (
            .O(N__30760),
            .I(N__30754));
    CascadeMux I__5429 (
            .O(N__30757),
            .I(N__30751));
    CascadeBuf I__5428 (
            .O(N__30754),
            .I(N__30748));
    CascadeBuf I__5427 (
            .O(N__30751),
            .I(N__30745));
    CascadeMux I__5426 (
            .O(N__30748),
            .I(N__30742));
    CascadeMux I__5425 (
            .O(N__30745),
            .I(N__30739));
    InMux I__5424 (
            .O(N__30742),
            .I(N__30736));
    CascadeBuf I__5423 (
            .O(N__30739),
            .I(N__30733));
    LocalMux I__5422 (
            .O(N__30736),
            .I(N__30730));
    CascadeMux I__5421 (
            .O(N__30733),
            .I(N__30727));
    Span4Mux_h I__5420 (
            .O(N__30730),
            .I(N__30724));
    InMux I__5419 (
            .O(N__30727),
            .I(N__30721));
    Span4Mux_v I__5418 (
            .O(N__30724),
            .I(N__30717));
    LocalMux I__5417 (
            .O(N__30721),
            .I(N__30714));
    InMux I__5416 (
            .O(N__30720),
            .I(N__30711));
    Span4Mux_h I__5415 (
            .O(N__30717),
            .I(N__30708));
    Span12Mux_h I__5414 (
            .O(N__30714),
            .I(N__30705));
    LocalMux I__5413 (
            .O(N__30711),
            .I(data_count_8));
    Odrv4 I__5412 (
            .O(N__30708),
            .I(data_count_8));
    Odrv12 I__5411 (
            .O(N__30705),
            .I(data_count_8));
    InMux I__5410 (
            .O(N__30698),
            .I(bfn_11_12_0_));
    InMux I__5409 (
            .O(N__30695),
            .I(n19353));
    CascadeMux I__5408 (
            .O(N__30692),
            .I(N__30689));
    CascadeBuf I__5407 (
            .O(N__30689),
            .I(N__30686));
    CascadeMux I__5406 (
            .O(N__30686),
            .I(N__30683));
    CascadeBuf I__5405 (
            .O(N__30683),
            .I(N__30680));
    CascadeMux I__5404 (
            .O(N__30680),
            .I(N__30677));
    CascadeBuf I__5403 (
            .O(N__30677),
            .I(N__30674));
    CascadeMux I__5402 (
            .O(N__30674),
            .I(N__30671));
    CascadeBuf I__5401 (
            .O(N__30671),
            .I(N__30668));
    CascadeMux I__5400 (
            .O(N__30668),
            .I(N__30665));
    CascadeBuf I__5399 (
            .O(N__30665),
            .I(N__30662));
    CascadeMux I__5398 (
            .O(N__30662),
            .I(N__30659));
    CascadeBuf I__5397 (
            .O(N__30659),
            .I(N__30656));
    CascadeMux I__5396 (
            .O(N__30656),
            .I(N__30653));
    CascadeBuf I__5395 (
            .O(N__30653),
            .I(N__30650));
    CascadeMux I__5394 (
            .O(N__30650),
            .I(N__30647));
    CascadeBuf I__5393 (
            .O(N__30647),
            .I(N__30643));
    CascadeMux I__5392 (
            .O(N__30646),
            .I(N__30640));
    CascadeMux I__5391 (
            .O(N__30643),
            .I(N__30637));
    CascadeBuf I__5390 (
            .O(N__30640),
            .I(N__30634));
    CascadeBuf I__5389 (
            .O(N__30637),
            .I(N__30631));
    CascadeMux I__5388 (
            .O(N__30634),
            .I(N__30628));
    CascadeMux I__5387 (
            .O(N__30631),
            .I(N__30625));
    InMux I__5386 (
            .O(N__30628),
            .I(N__30622));
    InMux I__5385 (
            .O(N__30625),
            .I(N__30619));
    LocalMux I__5384 (
            .O(N__30622),
            .I(N__30616));
    LocalMux I__5383 (
            .O(N__30619),
            .I(N__30613));
    Span4Mux_h I__5382 (
            .O(N__30616),
            .I(N__30610));
    Span4Mux_v I__5381 (
            .O(N__30613),
            .I(N__30607));
    Span4Mux_h I__5380 (
            .O(N__30610),
            .I(N__30603));
    Sp12to4 I__5379 (
            .O(N__30607),
            .I(N__30600));
    InMux I__5378 (
            .O(N__30606),
            .I(N__30597));
    Sp12to4 I__5377 (
            .O(N__30603),
            .I(N__30594));
    Span12Mux_h I__5376 (
            .O(N__30600),
            .I(N__30591));
    LocalMux I__5375 (
            .O(N__30597),
            .I(data_count_9));
    Odrv12 I__5374 (
            .O(N__30594),
            .I(data_count_9));
    Odrv12 I__5373 (
            .O(N__30591),
            .I(data_count_9));
    InMux I__5372 (
            .O(N__30584),
            .I(N__30581));
    LocalMux I__5371 (
            .O(N__30581),
            .I(N__30577));
    InMux I__5370 (
            .O(N__30580),
            .I(N__30573));
    Span4Mux_v I__5369 (
            .O(N__30577),
            .I(N__30570));
    CascadeMux I__5368 (
            .O(N__30576),
            .I(N__30567));
    LocalMux I__5367 (
            .O(N__30573),
            .I(N__30564));
    Span4Mux_h I__5366 (
            .O(N__30570),
            .I(N__30561));
    InMux I__5365 (
            .O(N__30567),
            .I(N__30558));
    Span4Mux_h I__5364 (
            .O(N__30564),
            .I(N__30555));
    Span4Mux_v I__5363 (
            .O(N__30561),
            .I(N__30552));
    LocalMux I__5362 (
            .O(N__30558),
            .I(cmd_rdadctmp_16));
    Odrv4 I__5361 (
            .O(N__30555),
            .I(cmd_rdadctmp_16));
    Odrv4 I__5360 (
            .O(N__30552),
            .I(cmd_rdadctmp_16));
    InMux I__5359 (
            .O(N__30545),
            .I(N__30542));
    LocalMux I__5358 (
            .O(N__30542),
            .I(N__30539));
    Span4Mux_v I__5357 (
            .O(N__30539),
            .I(N__30536));
    Span4Mux_h I__5356 (
            .O(N__30536),
            .I(N__30532));
    InMux I__5355 (
            .O(N__30535),
            .I(N__30529));
    Odrv4 I__5354 (
            .O(N__30532),
            .I(buf_adcdata_vdc_8));
    LocalMux I__5353 (
            .O(N__30529),
            .I(buf_adcdata_vdc_8));
    InMux I__5352 (
            .O(N__30524),
            .I(N__30521));
    LocalMux I__5351 (
            .O(N__30521),
            .I(N__30518));
    Span4Mux_v I__5350 (
            .O(N__30518),
            .I(N__30515));
    Sp12to4 I__5349 (
            .O(N__30515),
            .I(N__30512));
    Span12Mux_h I__5348 (
            .O(N__30512),
            .I(N__30507));
    InMux I__5347 (
            .O(N__30511),
            .I(N__30502));
    InMux I__5346 (
            .O(N__30510),
            .I(N__30502));
    Odrv12 I__5345 (
            .O(N__30507),
            .I(buf_adcdata_vac_8));
    LocalMux I__5344 (
            .O(N__30502),
            .I(buf_adcdata_vac_8));
    InMux I__5343 (
            .O(N__30497),
            .I(N__30494));
    LocalMux I__5342 (
            .O(N__30494),
            .I(N__30491));
    Span4Mux_v I__5341 (
            .O(N__30491),
            .I(N__30488));
    Span4Mux_v I__5340 (
            .O(N__30488),
            .I(N__30485));
    Span4Mux_h I__5339 (
            .O(N__30485),
            .I(N__30481));
    InMux I__5338 (
            .O(N__30484),
            .I(N__30478));
    Odrv4 I__5337 (
            .O(N__30481),
            .I(buf_adcdata_vdc_10));
    LocalMux I__5336 (
            .O(N__30478),
            .I(buf_adcdata_vdc_10));
    InMux I__5335 (
            .O(N__30473),
            .I(N__30470));
    LocalMux I__5334 (
            .O(N__30470),
            .I(N__30467));
    Span4Mux_v I__5333 (
            .O(N__30467),
            .I(N__30464));
    Span4Mux_v I__5332 (
            .O(N__30464),
            .I(N__30461));
    Sp12to4 I__5331 (
            .O(N__30461),
            .I(N__30456));
    InMux I__5330 (
            .O(N__30460),
            .I(N__30451));
    InMux I__5329 (
            .O(N__30459),
            .I(N__30451));
    Odrv12 I__5328 (
            .O(N__30456),
            .I(buf_adcdata_vac_10));
    LocalMux I__5327 (
            .O(N__30451),
            .I(buf_adcdata_vac_10));
    CascadeMux I__5326 (
            .O(N__30446),
            .I(N__30442));
    CascadeMux I__5325 (
            .O(N__30445),
            .I(N__30439));
    InMux I__5324 (
            .O(N__30442),
            .I(N__30434));
    InMux I__5323 (
            .O(N__30439),
            .I(N__30434));
    LocalMux I__5322 (
            .O(N__30434),
            .I(N__30431));
    Span4Mux_v I__5321 (
            .O(N__30431),
            .I(N__30427));
    CascadeMux I__5320 (
            .O(N__30430),
            .I(N__30424));
    Span4Mux_v I__5319 (
            .O(N__30427),
            .I(N__30421));
    InMux I__5318 (
            .O(N__30424),
            .I(N__30418));
    Odrv4 I__5317 (
            .O(N__30421),
            .I(cmd_rdadctmp_17));
    LocalMux I__5316 (
            .O(N__30418),
            .I(cmd_rdadctmp_17));
    CascadeMux I__5315 (
            .O(N__30413),
            .I(n20590_cascade_));
    InMux I__5314 (
            .O(N__30410),
            .I(N__30407));
    LocalMux I__5313 (
            .O(N__30407),
            .I(N__30404));
    Span4Mux_v I__5312 (
            .O(N__30404),
            .I(N__30401));
    Span4Mux_h I__5311 (
            .O(N__30401),
            .I(N__30398));
    Span4Mux_h I__5310 (
            .O(N__30398),
            .I(N__30393));
    InMux I__5309 (
            .O(N__30397),
            .I(N__30388));
    InMux I__5308 (
            .O(N__30396),
            .I(N__30388));
    Odrv4 I__5307 (
            .O(N__30393),
            .I(buf_adcdata_vac_16));
    LocalMux I__5306 (
            .O(N__30388),
            .I(buf_adcdata_vac_16));
    CascadeMux I__5305 (
            .O(N__30383),
            .I(N__30380));
    CascadeBuf I__5304 (
            .O(N__30380),
            .I(N__30377));
    CascadeMux I__5303 (
            .O(N__30377),
            .I(N__30374));
    CascadeBuf I__5302 (
            .O(N__30374),
            .I(N__30371));
    CascadeMux I__5301 (
            .O(N__30371),
            .I(N__30368));
    CascadeBuf I__5300 (
            .O(N__30368),
            .I(N__30365));
    CascadeMux I__5299 (
            .O(N__30365),
            .I(N__30362));
    CascadeBuf I__5298 (
            .O(N__30362),
            .I(N__30359));
    CascadeMux I__5297 (
            .O(N__30359),
            .I(N__30356));
    CascadeBuf I__5296 (
            .O(N__30356),
            .I(N__30353));
    CascadeMux I__5295 (
            .O(N__30353),
            .I(N__30350));
    CascadeBuf I__5294 (
            .O(N__30350),
            .I(N__30347));
    CascadeMux I__5293 (
            .O(N__30347),
            .I(N__30344));
    CascadeBuf I__5292 (
            .O(N__30344),
            .I(N__30341));
    CascadeMux I__5291 (
            .O(N__30341),
            .I(N__30338));
    CascadeBuf I__5290 (
            .O(N__30338),
            .I(N__30334));
    CascadeMux I__5289 (
            .O(N__30337),
            .I(N__30331));
    CascadeMux I__5288 (
            .O(N__30334),
            .I(N__30328));
    CascadeBuf I__5287 (
            .O(N__30331),
            .I(N__30325));
    CascadeBuf I__5286 (
            .O(N__30328),
            .I(N__30322));
    CascadeMux I__5285 (
            .O(N__30325),
            .I(N__30319));
    CascadeMux I__5284 (
            .O(N__30322),
            .I(N__30316));
    InMux I__5283 (
            .O(N__30319),
            .I(N__30313));
    InMux I__5282 (
            .O(N__30316),
            .I(N__30310));
    LocalMux I__5281 (
            .O(N__30313),
            .I(N__30307));
    LocalMux I__5280 (
            .O(N__30310),
            .I(N__30304));
    Span4Mux_v I__5279 (
            .O(N__30307),
            .I(N__30300));
    Span4Mux_v I__5278 (
            .O(N__30304),
            .I(N__30297));
    CascadeMux I__5277 (
            .O(N__30303),
            .I(N__30294));
    Sp12to4 I__5276 (
            .O(N__30300),
            .I(N__30291));
    Sp12to4 I__5275 (
            .O(N__30297),
            .I(N__30288));
    InMux I__5274 (
            .O(N__30294),
            .I(N__30285));
    Span12Mux_h I__5273 (
            .O(N__30291),
            .I(N__30280));
    Span12Mux_h I__5272 (
            .O(N__30288),
            .I(N__30280));
    LocalMux I__5271 (
            .O(N__30285),
            .I(data_count_0));
    Odrv12 I__5270 (
            .O(N__30280),
            .I(data_count_0));
    CascadeMux I__5269 (
            .O(N__30275),
            .I(N__30272));
    CascadeBuf I__5268 (
            .O(N__30272),
            .I(N__30269));
    CascadeMux I__5267 (
            .O(N__30269),
            .I(N__30266));
    CascadeBuf I__5266 (
            .O(N__30266),
            .I(N__30263));
    CascadeMux I__5265 (
            .O(N__30263),
            .I(N__30260));
    CascadeBuf I__5264 (
            .O(N__30260),
            .I(N__30257));
    CascadeMux I__5263 (
            .O(N__30257),
            .I(N__30254));
    CascadeBuf I__5262 (
            .O(N__30254),
            .I(N__30251));
    CascadeMux I__5261 (
            .O(N__30251),
            .I(N__30248));
    CascadeBuf I__5260 (
            .O(N__30248),
            .I(N__30245));
    CascadeMux I__5259 (
            .O(N__30245),
            .I(N__30242));
    CascadeBuf I__5258 (
            .O(N__30242),
            .I(N__30239));
    CascadeMux I__5257 (
            .O(N__30239),
            .I(N__30236));
    CascadeBuf I__5256 (
            .O(N__30236),
            .I(N__30233));
    CascadeMux I__5255 (
            .O(N__30233),
            .I(N__30230));
    CascadeBuf I__5254 (
            .O(N__30230),
            .I(N__30226));
    CascadeMux I__5253 (
            .O(N__30229),
            .I(N__30223));
    CascadeMux I__5252 (
            .O(N__30226),
            .I(N__30220));
    CascadeBuf I__5251 (
            .O(N__30223),
            .I(N__30217));
    CascadeBuf I__5250 (
            .O(N__30220),
            .I(N__30214));
    CascadeMux I__5249 (
            .O(N__30217),
            .I(N__30211));
    CascadeMux I__5248 (
            .O(N__30214),
            .I(N__30208));
    InMux I__5247 (
            .O(N__30211),
            .I(N__30205));
    InMux I__5246 (
            .O(N__30208),
            .I(N__30202));
    LocalMux I__5245 (
            .O(N__30205),
            .I(N__30199));
    LocalMux I__5244 (
            .O(N__30202),
            .I(N__30196));
    Span4Mux_h I__5243 (
            .O(N__30199),
            .I(N__30193));
    Span4Mux_h I__5242 (
            .O(N__30196),
            .I(N__30190));
    Sp12to4 I__5241 (
            .O(N__30193),
            .I(N__30186));
    Sp12to4 I__5240 (
            .O(N__30190),
            .I(N__30183));
    InMux I__5239 (
            .O(N__30189),
            .I(N__30180));
    Span12Mux_v I__5238 (
            .O(N__30186),
            .I(N__30175));
    Span12Mux_v I__5237 (
            .O(N__30183),
            .I(N__30175));
    LocalMux I__5236 (
            .O(N__30180),
            .I(data_count_1));
    Odrv12 I__5235 (
            .O(N__30175),
            .I(data_count_1));
    InMux I__5234 (
            .O(N__30170),
            .I(n19345));
    CascadeMux I__5233 (
            .O(N__30167),
            .I(N__30164));
    CascadeBuf I__5232 (
            .O(N__30164),
            .I(N__30161));
    CascadeMux I__5231 (
            .O(N__30161),
            .I(N__30158));
    CascadeBuf I__5230 (
            .O(N__30158),
            .I(N__30155));
    CascadeMux I__5229 (
            .O(N__30155),
            .I(N__30152));
    CascadeBuf I__5228 (
            .O(N__30152),
            .I(N__30149));
    CascadeMux I__5227 (
            .O(N__30149),
            .I(N__30146));
    CascadeBuf I__5226 (
            .O(N__30146),
            .I(N__30143));
    CascadeMux I__5225 (
            .O(N__30143),
            .I(N__30140));
    CascadeBuf I__5224 (
            .O(N__30140),
            .I(N__30137));
    CascadeMux I__5223 (
            .O(N__30137),
            .I(N__30134));
    CascadeBuf I__5222 (
            .O(N__30134),
            .I(N__30131));
    CascadeMux I__5221 (
            .O(N__30131),
            .I(N__30128));
    CascadeBuf I__5220 (
            .O(N__30128),
            .I(N__30125));
    CascadeMux I__5219 (
            .O(N__30125),
            .I(N__30122));
    CascadeBuf I__5218 (
            .O(N__30122),
            .I(N__30119));
    CascadeMux I__5217 (
            .O(N__30119),
            .I(N__30116));
    CascadeBuf I__5216 (
            .O(N__30116),
            .I(N__30112));
    CascadeMux I__5215 (
            .O(N__30115),
            .I(N__30109));
    CascadeMux I__5214 (
            .O(N__30112),
            .I(N__30106));
    CascadeBuf I__5213 (
            .O(N__30109),
            .I(N__30103));
    InMux I__5212 (
            .O(N__30106),
            .I(N__30100));
    CascadeMux I__5211 (
            .O(N__30103),
            .I(N__30097));
    LocalMux I__5210 (
            .O(N__30100),
            .I(N__30094));
    InMux I__5209 (
            .O(N__30097),
            .I(N__30091));
    Span4Mux_v I__5208 (
            .O(N__30094),
            .I(N__30088));
    LocalMux I__5207 (
            .O(N__30091),
            .I(N__30085));
    Span4Mux_v I__5206 (
            .O(N__30088),
            .I(N__30082));
    Span4Mux_v I__5205 (
            .O(N__30085),
            .I(N__30079));
    Sp12to4 I__5204 (
            .O(N__30082),
            .I(N__30076));
    Sp12to4 I__5203 (
            .O(N__30079),
            .I(N__30072));
    Span12Mux_h I__5202 (
            .O(N__30076),
            .I(N__30069));
    InMux I__5201 (
            .O(N__30075),
            .I(N__30066));
    Span12Mux_h I__5200 (
            .O(N__30072),
            .I(N__30061));
    Span12Mux_v I__5199 (
            .O(N__30069),
            .I(N__30061));
    LocalMux I__5198 (
            .O(N__30066),
            .I(data_count_2));
    Odrv12 I__5197 (
            .O(N__30061),
            .I(data_count_2));
    InMux I__5196 (
            .O(N__30056),
            .I(n19346));
    CascadeMux I__5195 (
            .O(N__30053),
            .I(N__30050));
    CascadeBuf I__5194 (
            .O(N__30050),
            .I(N__30047));
    CascadeMux I__5193 (
            .O(N__30047),
            .I(N__30044));
    CascadeBuf I__5192 (
            .O(N__30044),
            .I(N__30041));
    CascadeMux I__5191 (
            .O(N__30041),
            .I(N__30038));
    CascadeBuf I__5190 (
            .O(N__30038),
            .I(N__30035));
    CascadeMux I__5189 (
            .O(N__30035),
            .I(N__30032));
    CascadeBuf I__5188 (
            .O(N__30032),
            .I(N__30029));
    CascadeMux I__5187 (
            .O(N__30029),
            .I(N__30026));
    CascadeBuf I__5186 (
            .O(N__30026),
            .I(N__30023));
    CascadeMux I__5185 (
            .O(N__30023),
            .I(N__30020));
    CascadeBuf I__5184 (
            .O(N__30020),
            .I(N__30017));
    CascadeMux I__5183 (
            .O(N__30017),
            .I(N__30014));
    CascadeBuf I__5182 (
            .O(N__30014),
            .I(N__30011));
    CascadeMux I__5181 (
            .O(N__30011),
            .I(N__30008));
    CascadeBuf I__5180 (
            .O(N__30008),
            .I(N__30005));
    CascadeMux I__5179 (
            .O(N__30005),
            .I(N__30002));
    CascadeBuf I__5178 (
            .O(N__30002),
            .I(N__29998));
    CascadeMux I__5177 (
            .O(N__30001),
            .I(N__29995));
    CascadeMux I__5176 (
            .O(N__29998),
            .I(N__29992));
    CascadeBuf I__5175 (
            .O(N__29995),
            .I(N__29989));
    InMux I__5174 (
            .O(N__29992),
            .I(N__29986));
    CascadeMux I__5173 (
            .O(N__29989),
            .I(N__29983));
    LocalMux I__5172 (
            .O(N__29986),
            .I(N__29980));
    InMux I__5171 (
            .O(N__29983),
            .I(N__29977));
    Span4Mux_v I__5170 (
            .O(N__29980),
            .I(N__29974));
    LocalMux I__5169 (
            .O(N__29977),
            .I(N__29970));
    Sp12to4 I__5168 (
            .O(N__29974),
            .I(N__29967));
    InMux I__5167 (
            .O(N__29973),
            .I(N__29964));
    Span12Mux_v I__5166 (
            .O(N__29970),
            .I(N__29961));
    Span12Mux_h I__5165 (
            .O(N__29967),
            .I(N__29958));
    LocalMux I__5164 (
            .O(N__29964),
            .I(data_count_3));
    Odrv12 I__5163 (
            .O(N__29961),
            .I(data_count_3));
    Odrv12 I__5162 (
            .O(N__29958),
            .I(data_count_3));
    InMux I__5161 (
            .O(N__29951),
            .I(n19347));
    CascadeMux I__5160 (
            .O(N__29948),
            .I(N__29945));
    CascadeBuf I__5159 (
            .O(N__29945),
            .I(N__29942));
    CascadeMux I__5158 (
            .O(N__29942),
            .I(N__29939));
    CascadeBuf I__5157 (
            .O(N__29939),
            .I(N__29936));
    CascadeMux I__5156 (
            .O(N__29936),
            .I(N__29933));
    CascadeBuf I__5155 (
            .O(N__29933),
            .I(N__29930));
    CascadeMux I__5154 (
            .O(N__29930),
            .I(N__29927));
    CascadeBuf I__5153 (
            .O(N__29927),
            .I(N__29924));
    CascadeMux I__5152 (
            .O(N__29924),
            .I(N__29921));
    CascadeBuf I__5151 (
            .O(N__29921),
            .I(N__29918));
    CascadeMux I__5150 (
            .O(N__29918),
            .I(N__29915));
    CascadeBuf I__5149 (
            .O(N__29915),
            .I(N__29912));
    CascadeMux I__5148 (
            .O(N__29912),
            .I(N__29909));
    CascadeBuf I__5147 (
            .O(N__29909),
            .I(N__29906));
    CascadeMux I__5146 (
            .O(N__29906),
            .I(N__29903));
    CascadeBuf I__5145 (
            .O(N__29903),
            .I(N__29900));
    CascadeMux I__5144 (
            .O(N__29900),
            .I(N__29896));
    CascadeMux I__5143 (
            .O(N__29899),
            .I(N__29893));
    CascadeBuf I__5142 (
            .O(N__29896),
            .I(N__29890));
    CascadeBuf I__5141 (
            .O(N__29893),
            .I(N__29887));
    CascadeMux I__5140 (
            .O(N__29890),
            .I(N__29884));
    CascadeMux I__5139 (
            .O(N__29887),
            .I(N__29881));
    InMux I__5138 (
            .O(N__29884),
            .I(N__29878));
    InMux I__5137 (
            .O(N__29881),
            .I(N__29875));
    LocalMux I__5136 (
            .O(N__29878),
            .I(N__29872));
    LocalMux I__5135 (
            .O(N__29875),
            .I(N__29869));
    Span4Mux_v I__5134 (
            .O(N__29872),
            .I(N__29866));
    Span4Mux_v I__5133 (
            .O(N__29869),
            .I(N__29863));
    Span4Mux_v I__5132 (
            .O(N__29866),
            .I(N__29860));
    Span4Mux_h I__5131 (
            .O(N__29863),
            .I(N__29856));
    Span4Mux_v I__5130 (
            .O(N__29860),
            .I(N__29853));
    InMux I__5129 (
            .O(N__29859),
            .I(N__29850));
    Span4Mux_h I__5128 (
            .O(N__29856),
            .I(N__29847));
    Sp12to4 I__5127 (
            .O(N__29853),
            .I(N__29844));
    LocalMux I__5126 (
            .O(N__29850),
            .I(data_count_4));
    Odrv4 I__5125 (
            .O(N__29847),
            .I(data_count_4));
    Odrv12 I__5124 (
            .O(N__29844),
            .I(data_count_4));
    InMux I__5123 (
            .O(N__29837),
            .I(n19348));
    CascadeMux I__5122 (
            .O(N__29834),
            .I(N__29831));
    CascadeBuf I__5121 (
            .O(N__29831),
            .I(N__29828));
    CascadeMux I__5120 (
            .O(N__29828),
            .I(N__29825));
    CascadeBuf I__5119 (
            .O(N__29825),
            .I(N__29822));
    CascadeMux I__5118 (
            .O(N__29822),
            .I(N__29819));
    CascadeBuf I__5117 (
            .O(N__29819),
            .I(N__29816));
    CascadeMux I__5116 (
            .O(N__29816),
            .I(N__29813));
    CascadeBuf I__5115 (
            .O(N__29813),
            .I(N__29810));
    CascadeMux I__5114 (
            .O(N__29810),
            .I(N__29807));
    CascadeBuf I__5113 (
            .O(N__29807),
            .I(N__29804));
    CascadeMux I__5112 (
            .O(N__29804),
            .I(N__29801));
    CascadeBuf I__5111 (
            .O(N__29801),
            .I(N__29798));
    CascadeMux I__5110 (
            .O(N__29798),
            .I(N__29795));
    CascadeBuf I__5109 (
            .O(N__29795),
            .I(N__29792));
    CascadeMux I__5108 (
            .O(N__29792),
            .I(N__29789));
    CascadeBuf I__5107 (
            .O(N__29789),
            .I(N__29786));
    CascadeMux I__5106 (
            .O(N__29786),
            .I(N__29782));
    CascadeMux I__5105 (
            .O(N__29785),
            .I(N__29779));
    CascadeBuf I__5104 (
            .O(N__29782),
            .I(N__29776));
    CascadeBuf I__5103 (
            .O(N__29779),
            .I(N__29773));
    CascadeMux I__5102 (
            .O(N__29776),
            .I(N__29770));
    CascadeMux I__5101 (
            .O(N__29773),
            .I(N__29767));
    InMux I__5100 (
            .O(N__29770),
            .I(N__29764));
    InMux I__5099 (
            .O(N__29767),
            .I(N__29761));
    LocalMux I__5098 (
            .O(N__29764),
            .I(N__29758));
    LocalMux I__5097 (
            .O(N__29761),
            .I(N__29754));
    Sp12to4 I__5096 (
            .O(N__29758),
            .I(N__29751));
    InMux I__5095 (
            .O(N__29757),
            .I(N__29748));
    Span12Mux_h I__5094 (
            .O(N__29754),
            .I(N__29745));
    Span12Mux_v I__5093 (
            .O(N__29751),
            .I(N__29742));
    LocalMux I__5092 (
            .O(N__29748),
            .I(data_count_5));
    Odrv12 I__5091 (
            .O(N__29745),
            .I(data_count_5));
    Odrv12 I__5090 (
            .O(N__29742),
            .I(data_count_5));
    InMux I__5089 (
            .O(N__29735),
            .I(n19349));
    CascadeMux I__5088 (
            .O(N__29732),
            .I(N__29729));
    CascadeBuf I__5087 (
            .O(N__29729),
            .I(N__29726));
    CascadeMux I__5086 (
            .O(N__29726),
            .I(N__29723));
    CascadeBuf I__5085 (
            .O(N__29723),
            .I(N__29720));
    CascadeMux I__5084 (
            .O(N__29720),
            .I(N__29717));
    CascadeBuf I__5083 (
            .O(N__29717),
            .I(N__29714));
    CascadeMux I__5082 (
            .O(N__29714),
            .I(N__29711));
    CascadeBuf I__5081 (
            .O(N__29711),
            .I(N__29708));
    CascadeMux I__5080 (
            .O(N__29708),
            .I(N__29705));
    CascadeBuf I__5079 (
            .O(N__29705),
            .I(N__29702));
    CascadeMux I__5078 (
            .O(N__29702),
            .I(N__29699));
    CascadeBuf I__5077 (
            .O(N__29699),
            .I(N__29696));
    CascadeMux I__5076 (
            .O(N__29696),
            .I(N__29693));
    CascadeBuf I__5075 (
            .O(N__29693),
            .I(N__29690));
    CascadeMux I__5074 (
            .O(N__29690),
            .I(N__29686));
    CascadeMux I__5073 (
            .O(N__29689),
            .I(N__29683));
    CascadeBuf I__5072 (
            .O(N__29686),
            .I(N__29680));
    CascadeBuf I__5071 (
            .O(N__29683),
            .I(N__29677));
    CascadeMux I__5070 (
            .O(N__29680),
            .I(N__29674));
    CascadeMux I__5069 (
            .O(N__29677),
            .I(N__29671));
    CascadeBuf I__5068 (
            .O(N__29674),
            .I(N__29668));
    InMux I__5067 (
            .O(N__29671),
            .I(N__29665));
    CascadeMux I__5066 (
            .O(N__29668),
            .I(N__29662));
    LocalMux I__5065 (
            .O(N__29665),
            .I(N__29659));
    InMux I__5064 (
            .O(N__29662),
            .I(N__29656));
    Span4Mux_h I__5063 (
            .O(N__29659),
            .I(N__29653));
    LocalMux I__5062 (
            .O(N__29656),
            .I(N__29650));
    Span4Mux_v I__5061 (
            .O(N__29653),
            .I(N__29646));
    Sp12to4 I__5060 (
            .O(N__29650),
            .I(N__29643));
    InMux I__5059 (
            .O(N__29649),
            .I(N__29640));
    Span4Mux_h I__5058 (
            .O(N__29646),
            .I(N__29637));
    Span12Mux_v I__5057 (
            .O(N__29643),
            .I(N__29634));
    LocalMux I__5056 (
            .O(N__29640),
            .I(data_count_6));
    Odrv4 I__5055 (
            .O(N__29637),
            .I(data_count_6));
    Odrv12 I__5054 (
            .O(N__29634),
            .I(data_count_6));
    InMux I__5053 (
            .O(N__29627),
            .I(n19350));
    CascadeMux I__5052 (
            .O(N__29624),
            .I(N__29621));
    CascadeBuf I__5051 (
            .O(N__29621),
            .I(N__29618));
    CascadeMux I__5050 (
            .O(N__29618),
            .I(N__29615));
    CascadeBuf I__5049 (
            .O(N__29615),
            .I(N__29612));
    CascadeMux I__5048 (
            .O(N__29612),
            .I(N__29609));
    CascadeBuf I__5047 (
            .O(N__29609),
            .I(N__29606));
    CascadeMux I__5046 (
            .O(N__29606),
            .I(N__29603));
    CascadeBuf I__5045 (
            .O(N__29603),
            .I(N__29600));
    CascadeMux I__5044 (
            .O(N__29600),
            .I(N__29597));
    CascadeBuf I__5043 (
            .O(N__29597),
            .I(N__29594));
    CascadeMux I__5042 (
            .O(N__29594),
            .I(N__29591));
    CascadeBuf I__5041 (
            .O(N__29591),
            .I(N__29588));
    CascadeMux I__5040 (
            .O(N__29588),
            .I(N__29585));
    CascadeBuf I__5039 (
            .O(N__29585),
            .I(N__29582));
    CascadeMux I__5038 (
            .O(N__29582),
            .I(N__29579));
    CascadeBuf I__5037 (
            .O(N__29579),
            .I(N__29575));
    CascadeMux I__5036 (
            .O(N__29578),
            .I(N__29572));
    CascadeMux I__5035 (
            .O(N__29575),
            .I(N__29569));
    CascadeBuf I__5034 (
            .O(N__29572),
            .I(N__29566));
    CascadeBuf I__5033 (
            .O(N__29569),
            .I(N__29563));
    CascadeMux I__5032 (
            .O(N__29566),
            .I(N__29560));
    CascadeMux I__5031 (
            .O(N__29563),
            .I(N__29557));
    InMux I__5030 (
            .O(N__29560),
            .I(N__29554));
    InMux I__5029 (
            .O(N__29557),
            .I(N__29551));
    LocalMux I__5028 (
            .O(N__29554),
            .I(N__29548));
    LocalMux I__5027 (
            .O(N__29551),
            .I(N__29545));
    Span4Mux_h I__5026 (
            .O(N__29548),
            .I(N__29542));
    Span4Mux_h I__5025 (
            .O(N__29545),
            .I(N__29539));
    Sp12to4 I__5024 (
            .O(N__29542),
            .I(N__29535));
    Sp12to4 I__5023 (
            .O(N__29539),
            .I(N__29532));
    InMux I__5022 (
            .O(N__29538),
            .I(N__29529));
    Span12Mux_v I__5021 (
            .O(N__29535),
            .I(N__29524));
    Span12Mux_v I__5020 (
            .O(N__29532),
            .I(N__29524));
    LocalMux I__5019 (
            .O(N__29529),
            .I(data_count_7));
    Odrv12 I__5018 (
            .O(N__29524),
            .I(data_count_7));
    InMux I__5017 (
            .O(N__29519),
            .I(n19351));
    CascadeMux I__5016 (
            .O(N__29516),
            .I(N__29512));
    CascadeMux I__5015 (
            .O(N__29515),
            .I(N__29509));
    InMux I__5014 (
            .O(N__29512),
            .I(N__29505));
    InMux I__5013 (
            .O(N__29509),
            .I(N__29502));
    CascadeMux I__5012 (
            .O(N__29508),
            .I(N__29499));
    LocalMux I__5011 (
            .O(N__29505),
            .I(N__29496));
    LocalMux I__5010 (
            .O(N__29502),
            .I(N__29492));
    InMux I__5009 (
            .O(N__29499),
            .I(N__29489));
    Span4Mux_v I__5008 (
            .O(N__29496),
            .I(N__29485));
    InMux I__5007 (
            .O(N__29495),
            .I(N__29482));
    Span4Mux_v I__5006 (
            .O(N__29492),
            .I(N__29479));
    LocalMux I__5005 (
            .O(N__29489),
            .I(N__29476));
    InMux I__5004 (
            .O(N__29488),
            .I(N__29473));
    Span4Mux_h I__5003 (
            .O(N__29485),
            .I(N__29468));
    LocalMux I__5002 (
            .O(N__29482),
            .I(N__29468));
    Odrv4 I__5001 (
            .O(N__29479),
            .I(buf_cfgRTD_6));
    Odrv12 I__5000 (
            .O(N__29476),
            .I(buf_cfgRTD_6));
    LocalMux I__4999 (
            .O(N__29473),
            .I(buf_cfgRTD_6));
    Odrv4 I__4998 (
            .O(N__29468),
            .I(buf_cfgRTD_6));
    InMux I__4997 (
            .O(N__29459),
            .I(N__29456));
    LocalMux I__4996 (
            .O(N__29456),
            .I(N__29453));
    Span4Mux_v I__4995 (
            .O(N__29453),
            .I(N__29448));
    CascadeMux I__4994 (
            .O(N__29452),
            .I(N__29445));
    CascadeMux I__4993 (
            .O(N__29451),
            .I(N__29442));
    Span4Mux_h I__4992 (
            .O(N__29448),
            .I(N__29439));
    InMux I__4991 (
            .O(N__29445),
            .I(N__29434));
    InMux I__4990 (
            .O(N__29442),
            .I(N__29434));
    Odrv4 I__4989 (
            .O(N__29439),
            .I(cmd_rdadctmp_27));
    LocalMux I__4988 (
            .O(N__29434),
            .I(cmd_rdadctmp_27));
    InMux I__4987 (
            .O(N__29429),
            .I(N__29425));
    InMux I__4986 (
            .O(N__29428),
            .I(N__29422));
    LocalMux I__4985 (
            .O(N__29425),
            .I(N__29418));
    LocalMux I__4984 (
            .O(N__29422),
            .I(N__29415));
    InMux I__4983 (
            .O(N__29421),
            .I(N__29412));
    Span12Mux_h I__4982 (
            .O(N__29418),
            .I(N__29409));
    Span4Mux_h I__4981 (
            .O(N__29415),
            .I(N__29406));
    LocalMux I__4980 (
            .O(N__29412),
            .I(buf_adcdata_vac_19));
    Odrv12 I__4979 (
            .O(N__29409),
            .I(buf_adcdata_vac_19));
    Odrv4 I__4978 (
            .O(N__29406),
            .I(buf_adcdata_vac_19));
    InMux I__4977 (
            .O(N__29399),
            .I(N__29395));
    CascadeMux I__4976 (
            .O(N__29398),
            .I(N__29391));
    LocalMux I__4975 (
            .O(N__29395),
            .I(N__29388));
    CascadeMux I__4974 (
            .O(N__29394),
            .I(N__29385));
    InMux I__4973 (
            .O(N__29391),
            .I(N__29382));
    Span12Mux_h I__4972 (
            .O(N__29388),
            .I(N__29379));
    InMux I__4971 (
            .O(N__29385),
            .I(N__29376));
    LocalMux I__4970 (
            .O(N__29382),
            .I(cmd_rdadctmp_8_adj_1442));
    Odrv12 I__4969 (
            .O(N__29379),
            .I(cmd_rdadctmp_8_adj_1442));
    LocalMux I__4968 (
            .O(N__29376),
            .I(cmd_rdadctmp_8_adj_1442));
    CascadeMux I__4967 (
            .O(N__29369),
            .I(N__29366));
    InMux I__4966 (
            .O(N__29366),
            .I(N__29359));
    InMux I__4965 (
            .O(N__29365),
            .I(N__29359));
    CascadeMux I__4964 (
            .O(N__29364),
            .I(N__29356));
    LocalMux I__4963 (
            .O(N__29359),
            .I(N__29353));
    InMux I__4962 (
            .O(N__29356),
            .I(N__29350));
    Odrv4 I__4961 (
            .O(N__29353),
            .I(cmd_rdadctmp_9_adj_1441));
    LocalMux I__4960 (
            .O(N__29350),
            .I(cmd_rdadctmp_9_adj_1441));
    InMux I__4959 (
            .O(N__29345),
            .I(N__29342));
    LocalMux I__4958 (
            .O(N__29342),
            .I(N__29338));
    CascadeMux I__4957 (
            .O(N__29341),
            .I(N__29335));
    Span4Mux_v I__4956 (
            .O(N__29338),
            .I(N__29332));
    InMux I__4955 (
            .O(N__29335),
            .I(N__29329));
    Odrv4 I__4954 (
            .O(N__29332),
            .I(buf_adcdata_vdc_15));
    LocalMux I__4953 (
            .O(N__29329),
            .I(buf_adcdata_vdc_15));
    InMux I__4952 (
            .O(N__29324),
            .I(N__29321));
    LocalMux I__4951 (
            .O(N__29321),
            .I(N__29318));
    Span4Mux_v I__4950 (
            .O(N__29318),
            .I(N__29315));
    Span4Mux_h I__4949 (
            .O(N__29315),
            .I(N__29312));
    Span4Mux_h I__4948 (
            .O(N__29312),
            .I(N__29307));
    InMux I__4947 (
            .O(N__29311),
            .I(N__29302));
    InMux I__4946 (
            .O(N__29310),
            .I(N__29302));
    Odrv4 I__4945 (
            .O(N__29307),
            .I(buf_adcdata_vac_15));
    LocalMux I__4944 (
            .O(N__29302),
            .I(buf_adcdata_vac_15));
    InMux I__4943 (
            .O(N__29297),
            .I(N__29294));
    LocalMux I__4942 (
            .O(N__29294),
            .I(N__29291));
    Span4Mux_h I__4941 (
            .O(N__29291),
            .I(N__29288));
    Odrv4 I__4940 (
            .O(N__29288),
            .I(n22016));
    CascadeMux I__4939 (
            .O(N__29285),
            .I(N__29282));
    InMux I__4938 (
            .O(N__29282),
            .I(N__29279));
    LocalMux I__4937 (
            .O(N__29279),
            .I(N__29275));
    CascadeMux I__4936 (
            .O(N__29278),
            .I(N__29272));
    Span4Mux_v I__4935 (
            .O(N__29275),
            .I(N__29269));
    InMux I__4934 (
            .O(N__29272),
            .I(N__29266));
    Odrv4 I__4933 (
            .O(N__29269),
            .I(buf_adcdata_vdc_16));
    LocalMux I__4932 (
            .O(N__29266),
            .I(buf_adcdata_vdc_16));
    CascadeMux I__4931 (
            .O(N__29261),
            .I(N__29257));
    CascadeMux I__4930 (
            .O(N__29260),
            .I(N__29253));
    InMux I__4929 (
            .O(N__29257),
            .I(N__29250));
    InMux I__4928 (
            .O(N__29256),
            .I(N__29245));
    InMux I__4927 (
            .O(N__29253),
            .I(N__29245));
    LocalMux I__4926 (
            .O(N__29250),
            .I(cmd_rdadctmp_23));
    LocalMux I__4925 (
            .O(N__29245),
            .I(cmd_rdadctmp_23));
    CascadeMux I__4924 (
            .O(N__29240),
            .I(N__29235));
    InMux I__4923 (
            .O(N__29239),
            .I(N__29232));
    InMux I__4922 (
            .O(N__29238),
            .I(N__29229));
    InMux I__4921 (
            .O(N__29235),
            .I(N__29226));
    LocalMux I__4920 (
            .O(N__29232),
            .I(N__29223));
    LocalMux I__4919 (
            .O(N__29229),
            .I(cmd_rdadctmp_24));
    LocalMux I__4918 (
            .O(N__29226),
            .I(cmd_rdadctmp_24));
    Odrv4 I__4917 (
            .O(N__29223),
            .I(cmd_rdadctmp_24));
    InMux I__4916 (
            .O(N__29216),
            .I(N__29212));
    InMux I__4915 (
            .O(N__29215),
            .I(N__29209));
    LocalMux I__4914 (
            .O(N__29212),
            .I(cmd_rdadcbuf_27));
    LocalMux I__4913 (
            .O(N__29209),
            .I(cmd_rdadcbuf_27));
    InMux I__4912 (
            .O(N__29204),
            .I(N__29201));
    LocalMux I__4911 (
            .O(N__29201),
            .I(N__29197));
    InMux I__4910 (
            .O(N__29200),
            .I(N__29194));
    Odrv4 I__4909 (
            .O(N__29197),
            .I(cmd_rdadcbuf_11));
    LocalMux I__4908 (
            .O(N__29194),
            .I(cmd_rdadcbuf_11));
    InMux I__4907 (
            .O(N__29189),
            .I(N__29185));
    InMux I__4906 (
            .O(N__29188),
            .I(N__29182));
    LocalMux I__4905 (
            .O(N__29185),
            .I(cmd_rdadcbuf_33));
    LocalMux I__4904 (
            .O(N__29182),
            .I(cmd_rdadcbuf_33));
    CascadeMux I__4903 (
            .O(N__29177),
            .I(N__29174));
    InMux I__4902 (
            .O(N__29174),
            .I(N__29154));
    InMux I__4901 (
            .O(N__29173),
            .I(N__29154));
    CascadeMux I__4900 (
            .O(N__29172),
            .I(N__29151));
    InMux I__4899 (
            .O(N__29171),
            .I(N__29147));
    InMux I__4898 (
            .O(N__29170),
            .I(N__29132));
    InMux I__4897 (
            .O(N__29169),
            .I(N__29132));
    InMux I__4896 (
            .O(N__29168),
            .I(N__29132));
    InMux I__4895 (
            .O(N__29167),
            .I(N__29132));
    InMux I__4894 (
            .O(N__29166),
            .I(N__29132));
    InMux I__4893 (
            .O(N__29165),
            .I(N__29132));
    InMux I__4892 (
            .O(N__29164),
            .I(N__29132));
    CascadeMux I__4891 (
            .O(N__29163),
            .I(N__29128));
    CascadeMux I__4890 (
            .O(N__29162),
            .I(N__29121));
    CascadeMux I__4889 (
            .O(N__29161),
            .I(N__29118));
    CascadeMux I__4888 (
            .O(N__29160),
            .I(N__29115));
    CascadeMux I__4887 (
            .O(N__29159),
            .I(N__29112));
    LocalMux I__4886 (
            .O(N__29154),
            .I(N__29107));
    InMux I__4885 (
            .O(N__29151),
            .I(N__29102));
    InMux I__4884 (
            .O(N__29150),
            .I(N__29102));
    LocalMux I__4883 (
            .O(N__29147),
            .I(N__29099));
    LocalMux I__4882 (
            .O(N__29132),
            .I(N__29096));
    InMux I__4881 (
            .O(N__29131),
            .I(N__29093));
    InMux I__4880 (
            .O(N__29128),
            .I(N__29090));
    InMux I__4879 (
            .O(N__29127),
            .I(N__29073));
    InMux I__4878 (
            .O(N__29126),
            .I(N__29073));
    InMux I__4877 (
            .O(N__29125),
            .I(N__29073));
    InMux I__4876 (
            .O(N__29124),
            .I(N__29073));
    InMux I__4875 (
            .O(N__29121),
            .I(N__29073));
    InMux I__4874 (
            .O(N__29118),
            .I(N__29073));
    InMux I__4873 (
            .O(N__29115),
            .I(N__29073));
    InMux I__4872 (
            .O(N__29112),
            .I(N__29073));
    InMux I__4871 (
            .O(N__29111),
            .I(N__29068));
    InMux I__4870 (
            .O(N__29110),
            .I(N__29068));
    Span4Mux_v I__4869 (
            .O(N__29107),
            .I(N__29065));
    LocalMux I__4868 (
            .O(N__29102),
            .I(N__29058));
    Span4Mux_h I__4867 (
            .O(N__29099),
            .I(N__29058));
    Span4Mux_h I__4866 (
            .O(N__29096),
            .I(N__29058));
    LocalMux I__4865 (
            .O(N__29093),
            .I(n13109));
    LocalMux I__4864 (
            .O(N__29090),
            .I(n13109));
    LocalMux I__4863 (
            .O(N__29073),
            .I(n13109));
    LocalMux I__4862 (
            .O(N__29068),
            .I(n13109));
    Odrv4 I__4861 (
            .O(N__29065),
            .I(n13109));
    Odrv4 I__4860 (
            .O(N__29058),
            .I(n13109));
    InMux I__4859 (
            .O(N__29045),
            .I(N__29041));
    InMux I__4858 (
            .O(N__29044),
            .I(N__29038));
    LocalMux I__4857 (
            .O(N__29041),
            .I(cmd_rdadcbuf_20));
    LocalMux I__4856 (
            .O(N__29038),
            .I(cmd_rdadcbuf_20));
    InMux I__4855 (
            .O(N__29033),
            .I(N__29030));
    LocalMux I__4854 (
            .O(N__29030),
            .I(N__29025));
    InMux I__4853 (
            .O(N__29029),
            .I(N__29022));
    InMux I__4852 (
            .O(N__29028),
            .I(N__29019));
    Span12Mux_h I__4851 (
            .O(N__29025),
            .I(N__29016));
    LocalMux I__4850 (
            .O(N__29022),
            .I(N__29013));
    LocalMux I__4849 (
            .O(N__29019),
            .I(buf_adcdata_vac_18));
    Odrv12 I__4848 (
            .O(N__29016),
            .I(buf_adcdata_vac_18));
    Odrv4 I__4847 (
            .O(N__29013),
            .I(buf_adcdata_vac_18));
    InMux I__4846 (
            .O(N__29006),
            .I(N__29002));
    InMux I__4845 (
            .O(N__29005),
            .I(N__28997));
    LocalMux I__4844 (
            .O(N__29002),
            .I(N__28991));
    InMux I__4843 (
            .O(N__29001),
            .I(N__28986));
    InMux I__4842 (
            .O(N__29000),
            .I(N__28986));
    LocalMux I__4841 (
            .O(N__28997),
            .I(N__28983));
    InMux I__4840 (
            .O(N__28996),
            .I(N__28980));
    InMux I__4839 (
            .O(N__28995),
            .I(N__28974));
    InMux I__4838 (
            .O(N__28994),
            .I(N__28974));
    Span4Mux_h I__4837 (
            .O(N__28991),
            .I(N__28969));
    LocalMux I__4836 (
            .O(N__28986),
            .I(N__28969));
    Span4Mux_v I__4835 (
            .O(N__28983),
            .I(N__28964));
    LocalMux I__4834 (
            .O(N__28980),
            .I(N__28964));
    InMux I__4833 (
            .O(N__28979),
            .I(N__28961));
    LocalMux I__4832 (
            .O(N__28974),
            .I(N__28958));
    Span4Mux_v I__4831 (
            .O(N__28969),
            .I(N__28955));
    Span4Mux_h I__4830 (
            .O(N__28964),
            .I(N__28952));
    LocalMux I__4829 (
            .O(N__28961),
            .I(N__28947));
    Span4Mux_h I__4828 (
            .O(N__28958),
            .I(N__28947));
    Odrv4 I__4827 (
            .O(N__28955),
            .I(n12411));
    Odrv4 I__4826 (
            .O(N__28952),
            .I(n12411));
    Odrv4 I__4825 (
            .O(N__28947),
            .I(n12411));
    CascadeMux I__4824 (
            .O(N__28940),
            .I(n30_adj_1480_cascade_));
    InMux I__4823 (
            .O(N__28937),
            .I(N__28934));
    LocalMux I__4822 (
            .O(N__28934),
            .I(N__28930));
    CascadeMux I__4821 (
            .O(N__28933),
            .I(N__28927));
    Span4Mux_v I__4820 (
            .O(N__28930),
            .I(N__28924));
    InMux I__4819 (
            .O(N__28927),
            .I(N__28921));
    Odrv4 I__4818 (
            .O(N__28924),
            .I(buf_adcdata_vdc_1));
    LocalMux I__4817 (
            .O(N__28921),
            .I(buf_adcdata_vdc_1));
    CascadeMux I__4816 (
            .O(N__28916),
            .I(n19_adj_1491_cascade_));
    InMux I__4815 (
            .O(N__28913),
            .I(N__28910));
    LocalMux I__4814 (
            .O(N__28910),
            .I(N__28907));
    Span12Mux_h I__4813 (
            .O(N__28907),
            .I(N__28902));
    InMux I__4812 (
            .O(N__28906),
            .I(N__28897));
    InMux I__4811 (
            .O(N__28905),
            .I(N__28897));
    Odrv12 I__4810 (
            .O(N__28902),
            .I(buf_adcdata_iac_1));
    LocalMux I__4809 (
            .O(N__28897),
            .I(buf_adcdata_iac_1));
    CascadeMux I__4808 (
            .O(N__28892),
            .I(N__28889));
    InMux I__4807 (
            .O(N__28889),
            .I(N__28886));
    LocalMux I__4806 (
            .O(N__28886),
            .I(N__28882));
    InMux I__4805 (
            .O(N__28885),
            .I(N__28879));
    Span4Mux_v I__4804 (
            .O(N__28882),
            .I(N__28874));
    LocalMux I__4803 (
            .O(N__28879),
            .I(N__28874));
    Odrv4 I__4802 (
            .O(N__28874),
            .I(buf_readRTD_14));
    InMux I__4801 (
            .O(N__28871),
            .I(N__28867));
    InMux I__4800 (
            .O(N__28870),
            .I(N__28864));
    LocalMux I__4799 (
            .O(N__28867),
            .I(cmd_rdadcbuf_26));
    LocalMux I__4798 (
            .O(N__28864),
            .I(cmd_rdadcbuf_26));
    InMux I__4797 (
            .O(N__28859),
            .I(N__28855));
    InMux I__4796 (
            .O(N__28858),
            .I(N__28852));
    LocalMux I__4795 (
            .O(N__28855),
            .I(cmd_rdadcbuf_25));
    LocalMux I__4794 (
            .O(N__28852),
            .I(cmd_rdadcbuf_25));
    InMux I__4793 (
            .O(N__28847),
            .I(N__28843));
    InMux I__4792 (
            .O(N__28846),
            .I(N__28840));
    LocalMux I__4791 (
            .O(N__28843),
            .I(cmd_rdadcbuf_24));
    LocalMux I__4790 (
            .O(N__28840),
            .I(cmd_rdadcbuf_24));
    CascadeMux I__4789 (
            .O(N__28835),
            .I(N__28831));
    CascadeMux I__4788 (
            .O(N__28834),
            .I(N__28828));
    InMux I__4787 (
            .O(N__28831),
            .I(N__28825));
    InMux I__4786 (
            .O(N__28828),
            .I(N__28821));
    LocalMux I__4785 (
            .O(N__28825),
            .I(N__28818));
    CascadeMux I__4784 (
            .O(N__28824),
            .I(N__28815));
    LocalMux I__4783 (
            .O(N__28821),
            .I(N__28810));
    Span4Mux_h I__4782 (
            .O(N__28818),
            .I(N__28810));
    InMux I__4781 (
            .O(N__28815),
            .I(N__28807));
    Odrv4 I__4780 (
            .O(N__28810),
            .I(cmd_rdadctmp_11));
    LocalMux I__4779 (
            .O(N__28807),
            .I(cmd_rdadctmp_11));
    InMux I__4778 (
            .O(N__28802),
            .I(N__28799));
    LocalMux I__4777 (
            .O(N__28799),
            .I(N__28796));
    Span12Mux_h I__4776 (
            .O(N__28796),
            .I(N__28791));
    InMux I__4775 (
            .O(N__28795),
            .I(N__28786));
    InMux I__4774 (
            .O(N__28794),
            .I(N__28786));
    Odrv12 I__4773 (
            .O(N__28791),
            .I(buf_adcdata_vac_3));
    LocalMux I__4772 (
            .O(N__28786),
            .I(buf_adcdata_vac_3));
    CascadeMux I__4771 (
            .O(N__28781),
            .I(N__28777));
    CascadeMux I__4770 (
            .O(N__28780),
            .I(N__28773));
    InMux I__4769 (
            .O(N__28777),
            .I(N__28766));
    InMux I__4768 (
            .O(N__28776),
            .I(N__28766));
    InMux I__4767 (
            .O(N__28773),
            .I(N__28766));
    LocalMux I__4766 (
            .O(N__28766),
            .I(cmd_rdadctmp_11_adj_1439));
    CascadeMux I__4765 (
            .O(N__28763),
            .I(N__28759));
    CascadeMux I__4764 (
            .O(N__28762),
            .I(N__28756));
    InMux I__4763 (
            .O(N__28759),
            .I(N__28752));
    InMux I__4762 (
            .O(N__28756),
            .I(N__28749));
    CascadeMux I__4761 (
            .O(N__28755),
            .I(N__28746));
    LocalMux I__4760 (
            .O(N__28752),
            .I(N__28743));
    LocalMux I__4759 (
            .O(N__28749),
            .I(N__28740));
    InMux I__4758 (
            .O(N__28746),
            .I(N__28737));
    Span4Mux_h I__4757 (
            .O(N__28743),
            .I(N__28734));
    Span4Mux_v I__4756 (
            .O(N__28740),
            .I(N__28731));
    LocalMux I__4755 (
            .O(N__28737),
            .I(cmd_rdadctmp_12_adj_1438));
    Odrv4 I__4754 (
            .O(N__28734),
            .I(cmd_rdadctmp_12_adj_1438));
    Odrv4 I__4753 (
            .O(N__28731),
            .I(cmd_rdadctmp_12_adj_1438));
    InMux I__4752 (
            .O(N__28724),
            .I(N__28721));
    LocalMux I__4751 (
            .O(N__28721),
            .I(N__28718));
    Span4Mux_v I__4750 (
            .O(N__28718),
            .I(N__28715));
    Span4Mux_h I__4749 (
            .O(N__28715),
            .I(N__28712));
    Span4Mux_h I__4748 (
            .O(N__28712),
            .I(N__28709));
    Odrv4 I__4747 (
            .O(N__28709),
            .I(buf_data_vac_7));
    InMux I__4746 (
            .O(N__28706),
            .I(N__28703));
    LocalMux I__4745 (
            .O(N__28703),
            .I(N__28700));
    Span4Mux_v I__4744 (
            .O(N__28700),
            .I(N__28697));
    Span4Mux_h I__4743 (
            .O(N__28697),
            .I(N__28694));
    Odrv4 I__4742 (
            .O(N__28694),
            .I(buf_data_vac_6));
    InMux I__4741 (
            .O(N__28691),
            .I(N__28688));
    LocalMux I__4740 (
            .O(N__28688),
            .I(N__28685));
    Span4Mux_h I__4739 (
            .O(N__28685),
            .I(N__28682));
    Span4Mux_h I__4738 (
            .O(N__28682),
            .I(N__28679));
    Odrv4 I__4737 (
            .O(N__28679),
            .I(buf_data_vac_5));
    CascadeMux I__4736 (
            .O(N__28676),
            .I(N__28673));
    InMux I__4735 (
            .O(N__28673),
            .I(N__28670));
    LocalMux I__4734 (
            .O(N__28670),
            .I(N__28665));
    InMux I__4733 (
            .O(N__28669),
            .I(N__28662));
    CascadeMux I__4732 (
            .O(N__28668),
            .I(N__28659));
    Span4Mux_v I__4731 (
            .O(N__28665),
            .I(N__28656));
    LocalMux I__4730 (
            .O(N__28662),
            .I(N__28653));
    InMux I__4729 (
            .O(N__28659),
            .I(N__28650));
    Odrv4 I__4728 (
            .O(N__28656),
            .I(cmd_rdadctmp_10_adj_1440));
    Odrv12 I__4727 (
            .O(N__28653),
            .I(cmd_rdadctmp_10_adj_1440));
    LocalMux I__4726 (
            .O(N__28650),
            .I(cmd_rdadctmp_10_adj_1440));
    InMux I__4725 (
            .O(N__28643),
            .I(N__28640));
    LocalMux I__4724 (
            .O(N__28640),
            .I(N__28637));
    Span4Mux_h I__4723 (
            .O(N__28637),
            .I(N__28633));
    CascadeMux I__4722 (
            .O(N__28636),
            .I(N__28630));
    Span4Mux_h I__4721 (
            .O(N__28633),
            .I(N__28627));
    InMux I__4720 (
            .O(N__28630),
            .I(N__28624));
    Odrv4 I__4719 (
            .O(N__28627),
            .I(buf_adcdata_vdc_2));
    LocalMux I__4718 (
            .O(N__28624),
            .I(buf_adcdata_vdc_2));
    InMux I__4717 (
            .O(N__28619),
            .I(N__28616));
    LocalMux I__4716 (
            .O(N__28616),
            .I(N__28613));
    Span4Mux_v I__4715 (
            .O(N__28613),
            .I(N__28610));
    Span4Mux_h I__4714 (
            .O(N__28610),
            .I(N__28607));
    Span4Mux_h I__4713 (
            .O(N__28607),
            .I(N__28602));
    InMux I__4712 (
            .O(N__28606),
            .I(N__28597));
    InMux I__4711 (
            .O(N__28605),
            .I(N__28597));
    Odrv4 I__4710 (
            .O(N__28602),
            .I(buf_adcdata_vac_2));
    LocalMux I__4709 (
            .O(N__28597),
            .I(buf_adcdata_vac_2));
    InMux I__4708 (
            .O(N__28592),
            .I(N__28589));
    LocalMux I__4707 (
            .O(N__28589),
            .I(N__28586));
    Span4Mux_v I__4706 (
            .O(N__28586),
            .I(N__28582));
    InMux I__4705 (
            .O(N__28585),
            .I(N__28578));
    Sp12to4 I__4704 (
            .O(N__28582),
            .I(N__28575));
    InMux I__4703 (
            .O(N__28581),
            .I(N__28572));
    LocalMux I__4702 (
            .O(N__28578),
            .I(buf_adcdata_iac_2));
    Odrv12 I__4701 (
            .O(N__28575),
            .I(buf_adcdata_iac_2));
    LocalMux I__4700 (
            .O(N__28572),
            .I(buf_adcdata_iac_2));
    CascadeMux I__4699 (
            .O(N__28565),
            .I(n19_adj_1646_cascade_));
    InMux I__4698 (
            .O(N__28562),
            .I(N__28559));
    LocalMux I__4697 (
            .O(N__28559),
            .I(N__28556));
    Span4Mux_h I__4696 (
            .O(N__28556),
            .I(N__28553));
    Span4Mux_h I__4695 (
            .O(N__28553),
            .I(N__28550));
    Span4Mux_h I__4694 (
            .O(N__28550),
            .I(N__28547));
    Odrv4 I__4693 (
            .O(N__28547),
            .I(buf_data_iac_2));
    CascadeMux I__4692 (
            .O(N__28544),
            .I(n22_adj_1647_cascade_));
    CascadeMux I__4691 (
            .O(N__28541),
            .I(N__28538));
    InMux I__4690 (
            .O(N__28538),
            .I(N__28532));
    InMux I__4689 (
            .O(N__28537),
            .I(N__28532));
    LocalMux I__4688 (
            .O(N__28532),
            .I(N__28528));
    CascadeMux I__4687 (
            .O(N__28531),
            .I(N__28525));
    Span4Mux_v I__4686 (
            .O(N__28528),
            .I(N__28522));
    InMux I__4685 (
            .O(N__28525),
            .I(N__28519));
    Odrv4 I__4684 (
            .O(N__28522),
            .I(cmd_rdadctmp_10));
    LocalMux I__4683 (
            .O(N__28519),
            .I(cmd_rdadctmp_10));
    InMux I__4682 (
            .O(N__28514),
            .I(N__28511));
    LocalMux I__4681 (
            .O(N__28511),
            .I(N__28507));
    InMux I__4680 (
            .O(N__28510),
            .I(N__28504));
    Span4Mux_v I__4679 (
            .O(N__28507),
            .I(N__28501));
    LocalMux I__4678 (
            .O(N__28504),
            .I(N__28498));
    Odrv4 I__4677 (
            .O(N__28501),
            .I(buf_adcdata_vdc_3));
    Odrv4 I__4676 (
            .O(N__28498),
            .I(buf_adcdata_vdc_3));
    CascadeMux I__4675 (
            .O(N__28493),
            .I(n19_adj_1642_cascade_));
    InMux I__4674 (
            .O(N__28490),
            .I(N__28487));
    LocalMux I__4673 (
            .O(N__28487),
            .I(N__28484));
    Span4Mux_h I__4672 (
            .O(N__28484),
            .I(N__28481));
    Span4Mux_h I__4671 (
            .O(N__28481),
            .I(N__28478));
    Odrv4 I__4670 (
            .O(N__28478),
            .I(buf_data_iac_3));
    CascadeMux I__4669 (
            .O(N__28475),
            .I(n22_adj_1643_cascade_));
    InMux I__4668 (
            .O(N__28472),
            .I(N__28469));
    LocalMux I__4667 (
            .O(N__28469),
            .I(N__28466));
    Span12Mux_h I__4666 (
            .O(N__28466),
            .I(N__28461));
    InMux I__4665 (
            .O(N__28465),
            .I(N__28456));
    InMux I__4664 (
            .O(N__28464),
            .I(N__28456));
    Odrv12 I__4663 (
            .O(N__28461),
            .I(buf_adcdata_iac_3));
    LocalMux I__4662 (
            .O(N__28456),
            .I(buf_adcdata_iac_3));
    CascadeMux I__4661 (
            .O(N__28451),
            .I(N__28448));
    InMux I__4660 (
            .O(N__28448),
            .I(N__28445));
    LocalMux I__4659 (
            .O(N__28445),
            .I(\SIG_DDS.tmp_buf_5 ));
    InMux I__4658 (
            .O(N__28442),
            .I(N__28437));
    InMux I__4657 (
            .O(N__28441),
            .I(N__28434));
    InMux I__4656 (
            .O(N__28440),
            .I(N__28431));
    LocalMux I__4655 (
            .O(N__28437),
            .I(N__28428));
    LocalMux I__4654 (
            .O(N__28434),
            .I(buf_dds0_2));
    LocalMux I__4653 (
            .O(N__28431),
            .I(buf_dds0_2));
    Odrv4 I__4652 (
            .O(N__28428),
            .I(buf_dds0_2));
    CascadeMux I__4651 (
            .O(N__28421),
            .I(N__28418));
    InMux I__4650 (
            .O(N__28418),
            .I(N__28415));
    LocalMux I__4649 (
            .O(N__28415),
            .I(N__28410));
    InMux I__4648 (
            .O(N__28414),
            .I(N__28407));
    InMux I__4647 (
            .O(N__28413),
            .I(N__28404));
    Span4Mux_h I__4646 (
            .O(N__28410),
            .I(N__28401));
    LocalMux I__4645 (
            .O(N__28407),
            .I(N__28398));
    LocalMux I__4644 (
            .O(N__28404),
            .I(buf_dds0_4));
    Odrv4 I__4643 (
            .O(N__28401),
            .I(buf_dds0_4));
    Odrv4 I__4642 (
            .O(N__28398),
            .I(buf_dds0_4));
    CascadeMux I__4641 (
            .O(N__28391),
            .I(N__28388));
    InMux I__4640 (
            .O(N__28388),
            .I(N__28385));
    LocalMux I__4639 (
            .O(N__28385),
            .I(\SIG_DDS.tmp_buf_4 ));
    CascadeMux I__4638 (
            .O(N__28382),
            .I(N__28379));
    InMux I__4637 (
            .O(N__28379),
            .I(N__28376));
    LocalMux I__4636 (
            .O(N__28376),
            .I(\SIG_DDS.tmp_buf_7 ));
    InMux I__4635 (
            .O(N__28373),
            .I(N__28369));
    CascadeMux I__4634 (
            .O(N__28372),
            .I(N__28365));
    LocalMux I__4633 (
            .O(N__28369),
            .I(N__28362));
    InMux I__4632 (
            .O(N__28368),
            .I(N__28357));
    InMux I__4631 (
            .O(N__28365),
            .I(N__28357));
    Odrv4 I__4630 (
            .O(N__28362),
            .I(buf_dds0_8));
    LocalMux I__4629 (
            .O(N__28357),
            .I(buf_dds0_8));
    CascadeMux I__4628 (
            .O(N__28352),
            .I(N__28349));
    InMux I__4627 (
            .O(N__28349),
            .I(N__28346));
    LocalMux I__4626 (
            .O(N__28346),
            .I(N__28343));
    Odrv4 I__4625 (
            .O(N__28343),
            .I(\SIG_DDS.tmp_buf_8 ));
    InMux I__4624 (
            .O(N__28340),
            .I(N__28336));
    InMux I__4623 (
            .O(N__28339),
            .I(N__28332));
    LocalMux I__4622 (
            .O(N__28336),
            .I(N__28329));
    InMux I__4621 (
            .O(N__28335),
            .I(N__28326));
    LocalMux I__4620 (
            .O(N__28332),
            .I(N__28323));
    Odrv4 I__4619 (
            .O(N__28329),
            .I(buf_dds0_1));
    LocalMux I__4618 (
            .O(N__28326),
            .I(buf_dds0_1));
    Odrv4 I__4617 (
            .O(N__28323),
            .I(buf_dds0_1));
    CascadeMux I__4616 (
            .O(N__28316),
            .I(N__28313));
    InMux I__4615 (
            .O(N__28313),
            .I(N__28310));
    LocalMux I__4614 (
            .O(N__28310),
            .I(\SIG_DDS.tmp_buf_1 ));
    CascadeMux I__4613 (
            .O(N__28307),
            .I(N__28304));
    InMux I__4612 (
            .O(N__28304),
            .I(N__28301));
    LocalMux I__4611 (
            .O(N__28301),
            .I(\SIG_DDS.tmp_buf_2 ));
    InMux I__4610 (
            .O(N__28298),
            .I(N__28295));
    LocalMux I__4609 (
            .O(N__28295),
            .I(N__28292));
    Span4Mux_h I__4608 (
            .O(N__28292),
            .I(N__28289));
    Span4Mux_v I__4607 (
            .O(N__28289),
            .I(N__28284));
    InMux I__4606 (
            .O(N__28288),
            .I(N__28281));
    InMux I__4605 (
            .O(N__28287),
            .I(N__28278));
    Odrv4 I__4604 (
            .O(N__28284),
            .I(buf_dds0_3));
    LocalMux I__4603 (
            .O(N__28281),
            .I(buf_dds0_3));
    LocalMux I__4602 (
            .O(N__28278),
            .I(buf_dds0_3));
    InMux I__4601 (
            .O(N__28271),
            .I(N__28268));
    LocalMux I__4600 (
            .O(N__28268),
            .I(\SIG_DDS.tmp_buf_3 ));
    InMux I__4599 (
            .O(N__28265),
            .I(N__28262));
    LocalMux I__4598 (
            .O(N__28262),
            .I(N__28259));
    Odrv12 I__4597 (
            .O(N__28259),
            .I(n8_adj_1553));
    InMux I__4596 (
            .O(N__28256),
            .I(N__28252));
    InMux I__4595 (
            .O(N__28255),
            .I(N__28249));
    LocalMux I__4594 (
            .O(N__28252),
            .I(N__28246));
    LocalMux I__4593 (
            .O(N__28249),
            .I(n7_adj_1552));
    Odrv12 I__4592 (
            .O(N__28246),
            .I(n7_adj_1552));
    CascadeMux I__4591 (
            .O(N__28241),
            .I(N__28238));
    CascadeBuf I__4590 (
            .O(N__28238),
            .I(N__28235));
    CascadeMux I__4589 (
            .O(N__28235),
            .I(N__28232));
    CascadeBuf I__4588 (
            .O(N__28232),
            .I(N__28229));
    CascadeMux I__4587 (
            .O(N__28229),
            .I(N__28226));
    CascadeBuf I__4586 (
            .O(N__28226),
            .I(N__28223));
    CascadeMux I__4585 (
            .O(N__28223),
            .I(N__28220));
    CascadeBuf I__4584 (
            .O(N__28220),
            .I(N__28217));
    CascadeMux I__4583 (
            .O(N__28217),
            .I(N__28214));
    CascadeBuf I__4582 (
            .O(N__28214),
            .I(N__28211));
    CascadeMux I__4581 (
            .O(N__28211),
            .I(N__28208));
    CascadeBuf I__4580 (
            .O(N__28208),
            .I(N__28205));
    CascadeMux I__4579 (
            .O(N__28205),
            .I(N__28201));
    CascadeMux I__4578 (
            .O(N__28204),
            .I(N__28198));
    CascadeBuf I__4577 (
            .O(N__28201),
            .I(N__28195));
    CascadeBuf I__4576 (
            .O(N__28198),
            .I(N__28192));
    CascadeMux I__4575 (
            .O(N__28195),
            .I(N__28189));
    CascadeMux I__4574 (
            .O(N__28192),
            .I(N__28186));
    CascadeBuf I__4573 (
            .O(N__28189),
            .I(N__28183));
    InMux I__4572 (
            .O(N__28186),
            .I(N__28180));
    CascadeMux I__4571 (
            .O(N__28183),
            .I(N__28177));
    LocalMux I__4570 (
            .O(N__28180),
            .I(N__28174));
    CascadeBuf I__4569 (
            .O(N__28177),
            .I(N__28171));
    Span4Mux_h I__4568 (
            .O(N__28174),
            .I(N__28168));
    CascadeMux I__4567 (
            .O(N__28171),
            .I(N__28165));
    Span4Mux_v I__4566 (
            .O(N__28168),
            .I(N__28162));
    InMux I__4565 (
            .O(N__28165),
            .I(N__28159));
    Sp12to4 I__4564 (
            .O(N__28162),
            .I(N__28156));
    LocalMux I__4563 (
            .O(N__28159),
            .I(N__28153));
    Span12Mux_v I__4562 (
            .O(N__28156),
            .I(N__28148));
    Span12Mux_s8_h I__4561 (
            .O(N__28153),
            .I(N__28148));
    Odrv12 I__4560 (
            .O(N__28148),
            .I(data_index_9_N_216_9));
    InMux I__4559 (
            .O(N__28145),
            .I(N__28140));
    InMux I__4558 (
            .O(N__28144),
            .I(N__28135));
    InMux I__4557 (
            .O(N__28143),
            .I(N__28135));
    LocalMux I__4556 (
            .O(N__28140),
            .I(buf_dds0_10));
    LocalMux I__4555 (
            .O(N__28135),
            .I(buf_dds0_10));
    CascadeMux I__4554 (
            .O(N__28130),
            .I(N__28127));
    InMux I__4553 (
            .O(N__28127),
            .I(N__28124));
    LocalMux I__4552 (
            .O(N__28124),
            .I(\SIG_DDS.tmp_buf_10 ));
    InMux I__4551 (
            .O(N__28121),
            .I(N__28118));
    LocalMux I__4550 (
            .O(N__28118),
            .I(N__28113));
    InMux I__4549 (
            .O(N__28117),
            .I(N__28110));
    InMux I__4548 (
            .O(N__28116),
            .I(N__28107));
    Span4Mux_h I__4547 (
            .O(N__28113),
            .I(N__28102));
    LocalMux I__4546 (
            .O(N__28110),
            .I(N__28102));
    LocalMux I__4545 (
            .O(N__28107),
            .I(buf_dds0_13));
    Odrv4 I__4544 (
            .O(N__28102),
            .I(buf_dds0_13));
    InMux I__4543 (
            .O(N__28097),
            .I(N__28094));
    LocalMux I__4542 (
            .O(N__28094),
            .I(\SIG_DDS.tmp_buf_13 ));
    InMux I__4541 (
            .O(N__28091),
            .I(N__28088));
    LocalMux I__4540 (
            .O(N__28088),
            .I(\SIG_DDS.tmp_buf_11 ));
    CascadeMux I__4539 (
            .O(N__28085),
            .I(N__28082));
    InMux I__4538 (
            .O(N__28082),
            .I(N__28079));
    LocalMux I__4537 (
            .O(N__28079),
            .I(N__28076));
    Odrv12 I__4536 (
            .O(N__28076),
            .I(\SIG_DDS.tmp_buf_12 ));
    CascadeMux I__4535 (
            .O(N__28073),
            .I(N__28070));
    InMux I__4534 (
            .O(N__28070),
            .I(N__28067));
    LocalMux I__4533 (
            .O(N__28067),
            .I(\SIG_DDS.tmp_buf_14 ));
    InMux I__4532 (
            .O(N__28064),
            .I(N__28061));
    LocalMux I__4531 (
            .O(N__28061),
            .I(N__28057));
    InMux I__4530 (
            .O(N__28060),
            .I(N__28053));
    Span4Mux_v I__4529 (
            .O(N__28057),
            .I(N__28050));
    InMux I__4528 (
            .O(N__28056),
            .I(N__28047));
    LocalMux I__4527 (
            .O(N__28053),
            .I(N__28044));
    Span4Mux_v I__4526 (
            .O(N__28050),
            .I(N__28041));
    LocalMux I__4525 (
            .O(N__28047),
            .I(buf_dds0_15));
    Odrv4 I__4524 (
            .O(N__28044),
            .I(buf_dds0_15));
    Odrv4 I__4523 (
            .O(N__28041),
            .I(buf_dds0_15));
    InMux I__4522 (
            .O(N__28034),
            .I(N__28031));
    LocalMux I__4521 (
            .O(N__28031),
            .I(N__28027));
    InMux I__4520 (
            .O(N__28030),
            .I(N__28024));
    Span4Mux_h I__4519 (
            .O(N__28027),
            .I(N__28020));
    LocalMux I__4518 (
            .O(N__28024),
            .I(N__28017));
    InMux I__4517 (
            .O(N__28023),
            .I(N__28014));
    Odrv4 I__4516 (
            .O(N__28020),
            .I(buf_dds0_9));
    Odrv4 I__4515 (
            .O(N__28017),
            .I(buf_dds0_9));
    LocalMux I__4514 (
            .O(N__28014),
            .I(buf_dds0_9));
    CascadeMux I__4513 (
            .O(N__28007),
            .I(N__28004));
    InMux I__4512 (
            .O(N__28004),
            .I(N__28001));
    LocalMux I__4511 (
            .O(N__28001),
            .I(\SIG_DDS.tmp_buf_9 ));
    CascadeMux I__4510 (
            .O(N__27998),
            .I(N__27995));
    InMux I__4509 (
            .O(N__27995),
            .I(N__27992));
    LocalMux I__4508 (
            .O(N__27992),
            .I(\SIG_DDS.tmp_buf_6 ));
    CascadeMux I__4507 (
            .O(N__27989),
            .I(n8_adj_1553_cascade_));
    InMux I__4506 (
            .O(N__27986),
            .I(N__27981));
    InMux I__4505 (
            .O(N__27985),
            .I(N__27976));
    InMux I__4504 (
            .O(N__27984),
            .I(N__27976));
    LocalMux I__4503 (
            .O(N__27981),
            .I(data_index_9));
    LocalMux I__4502 (
            .O(N__27976),
            .I(data_index_9));
    IoInMux I__4501 (
            .O(N__27971),
            .I(N__27968));
    LocalMux I__4500 (
            .O(N__27968),
            .I(N__27965));
    IoSpan4Mux I__4499 (
            .O(N__27965),
            .I(N__27962));
    Span4Mux_s2_h I__4498 (
            .O(N__27962),
            .I(N__27959));
    Span4Mux_h I__4497 (
            .O(N__27959),
            .I(N__27956));
    Sp12to4 I__4496 (
            .O(N__27956),
            .I(N__27953));
    Span12Mux_v I__4495 (
            .O(N__27953),
            .I(N__27950));
    Span12Mux_h I__4494 (
            .O(N__27950),
            .I(N__27947));
    Odrv12 I__4493 (
            .O(N__27947),
            .I(ICE_GPMI_0));
    CEMux I__4492 (
            .O(N__27944),
            .I(N__27941));
    LocalMux I__4491 (
            .O(N__27941),
            .I(N__27938));
    Odrv4 I__4490 (
            .O(N__27938),
            .I(n11401));
    CascadeMux I__4489 (
            .O(N__27935),
            .I(n20772_cascade_));
    CascadeMux I__4488 (
            .O(N__27932),
            .I(n11835_cascade_));
    InMux I__4487 (
            .O(N__27929),
            .I(n19388));
    InMux I__4486 (
            .O(N__27926),
            .I(n19389));
    InMux I__4485 (
            .O(N__27923),
            .I(n19390));
    InMux I__4484 (
            .O(N__27920),
            .I(N__27916));
    InMux I__4483 (
            .O(N__27919),
            .I(N__27913));
    LocalMux I__4482 (
            .O(N__27916),
            .I(N__27907));
    LocalMux I__4481 (
            .O(N__27913),
            .I(N__27907));
    InMux I__4480 (
            .O(N__27912),
            .I(N__27904));
    Odrv4 I__4479 (
            .O(N__27907),
            .I(data_index_8));
    LocalMux I__4478 (
            .O(N__27904),
            .I(data_index_8));
    InMux I__4477 (
            .O(N__27899),
            .I(N__27893));
    InMux I__4476 (
            .O(N__27898),
            .I(N__27893));
    LocalMux I__4475 (
            .O(N__27893),
            .I(n7_adj_1554));
    InMux I__4474 (
            .O(N__27890),
            .I(bfn_10_15_0_));
    InMux I__4473 (
            .O(N__27887),
            .I(n19392));
    InMux I__4472 (
            .O(N__27884),
            .I(N__27880));
    InMux I__4471 (
            .O(N__27883),
            .I(N__27876));
    LocalMux I__4470 (
            .O(N__27880),
            .I(N__27873));
    InMux I__4469 (
            .O(N__27879),
            .I(N__27870));
    LocalMux I__4468 (
            .O(N__27876),
            .I(buf_dds1_2));
    Odrv4 I__4467 (
            .O(N__27873),
            .I(buf_dds1_2));
    LocalMux I__4466 (
            .O(N__27870),
            .I(buf_dds1_2));
    InMux I__4465 (
            .O(N__27863),
            .I(N__27858));
    InMux I__4464 (
            .O(N__27862),
            .I(N__27855));
    InMux I__4463 (
            .O(N__27861),
            .I(N__27852));
    LocalMux I__4462 (
            .O(N__27858),
            .I(data_index_7));
    LocalMux I__4461 (
            .O(N__27855),
            .I(data_index_7));
    LocalMux I__4460 (
            .O(N__27852),
            .I(data_index_7));
    InMux I__4459 (
            .O(N__27845),
            .I(N__27842));
    LocalMux I__4458 (
            .O(N__27842),
            .I(n8_adj_1557));
    CascadeMux I__4457 (
            .O(N__27839),
            .I(n8_adj_1557_cascade_));
    InMux I__4456 (
            .O(N__27836),
            .I(N__27832));
    InMux I__4455 (
            .O(N__27835),
            .I(N__27829));
    LocalMux I__4454 (
            .O(N__27832),
            .I(n7_adj_1556));
    LocalMux I__4453 (
            .O(N__27829),
            .I(n7_adj_1556));
    CascadeMux I__4452 (
            .O(N__27824),
            .I(N__27821));
    CascadeBuf I__4451 (
            .O(N__27821),
            .I(N__27818));
    CascadeMux I__4450 (
            .O(N__27818),
            .I(N__27815));
    CascadeBuf I__4449 (
            .O(N__27815),
            .I(N__27812));
    CascadeMux I__4448 (
            .O(N__27812),
            .I(N__27809));
    CascadeBuf I__4447 (
            .O(N__27809),
            .I(N__27806));
    CascadeMux I__4446 (
            .O(N__27806),
            .I(N__27803));
    CascadeBuf I__4445 (
            .O(N__27803),
            .I(N__27800));
    CascadeMux I__4444 (
            .O(N__27800),
            .I(N__27797));
    CascadeBuf I__4443 (
            .O(N__27797),
            .I(N__27794));
    CascadeMux I__4442 (
            .O(N__27794),
            .I(N__27791));
    CascadeBuf I__4441 (
            .O(N__27791),
            .I(N__27788));
    CascadeMux I__4440 (
            .O(N__27788),
            .I(N__27785));
    CascadeBuf I__4439 (
            .O(N__27785),
            .I(N__27782));
    CascadeMux I__4438 (
            .O(N__27782),
            .I(N__27778));
    CascadeMux I__4437 (
            .O(N__27781),
            .I(N__27775));
    CascadeBuf I__4436 (
            .O(N__27778),
            .I(N__27772));
    CascadeBuf I__4435 (
            .O(N__27775),
            .I(N__27769));
    CascadeMux I__4434 (
            .O(N__27772),
            .I(N__27766));
    CascadeMux I__4433 (
            .O(N__27769),
            .I(N__27763));
    CascadeBuf I__4432 (
            .O(N__27766),
            .I(N__27760));
    InMux I__4431 (
            .O(N__27763),
            .I(N__27757));
    CascadeMux I__4430 (
            .O(N__27760),
            .I(N__27754));
    LocalMux I__4429 (
            .O(N__27757),
            .I(N__27751));
    InMux I__4428 (
            .O(N__27754),
            .I(N__27748));
    Span12Mux_h I__4427 (
            .O(N__27751),
            .I(N__27745));
    LocalMux I__4426 (
            .O(N__27748),
            .I(N__27742));
    Span12Mux_v I__4425 (
            .O(N__27745),
            .I(N__27739));
    Span12Mux_s11_v I__4424 (
            .O(N__27742),
            .I(N__27736));
    Odrv12 I__4423 (
            .O(N__27739),
            .I(data_index_9_N_216_7));
    Odrv12 I__4422 (
            .O(N__27736),
            .I(data_index_9_N_216_7));
    CascadeMux I__4421 (
            .O(N__27731),
            .I(n20663_cascade_));
    InMux I__4420 (
            .O(N__27728),
            .I(bfn_10_14_0_));
    InMux I__4419 (
            .O(N__27725),
            .I(n19384));
    InMux I__4418 (
            .O(N__27722),
            .I(n19385));
    InMux I__4417 (
            .O(N__27719),
            .I(n19386));
    InMux I__4416 (
            .O(N__27716),
            .I(n19387));
    IoInMux I__4415 (
            .O(N__27713),
            .I(N__27710));
    LocalMux I__4414 (
            .O(N__27710),
            .I(N__27707));
    Span4Mux_s2_v I__4413 (
            .O(N__27707),
            .I(N__27704));
    Sp12to4 I__4412 (
            .O(N__27704),
            .I(N__27700));
    InMux I__4411 (
            .O(N__27703),
            .I(N__27697));
    Span12Mux_h I__4410 (
            .O(N__27700),
            .I(N__27694));
    LocalMux I__4409 (
            .O(N__27697),
            .I(N__27690));
    Span12Mux_v I__4408 (
            .O(N__27694),
            .I(N__27687));
    InMux I__4407 (
            .O(N__27693),
            .I(N__27684));
    Span4Mux_h I__4406 (
            .O(N__27690),
            .I(N__27681));
    Odrv12 I__4405 (
            .O(N__27687),
            .I(IAC_OSR1));
    LocalMux I__4404 (
            .O(N__27684),
            .I(IAC_OSR1));
    Odrv4 I__4403 (
            .O(N__27681),
            .I(IAC_OSR1));
    InMux I__4402 (
            .O(N__27674),
            .I(N__27669));
    InMux I__4401 (
            .O(N__27673),
            .I(N__27666));
    InMux I__4400 (
            .O(N__27672),
            .I(N__27663));
    LocalMux I__4399 (
            .O(N__27669),
            .I(comm_cmd_4));
    LocalMux I__4398 (
            .O(N__27666),
            .I(comm_cmd_4));
    LocalMux I__4397 (
            .O(N__27663),
            .I(comm_cmd_4));
    InMux I__4396 (
            .O(N__27656),
            .I(N__27652));
    CascadeMux I__4395 (
            .O(N__27655),
            .I(N__27649));
    LocalMux I__4394 (
            .O(N__27652),
            .I(N__27645));
    InMux I__4393 (
            .O(N__27649),
            .I(N__27642));
    InMux I__4392 (
            .O(N__27648),
            .I(N__27639));
    Span4Mux_h I__4391 (
            .O(N__27645),
            .I(N__27636));
    LocalMux I__4390 (
            .O(N__27642),
            .I(N__27633));
    LocalMux I__4389 (
            .O(N__27639),
            .I(buf_dds1_3));
    Odrv4 I__4388 (
            .O(N__27636),
            .I(buf_dds1_3));
    Odrv12 I__4387 (
            .O(N__27633),
            .I(buf_dds1_3));
    CascadeMux I__4386 (
            .O(N__27626),
            .I(N__27623));
    InMux I__4385 (
            .O(N__27623),
            .I(N__27619));
    CascadeMux I__4384 (
            .O(N__27622),
            .I(N__27616));
    LocalMux I__4383 (
            .O(N__27619),
            .I(N__27612));
    InMux I__4382 (
            .O(N__27616),
            .I(N__27609));
    InMux I__4381 (
            .O(N__27615),
            .I(N__27606));
    Span4Mux_h I__4380 (
            .O(N__27612),
            .I(N__27603));
    LocalMux I__4379 (
            .O(N__27609),
            .I(N__27600));
    LocalMux I__4378 (
            .O(N__27606),
            .I(N__27597));
    Span4Mux_v I__4377 (
            .O(N__27603),
            .I(N__27592));
    Span4Mux_v I__4376 (
            .O(N__27600),
            .I(N__27587));
    Span4Mux_h I__4375 (
            .O(N__27597),
            .I(N__27587));
    InMux I__4374 (
            .O(N__27596),
            .I(N__27584));
    InMux I__4373 (
            .O(N__27595),
            .I(N__27581));
    Odrv4 I__4372 (
            .O(N__27592),
            .I(buf_cfgRTD_1));
    Odrv4 I__4371 (
            .O(N__27587),
            .I(buf_cfgRTD_1));
    LocalMux I__4370 (
            .O(N__27584),
            .I(buf_cfgRTD_1));
    LocalMux I__4369 (
            .O(N__27581),
            .I(buf_cfgRTD_1));
    CascadeMux I__4368 (
            .O(N__27572),
            .I(N__27569));
    InMux I__4367 (
            .O(N__27569),
            .I(N__27566));
    LocalMux I__4366 (
            .O(N__27566),
            .I(N__27563));
    Span4Mux_h I__4365 (
            .O(N__27563),
            .I(N__27559));
    InMux I__4364 (
            .O(N__27562),
            .I(N__27556));
    Odrv4 I__4363 (
            .O(N__27559),
            .I(buf_readRTD_9));
    LocalMux I__4362 (
            .O(N__27556),
            .I(buf_readRTD_9));
    InMux I__4361 (
            .O(N__27551),
            .I(N__27548));
    LocalMux I__4360 (
            .O(N__27548),
            .I(N__27545));
    Span4Mux_h I__4359 (
            .O(N__27545),
            .I(N__27542));
    Odrv4 I__4358 (
            .O(N__27542),
            .I(n9_adj_1416));
    InMux I__4357 (
            .O(N__27539),
            .I(N__27534));
    CascadeMux I__4356 (
            .O(N__27538),
            .I(N__27531));
    CascadeMux I__4355 (
            .O(N__27537),
            .I(N__27528));
    LocalMux I__4354 (
            .O(N__27534),
            .I(N__27525));
    InMux I__4353 (
            .O(N__27531),
            .I(N__27522));
    InMux I__4352 (
            .O(N__27528),
            .I(N__27519));
    Span12Mux_v I__4351 (
            .O(N__27525),
            .I(N__27516));
    LocalMux I__4350 (
            .O(N__27522),
            .I(N__27513));
    LocalMux I__4349 (
            .O(N__27519),
            .I(buf_dds1_0));
    Odrv12 I__4348 (
            .O(N__27516),
            .I(buf_dds1_0));
    Odrv4 I__4347 (
            .O(N__27513),
            .I(buf_dds1_0));
    CascadeMux I__4346 (
            .O(N__27506),
            .I(N__27502));
    CascadeMux I__4345 (
            .O(N__27505),
            .I(N__27498));
    InMux I__4344 (
            .O(N__27502),
            .I(N__27495));
    InMux I__4343 (
            .O(N__27501),
            .I(N__27492));
    InMux I__4342 (
            .O(N__27498),
            .I(N__27489));
    LocalMux I__4341 (
            .O(N__27495),
            .I(N__27484));
    LocalMux I__4340 (
            .O(N__27492),
            .I(N__27484));
    LocalMux I__4339 (
            .O(N__27489),
            .I(N__27480));
    Span4Mux_v I__4338 (
            .O(N__27484),
            .I(N__27477));
    CascadeMux I__4337 (
            .O(N__27483),
            .I(N__27474));
    Span4Mux_h I__4336 (
            .O(N__27480),
            .I(N__27468));
    Span4Mux_h I__4335 (
            .O(N__27477),
            .I(N__27468));
    InMux I__4334 (
            .O(N__27474),
            .I(N__27465));
    InMux I__4333 (
            .O(N__27473),
            .I(N__27462));
    Odrv4 I__4332 (
            .O(N__27468),
            .I(buf_cfgRTD_5));
    LocalMux I__4331 (
            .O(N__27465),
            .I(buf_cfgRTD_5));
    LocalMux I__4330 (
            .O(N__27462),
            .I(buf_cfgRTD_5));
    InMux I__4329 (
            .O(N__27455),
            .I(N__27452));
    LocalMux I__4328 (
            .O(N__27452),
            .I(N__27448));
    InMux I__4327 (
            .O(N__27451),
            .I(N__27444));
    Span4Mux_v I__4326 (
            .O(N__27448),
            .I(N__27441));
    CascadeMux I__4325 (
            .O(N__27447),
            .I(N__27438));
    LocalMux I__4324 (
            .O(N__27444),
            .I(N__27435));
    Sp12to4 I__4323 (
            .O(N__27441),
            .I(N__27432));
    InMux I__4322 (
            .O(N__27438),
            .I(N__27429));
    Span4Mux_h I__4321 (
            .O(N__27435),
            .I(N__27426));
    Span12Mux_h I__4320 (
            .O(N__27432),
            .I(N__27423));
    LocalMux I__4319 (
            .O(N__27429),
            .I(buf_adcdata_iac_18));
    Odrv4 I__4318 (
            .O(N__27426),
            .I(buf_adcdata_iac_18));
    Odrv12 I__4317 (
            .O(N__27423),
            .I(buf_adcdata_iac_18));
    IoInMux I__4316 (
            .O(N__27416),
            .I(N__27413));
    LocalMux I__4315 (
            .O(N__27413),
            .I(N__27410));
    IoSpan4Mux I__4314 (
            .O(N__27410),
            .I(N__27407));
    Span4Mux_s2_v I__4313 (
            .O(N__27407),
            .I(N__27404));
    Sp12to4 I__4312 (
            .O(N__27404),
            .I(N__27400));
    InMux I__4311 (
            .O(N__27403),
            .I(N__27396));
    Span12Mux_v I__4310 (
            .O(N__27400),
            .I(N__27393));
    InMux I__4309 (
            .O(N__27399),
            .I(N__27390));
    LocalMux I__4308 (
            .O(N__27396),
            .I(N__27387));
    Odrv12 I__4307 (
            .O(N__27393),
            .I(IAC_FLT0));
    LocalMux I__4306 (
            .O(N__27390),
            .I(IAC_FLT0));
    Odrv4 I__4305 (
            .O(N__27387),
            .I(IAC_FLT0));
    InMux I__4304 (
            .O(N__27380),
            .I(N__27377));
    LocalMux I__4303 (
            .O(N__27377),
            .I(n20825));
    CascadeMux I__4302 (
            .O(N__27374),
            .I(N__27371));
    CascadeBuf I__4301 (
            .O(N__27371),
            .I(N__27368));
    CascadeMux I__4300 (
            .O(N__27368),
            .I(N__27365));
    CascadeBuf I__4299 (
            .O(N__27365),
            .I(N__27362));
    CascadeMux I__4298 (
            .O(N__27362),
            .I(N__27359));
    CascadeBuf I__4297 (
            .O(N__27359),
            .I(N__27356));
    CascadeMux I__4296 (
            .O(N__27356),
            .I(N__27353));
    CascadeBuf I__4295 (
            .O(N__27353),
            .I(N__27350));
    CascadeMux I__4294 (
            .O(N__27350),
            .I(N__27347));
    CascadeBuf I__4293 (
            .O(N__27347),
            .I(N__27344));
    CascadeMux I__4292 (
            .O(N__27344),
            .I(N__27341));
    CascadeBuf I__4291 (
            .O(N__27341),
            .I(N__27338));
    CascadeMux I__4290 (
            .O(N__27338),
            .I(N__27335));
    CascadeBuf I__4289 (
            .O(N__27335),
            .I(N__27332));
    CascadeMux I__4288 (
            .O(N__27332),
            .I(N__27329));
    CascadeBuf I__4287 (
            .O(N__27329),
            .I(N__27325));
    CascadeMux I__4286 (
            .O(N__27328),
            .I(N__27322));
    CascadeMux I__4285 (
            .O(N__27325),
            .I(N__27319));
    CascadeBuf I__4284 (
            .O(N__27322),
            .I(N__27316));
    CascadeBuf I__4283 (
            .O(N__27319),
            .I(N__27313));
    CascadeMux I__4282 (
            .O(N__27316),
            .I(N__27310));
    CascadeMux I__4281 (
            .O(N__27313),
            .I(N__27307));
    InMux I__4280 (
            .O(N__27310),
            .I(N__27304));
    InMux I__4279 (
            .O(N__27307),
            .I(N__27301));
    LocalMux I__4278 (
            .O(N__27304),
            .I(N__27298));
    LocalMux I__4277 (
            .O(N__27301),
            .I(N__27295));
    Span4Mux_h I__4276 (
            .O(N__27298),
            .I(N__27292));
    Span4Mux_v I__4275 (
            .O(N__27295),
            .I(N__27289));
    Span4Mux_v I__4274 (
            .O(N__27292),
            .I(N__27286));
    Sp12to4 I__4273 (
            .O(N__27289),
            .I(N__27283));
    Span4Mux_h I__4272 (
            .O(N__27286),
            .I(N__27280));
    Span12Mux_h I__4271 (
            .O(N__27283),
            .I(N__27277));
    Odrv4 I__4270 (
            .O(N__27280),
            .I(data_index_9_N_216_0));
    Odrv12 I__4269 (
            .O(N__27277),
            .I(data_index_9_N_216_0));
    InMux I__4268 (
            .O(N__27272),
            .I(N__27265));
    InMux I__4267 (
            .O(N__27271),
            .I(N__27265));
    InMux I__4266 (
            .O(N__27270),
            .I(N__27262));
    LocalMux I__4265 (
            .O(N__27265),
            .I(comm_cmd_5));
    LocalMux I__4264 (
            .O(N__27262),
            .I(comm_cmd_5));
    InMux I__4263 (
            .O(N__27257),
            .I(N__27252));
    InMux I__4262 (
            .O(N__27256),
            .I(N__27249));
    InMux I__4261 (
            .O(N__27255),
            .I(N__27246));
    LocalMux I__4260 (
            .O(N__27252),
            .I(comm_cmd_6));
    LocalMux I__4259 (
            .O(N__27249),
            .I(comm_cmd_6));
    LocalMux I__4258 (
            .O(N__27246),
            .I(comm_cmd_6));
    InMux I__4257 (
            .O(N__27239),
            .I(N__27236));
    LocalMux I__4256 (
            .O(N__27236),
            .I(N__27233));
    Span4Mux_h I__4255 (
            .O(N__27233),
            .I(N__27229));
    InMux I__4254 (
            .O(N__27232),
            .I(N__27226));
    Odrv4 I__4253 (
            .O(N__27229),
            .I(cmd_rdadcbuf_31));
    LocalMux I__4252 (
            .O(N__27226),
            .I(cmd_rdadcbuf_31));
    InMux I__4251 (
            .O(N__27221),
            .I(\ADC_VDC.n19452 ));
    CascadeMux I__4250 (
            .O(N__27218),
            .I(N__27215));
    InMux I__4249 (
            .O(N__27215),
            .I(N__27212));
    LocalMux I__4248 (
            .O(N__27212),
            .I(N__27209));
    Span4Mux_h I__4247 (
            .O(N__27209),
            .I(N__27205));
    InMux I__4246 (
            .O(N__27208),
            .I(N__27202));
    Odrv4 I__4245 (
            .O(N__27205),
            .I(cmd_rdadcbuf_32));
    LocalMux I__4244 (
            .O(N__27202),
            .I(cmd_rdadcbuf_32));
    InMux I__4243 (
            .O(N__27197),
            .I(bfn_10_9_0_));
    InMux I__4242 (
            .O(N__27194),
            .I(\ADC_VDC.n19454 ));
    CEMux I__4241 (
            .O(N__27191),
            .I(N__27187));
    CEMux I__4240 (
            .O(N__27190),
            .I(N__27184));
    LocalMux I__4239 (
            .O(N__27187),
            .I(N__27180));
    LocalMux I__4238 (
            .O(N__27184),
            .I(N__27177));
    CEMux I__4237 (
            .O(N__27183),
            .I(N__27174));
    Span4Mux_v I__4236 (
            .O(N__27180),
            .I(N__27166));
    Span4Mux_v I__4235 (
            .O(N__27177),
            .I(N__27166));
    LocalMux I__4234 (
            .O(N__27174),
            .I(N__27163));
    CEMux I__4233 (
            .O(N__27173),
            .I(N__27160));
    CEMux I__4232 (
            .O(N__27172),
            .I(N__27156));
    CEMux I__4231 (
            .O(N__27171),
            .I(N__27153));
    Span4Mux_h I__4230 (
            .O(N__27166),
            .I(N__27148));
    Span4Mux_v I__4229 (
            .O(N__27163),
            .I(N__27148));
    LocalMux I__4228 (
            .O(N__27160),
            .I(N__27145));
    CEMux I__4227 (
            .O(N__27159),
            .I(N__27142));
    LocalMux I__4226 (
            .O(N__27156),
            .I(N__27139));
    LocalMux I__4225 (
            .O(N__27153),
            .I(N__27136));
    Span4Mux_h I__4224 (
            .O(N__27148),
            .I(N__27133));
    Span4Mux_v I__4223 (
            .O(N__27145),
            .I(N__27130));
    LocalMux I__4222 (
            .O(N__27142),
            .I(N__27127));
    Span4Mux_h I__4221 (
            .O(N__27139),
            .I(N__27124));
    Span4Mux_v I__4220 (
            .O(N__27136),
            .I(N__27117));
    Span4Mux_h I__4219 (
            .O(N__27133),
            .I(N__27117));
    Span4Mux_h I__4218 (
            .O(N__27130),
            .I(N__27117));
    Span4Mux_h I__4217 (
            .O(N__27127),
            .I(N__27114));
    Odrv4 I__4216 (
            .O(N__27124),
            .I(\ADC_VDC.n13038 ));
    Odrv4 I__4215 (
            .O(N__27117),
            .I(\ADC_VDC.n13038 ));
    Odrv4 I__4214 (
            .O(N__27114),
            .I(\ADC_VDC.n13038 ));
    SRMux I__4213 (
            .O(N__27107),
            .I(N__27101));
    SRMux I__4212 (
            .O(N__27106),
            .I(N__27096));
    SRMux I__4211 (
            .O(N__27105),
            .I(N__27092));
    SRMux I__4210 (
            .O(N__27104),
            .I(N__27089));
    LocalMux I__4209 (
            .O(N__27101),
            .I(N__27086));
    SRMux I__4208 (
            .O(N__27100),
            .I(N__27083));
    SRMux I__4207 (
            .O(N__27099),
            .I(N__27080));
    LocalMux I__4206 (
            .O(N__27096),
            .I(N__27077));
    SRMux I__4205 (
            .O(N__27095),
            .I(N__27074));
    LocalMux I__4204 (
            .O(N__27092),
            .I(N__27071));
    LocalMux I__4203 (
            .O(N__27089),
            .I(N__27066));
    Span4Mux_v I__4202 (
            .O(N__27086),
            .I(N__27066));
    LocalMux I__4201 (
            .O(N__27083),
            .I(N__27063));
    LocalMux I__4200 (
            .O(N__27080),
            .I(N__27060));
    Span4Mux_h I__4199 (
            .O(N__27077),
            .I(N__27055));
    LocalMux I__4198 (
            .O(N__27074),
            .I(N__27055));
    Span4Mux_h I__4197 (
            .O(N__27071),
            .I(N__27052));
    Span4Mux_v I__4196 (
            .O(N__27066),
            .I(N__27047));
    Span4Mux_v I__4195 (
            .O(N__27063),
            .I(N__27047));
    Span4Mux_h I__4194 (
            .O(N__27060),
            .I(N__27044));
    Span4Mux_h I__4193 (
            .O(N__27055),
            .I(N__27041));
    Span4Mux_h I__4192 (
            .O(N__27052),
            .I(N__27038));
    Odrv4 I__4191 (
            .O(N__27047),
            .I(\ADC_VDC.n14931 ));
    Odrv4 I__4190 (
            .O(N__27044),
            .I(\ADC_VDC.n14931 ));
    Odrv4 I__4189 (
            .O(N__27041),
            .I(\ADC_VDC.n14931 ));
    Odrv4 I__4188 (
            .O(N__27038),
            .I(\ADC_VDC.n14931 ));
    InMux I__4187 (
            .O(N__27029),
            .I(N__27026));
    LocalMux I__4186 (
            .O(N__27026),
            .I(N__27023));
    Span12Mux_h I__4185 (
            .O(N__27023),
            .I(N__27018));
    InMux I__4184 (
            .O(N__27022),
            .I(N__27015));
    InMux I__4183 (
            .O(N__27021),
            .I(N__27012));
    Odrv12 I__4182 (
            .O(N__27018),
            .I(cmd_rdadcbuf_34));
    LocalMux I__4181 (
            .O(N__27015),
            .I(cmd_rdadcbuf_34));
    LocalMux I__4180 (
            .O(N__27012),
            .I(cmd_rdadcbuf_34));
    InMux I__4179 (
            .O(N__27005),
            .I(\ADC_VDC.n19455 ));
    InMux I__4178 (
            .O(N__27002),
            .I(N__26999));
    LocalMux I__4177 (
            .O(N__26999),
            .I(\ADC_VDC.cmd_rdadcbuf_35_N_1139_34 ));
    CascadeMux I__4176 (
            .O(N__26996),
            .I(N__26993));
    InMux I__4175 (
            .O(N__26993),
            .I(N__26990));
    LocalMux I__4174 (
            .O(N__26990),
            .I(N__26987));
    Span4Mux_h I__4173 (
            .O(N__26987),
            .I(N__26984));
    Span4Mux_v I__4172 (
            .O(N__26984),
            .I(N__26981));
    Odrv4 I__4171 (
            .O(N__26981),
            .I(n20824));
    InMux I__4170 (
            .O(N__26978),
            .I(N__26975));
    LocalMux I__4169 (
            .O(N__26975),
            .I(n22118));
    InMux I__4168 (
            .O(N__26972),
            .I(N__26967));
    CascadeMux I__4167 (
            .O(N__26971),
            .I(N__26964));
    InMux I__4166 (
            .O(N__26970),
            .I(N__26961));
    LocalMux I__4165 (
            .O(N__26967),
            .I(N__26958));
    InMux I__4164 (
            .O(N__26964),
            .I(N__26955));
    LocalMux I__4163 (
            .O(N__26961),
            .I(cmd_rdadctmp_8));
    Odrv12 I__4162 (
            .O(N__26958),
            .I(cmd_rdadctmp_8));
    LocalMux I__4161 (
            .O(N__26955),
            .I(cmd_rdadctmp_8));
    InMux I__4160 (
            .O(N__26948),
            .I(N__26944));
    InMux I__4159 (
            .O(N__26947),
            .I(N__26941));
    LocalMux I__4158 (
            .O(N__26944),
            .I(cmd_rdadcbuf_22));
    LocalMux I__4157 (
            .O(N__26941),
            .I(cmd_rdadcbuf_22));
    InMux I__4156 (
            .O(N__26936),
            .I(\ADC_VDC.n19443 ));
    InMux I__4155 (
            .O(N__26933),
            .I(N__26930));
    LocalMux I__4154 (
            .O(N__26930),
            .I(N__26926));
    InMux I__4153 (
            .O(N__26929),
            .I(N__26923));
    Odrv4 I__4152 (
            .O(N__26926),
            .I(cmd_rdadcbuf_23));
    LocalMux I__4151 (
            .O(N__26923),
            .I(cmd_rdadcbuf_23));
    InMux I__4150 (
            .O(N__26918),
            .I(\ADC_VDC.n19444 ));
    InMux I__4149 (
            .O(N__26915),
            .I(bfn_10_8_0_));
    InMux I__4148 (
            .O(N__26912),
            .I(\ADC_VDC.n19446 ));
    InMux I__4147 (
            .O(N__26909),
            .I(\ADC_VDC.n19447 ));
    InMux I__4146 (
            .O(N__26906),
            .I(\ADC_VDC.n19448 ));
    CascadeMux I__4145 (
            .O(N__26903),
            .I(N__26900));
    InMux I__4144 (
            .O(N__26900),
            .I(N__26897));
    LocalMux I__4143 (
            .O(N__26897),
            .I(N__26894));
    Span4Mux_h I__4142 (
            .O(N__26894),
            .I(N__26890));
    InMux I__4141 (
            .O(N__26893),
            .I(N__26887));
    Odrv4 I__4140 (
            .O(N__26890),
            .I(cmd_rdadcbuf_28));
    LocalMux I__4139 (
            .O(N__26887),
            .I(cmd_rdadcbuf_28));
    InMux I__4138 (
            .O(N__26882),
            .I(\ADC_VDC.n19449 ));
    InMux I__4137 (
            .O(N__26879),
            .I(N__26876));
    LocalMux I__4136 (
            .O(N__26876),
            .I(N__26872));
    InMux I__4135 (
            .O(N__26875),
            .I(N__26869));
    Odrv4 I__4134 (
            .O(N__26872),
            .I(cmd_rdadcbuf_29));
    LocalMux I__4133 (
            .O(N__26869),
            .I(cmd_rdadcbuf_29));
    InMux I__4132 (
            .O(N__26864),
            .I(\ADC_VDC.n19450 ));
    InMux I__4131 (
            .O(N__26861),
            .I(N__26858));
    LocalMux I__4130 (
            .O(N__26858),
            .I(N__26854));
    InMux I__4129 (
            .O(N__26857),
            .I(N__26851));
    Odrv12 I__4128 (
            .O(N__26854),
            .I(cmd_rdadcbuf_30));
    LocalMux I__4127 (
            .O(N__26851),
            .I(cmd_rdadcbuf_30));
    InMux I__4126 (
            .O(N__26846),
            .I(\ADC_VDC.n19451 ));
    InMux I__4125 (
            .O(N__26843),
            .I(N__26838));
    InMux I__4124 (
            .O(N__26842),
            .I(N__26835));
    InMux I__4123 (
            .O(N__26841),
            .I(N__26832));
    LocalMux I__4122 (
            .O(N__26838),
            .I(cmd_rdadctmp_14_adj_1465));
    LocalMux I__4121 (
            .O(N__26835),
            .I(cmd_rdadctmp_14_adj_1465));
    LocalMux I__4120 (
            .O(N__26832),
            .I(cmd_rdadctmp_14_adj_1465));
    InMux I__4119 (
            .O(N__26825),
            .I(N__26821));
    CascadeMux I__4118 (
            .O(N__26824),
            .I(N__26818));
    LocalMux I__4117 (
            .O(N__26821),
            .I(N__26815));
    InMux I__4116 (
            .O(N__26818),
            .I(N__26812));
    Odrv12 I__4115 (
            .O(N__26815),
            .I(cmd_rdadcbuf_14));
    LocalMux I__4114 (
            .O(N__26812),
            .I(cmd_rdadcbuf_14));
    InMux I__4113 (
            .O(N__26807),
            .I(\ADC_VDC.n19435 ));
    CascadeMux I__4112 (
            .O(N__26804),
            .I(N__26799));
    InMux I__4111 (
            .O(N__26803),
            .I(N__26794));
    InMux I__4110 (
            .O(N__26802),
            .I(N__26794));
    InMux I__4109 (
            .O(N__26799),
            .I(N__26791));
    LocalMux I__4108 (
            .O(N__26794),
            .I(cmd_rdadctmp_15_adj_1464));
    LocalMux I__4107 (
            .O(N__26791),
            .I(cmd_rdadctmp_15_adj_1464));
    InMux I__4106 (
            .O(N__26786),
            .I(N__26783));
    LocalMux I__4105 (
            .O(N__26783),
            .I(N__26779));
    InMux I__4104 (
            .O(N__26782),
            .I(N__26776));
    Odrv4 I__4103 (
            .O(N__26779),
            .I(cmd_rdadcbuf_15));
    LocalMux I__4102 (
            .O(N__26776),
            .I(cmd_rdadcbuf_15));
    InMux I__4101 (
            .O(N__26771),
            .I(\ADC_VDC.n19436 ));
    CascadeMux I__4100 (
            .O(N__26768),
            .I(N__26763));
    CascadeMux I__4099 (
            .O(N__26767),
            .I(N__26760));
    CascadeMux I__4098 (
            .O(N__26766),
            .I(N__26757));
    InMux I__4097 (
            .O(N__26763),
            .I(N__26752));
    InMux I__4096 (
            .O(N__26760),
            .I(N__26752));
    InMux I__4095 (
            .O(N__26757),
            .I(N__26749));
    LocalMux I__4094 (
            .O(N__26752),
            .I(cmd_rdadctmp_16_adj_1463));
    LocalMux I__4093 (
            .O(N__26749),
            .I(cmd_rdadctmp_16_adj_1463));
    InMux I__4092 (
            .O(N__26744),
            .I(N__26741));
    LocalMux I__4091 (
            .O(N__26741),
            .I(N__26738));
    Span4Mux_v I__4090 (
            .O(N__26738),
            .I(N__26734));
    InMux I__4089 (
            .O(N__26737),
            .I(N__26731));
    Odrv4 I__4088 (
            .O(N__26734),
            .I(cmd_rdadcbuf_16));
    LocalMux I__4087 (
            .O(N__26731),
            .I(cmd_rdadcbuf_16));
    InMux I__4086 (
            .O(N__26726),
            .I(bfn_10_7_0_));
    CascadeMux I__4085 (
            .O(N__26723),
            .I(N__26718));
    InMux I__4084 (
            .O(N__26722),
            .I(N__26713));
    InMux I__4083 (
            .O(N__26721),
            .I(N__26713));
    InMux I__4082 (
            .O(N__26718),
            .I(N__26710));
    LocalMux I__4081 (
            .O(N__26713),
            .I(cmd_rdadctmp_17_adj_1462));
    LocalMux I__4080 (
            .O(N__26710),
            .I(cmd_rdadctmp_17_adj_1462));
    CascadeMux I__4079 (
            .O(N__26705),
            .I(N__26702));
    InMux I__4078 (
            .O(N__26702),
            .I(N__26699));
    LocalMux I__4077 (
            .O(N__26699),
            .I(N__26696));
    Span4Mux_v I__4076 (
            .O(N__26696),
            .I(N__26692));
    InMux I__4075 (
            .O(N__26695),
            .I(N__26689));
    Odrv4 I__4074 (
            .O(N__26692),
            .I(cmd_rdadcbuf_17));
    LocalMux I__4073 (
            .O(N__26689),
            .I(cmd_rdadcbuf_17));
    InMux I__4072 (
            .O(N__26684),
            .I(\ADC_VDC.n19438 ));
    CascadeMux I__4071 (
            .O(N__26681),
            .I(N__26676));
    InMux I__4070 (
            .O(N__26680),
            .I(N__26673));
    InMux I__4069 (
            .O(N__26679),
            .I(N__26670));
    InMux I__4068 (
            .O(N__26676),
            .I(N__26667));
    LocalMux I__4067 (
            .O(N__26673),
            .I(cmd_rdadctmp_18_adj_1461));
    LocalMux I__4066 (
            .O(N__26670),
            .I(cmd_rdadctmp_18_adj_1461));
    LocalMux I__4065 (
            .O(N__26667),
            .I(cmd_rdadctmp_18_adj_1461));
    InMux I__4064 (
            .O(N__26660),
            .I(N__26657));
    LocalMux I__4063 (
            .O(N__26657),
            .I(N__26654));
    Span4Mux_h I__4062 (
            .O(N__26654),
            .I(N__26650));
    InMux I__4061 (
            .O(N__26653),
            .I(N__26647));
    Odrv4 I__4060 (
            .O(N__26650),
            .I(cmd_rdadcbuf_18));
    LocalMux I__4059 (
            .O(N__26647),
            .I(cmd_rdadcbuf_18));
    InMux I__4058 (
            .O(N__26642),
            .I(\ADC_VDC.n19439 ));
    CascadeMux I__4057 (
            .O(N__26639),
            .I(N__26634));
    InMux I__4056 (
            .O(N__26638),
            .I(N__26629));
    InMux I__4055 (
            .O(N__26637),
            .I(N__26629));
    InMux I__4054 (
            .O(N__26634),
            .I(N__26626));
    LocalMux I__4053 (
            .O(N__26629),
            .I(cmd_rdadctmp_19_adj_1460));
    LocalMux I__4052 (
            .O(N__26626),
            .I(cmd_rdadctmp_19_adj_1460));
    InMux I__4051 (
            .O(N__26621),
            .I(N__26618));
    LocalMux I__4050 (
            .O(N__26618),
            .I(N__26614));
    InMux I__4049 (
            .O(N__26617),
            .I(N__26611));
    Odrv12 I__4048 (
            .O(N__26614),
            .I(cmd_rdadcbuf_19));
    LocalMux I__4047 (
            .O(N__26611),
            .I(cmd_rdadcbuf_19));
    InMux I__4046 (
            .O(N__26606),
            .I(\ADC_VDC.n19440 ));
    CascadeMux I__4045 (
            .O(N__26603),
            .I(N__26598));
    InMux I__4044 (
            .O(N__26602),
            .I(N__26595));
    CascadeMux I__4043 (
            .O(N__26601),
            .I(N__26592));
    InMux I__4042 (
            .O(N__26598),
            .I(N__26589));
    LocalMux I__4041 (
            .O(N__26595),
            .I(N__26586));
    InMux I__4040 (
            .O(N__26592),
            .I(N__26583));
    LocalMux I__4039 (
            .O(N__26589),
            .I(cmd_rdadctmp_20_adj_1459));
    Odrv4 I__4038 (
            .O(N__26586),
            .I(cmd_rdadctmp_20_adj_1459));
    LocalMux I__4037 (
            .O(N__26583),
            .I(cmd_rdadctmp_20_adj_1459));
    InMux I__4036 (
            .O(N__26576),
            .I(\ADC_VDC.n19441 ));
    CascadeMux I__4035 (
            .O(N__26573),
            .I(N__26570));
    InMux I__4034 (
            .O(N__26570),
            .I(N__26565));
    InMux I__4033 (
            .O(N__26569),
            .I(N__26560));
    InMux I__4032 (
            .O(N__26568),
            .I(N__26560));
    LocalMux I__4031 (
            .O(N__26565),
            .I(N__26557));
    LocalMux I__4030 (
            .O(N__26560),
            .I(cmd_rdadctmp_21_adj_1458));
    Odrv4 I__4029 (
            .O(N__26557),
            .I(cmd_rdadctmp_21_adj_1458));
    CascadeMux I__4028 (
            .O(N__26552),
            .I(N__26549));
    InMux I__4027 (
            .O(N__26549),
            .I(N__26546));
    LocalMux I__4026 (
            .O(N__26546),
            .I(N__26543));
    Span4Mux_h I__4025 (
            .O(N__26543),
            .I(N__26539));
    InMux I__4024 (
            .O(N__26542),
            .I(N__26536));
    Odrv4 I__4023 (
            .O(N__26539),
            .I(cmd_rdadcbuf_21));
    LocalMux I__4022 (
            .O(N__26536),
            .I(cmd_rdadcbuf_21));
    InMux I__4021 (
            .O(N__26531),
            .I(\ADC_VDC.n19442 ));
    InMux I__4020 (
            .O(N__26528),
            .I(\ADC_VDC.n19427 ));
    InMux I__4019 (
            .O(N__26525),
            .I(N__26521));
    CascadeMux I__4018 (
            .O(N__26524),
            .I(N__26517));
    LocalMux I__4017 (
            .O(N__26521),
            .I(N__26514));
    InMux I__4016 (
            .O(N__26520),
            .I(N__26511));
    InMux I__4015 (
            .O(N__26517),
            .I(N__26508));
    Odrv4 I__4014 (
            .O(N__26514),
            .I(cmd_rdadctmp_7_adj_1472));
    LocalMux I__4013 (
            .O(N__26511),
            .I(cmd_rdadctmp_7_adj_1472));
    LocalMux I__4012 (
            .O(N__26508),
            .I(cmd_rdadctmp_7_adj_1472));
    InMux I__4011 (
            .O(N__26501),
            .I(N__26498));
    LocalMux I__4010 (
            .O(N__26498),
            .I(\ADC_VDC.cmd_rdadcbuf_7 ));
    InMux I__4009 (
            .O(N__26495),
            .I(\ADC_VDC.n19428 ));
    InMux I__4008 (
            .O(N__26492),
            .I(N__26488));
    CascadeMux I__4007 (
            .O(N__26491),
            .I(N__26484));
    LocalMux I__4006 (
            .O(N__26488),
            .I(N__26481));
    InMux I__4005 (
            .O(N__26487),
            .I(N__26478));
    InMux I__4004 (
            .O(N__26484),
            .I(N__26475));
    Odrv4 I__4003 (
            .O(N__26481),
            .I(cmd_rdadctmp_8_adj_1471));
    LocalMux I__4002 (
            .O(N__26478),
            .I(cmd_rdadctmp_8_adj_1471));
    LocalMux I__4001 (
            .O(N__26475),
            .I(cmd_rdadctmp_8_adj_1471));
    InMux I__4000 (
            .O(N__26468),
            .I(N__26465));
    LocalMux I__3999 (
            .O(N__26465),
            .I(\ADC_VDC.cmd_rdadcbuf_8 ));
    InMux I__3998 (
            .O(N__26462),
            .I(bfn_10_6_0_));
    CascadeMux I__3997 (
            .O(N__26459),
            .I(N__26455));
    CascadeMux I__3996 (
            .O(N__26458),
            .I(N__26451));
    InMux I__3995 (
            .O(N__26455),
            .I(N__26448));
    InMux I__3994 (
            .O(N__26454),
            .I(N__26445));
    InMux I__3993 (
            .O(N__26451),
            .I(N__26442));
    LocalMux I__3992 (
            .O(N__26448),
            .I(cmd_rdadctmp_9_adj_1470));
    LocalMux I__3991 (
            .O(N__26445),
            .I(cmd_rdadctmp_9_adj_1470));
    LocalMux I__3990 (
            .O(N__26442),
            .I(cmd_rdadctmp_9_adj_1470));
    InMux I__3989 (
            .O(N__26435),
            .I(N__26432));
    LocalMux I__3988 (
            .O(N__26432),
            .I(\ADC_VDC.cmd_rdadcbuf_9 ));
    InMux I__3987 (
            .O(N__26429),
            .I(\ADC_VDC.n19430 ));
    CascadeMux I__3986 (
            .O(N__26426),
            .I(N__26422));
    CascadeMux I__3985 (
            .O(N__26425),
            .I(N__26418));
    InMux I__3984 (
            .O(N__26422),
            .I(N__26415));
    InMux I__3983 (
            .O(N__26421),
            .I(N__26412));
    InMux I__3982 (
            .O(N__26418),
            .I(N__26409));
    LocalMux I__3981 (
            .O(N__26415),
            .I(cmd_rdadctmp_10_adj_1469));
    LocalMux I__3980 (
            .O(N__26412),
            .I(cmd_rdadctmp_10_adj_1469));
    LocalMux I__3979 (
            .O(N__26409),
            .I(cmd_rdadctmp_10_adj_1469));
    InMux I__3978 (
            .O(N__26402),
            .I(N__26399));
    LocalMux I__3977 (
            .O(N__26399),
            .I(\ADC_VDC.cmd_rdadcbuf_10 ));
    InMux I__3976 (
            .O(N__26396),
            .I(\ADC_VDC.n19431 ));
    CascadeMux I__3975 (
            .O(N__26393),
            .I(N__26388));
    InMux I__3974 (
            .O(N__26392),
            .I(N__26383));
    InMux I__3973 (
            .O(N__26391),
            .I(N__26383));
    InMux I__3972 (
            .O(N__26388),
            .I(N__26380));
    LocalMux I__3971 (
            .O(N__26383),
            .I(cmd_rdadctmp_11_adj_1468));
    LocalMux I__3970 (
            .O(N__26380),
            .I(cmd_rdadctmp_11_adj_1468));
    InMux I__3969 (
            .O(N__26375),
            .I(\ADC_VDC.n19432 ));
    CascadeMux I__3968 (
            .O(N__26372),
            .I(N__26368));
    CascadeMux I__3967 (
            .O(N__26371),
            .I(N__26365));
    InMux I__3966 (
            .O(N__26368),
            .I(N__26361));
    InMux I__3965 (
            .O(N__26365),
            .I(N__26356));
    InMux I__3964 (
            .O(N__26364),
            .I(N__26356));
    LocalMux I__3963 (
            .O(N__26361),
            .I(N__26353));
    LocalMux I__3962 (
            .O(N__26356),
            .I(cmd_rdadctmp_12_adj_1467));
    Odrv4 I__3961 (
            .O(N__26353),
            .I(cmd_rdadctmp_12_adj_1467));
    InMux I__3960 (
            .O(N__26348),
            .I(N__26345));
    LocalMux I__3959 (
            .O(N__26345),
            .I(N__26341));
    InMux I__3958 (
            .O(N__26344),
            .I(N__26338));
    Odrv12 I__3957 (
            .O(N__26341),
            .I(cmd_rdadcbuf_12));
    LocalMux I__3956 (
            .O(N__26338),
            .I(cmd_rdadcbuf_12));
    InMux I__3955 (
            .O(N__26333),
            .I(\ADC_VDC.n19433 ));
    InMux I__3954 (
            .O(N__26330),
            .I(N__26323));
    InMux I__3953 (
            .O(N__26329),
            .I(N__26323));
    InMux I__3952 (
            .O(N__26328),
            .I(N__26320));
    LocalMux I__3951 (
            .O(N__26323),
            .I(cmd_rdadctmp_13_adj_1466));
    LocalMux I__3950 (
            .O(N__26320),
            .I(cmd_rdadctmp_13_adj_1466));
    InMux I__3949 (
            .O(N__26315),
            .I(N__26312));
    LocalMux I__3948 (
            .O(N__26312),
            .I(N__26308));
    CascadeMux I__3947 (
            .O(N__26311),
            .I(N__26305));
    Span4Mux_h I__3946 (
            .O(N__26308),
            .I(N__26302));
    InMux I__3945 (
            .O(N__26305),
            .I(N__26299));
    Odrv4 I__3944 (
            .O(N__26302),
            .I(cmd_rdadcbuf_13));
    LocalMux I__3943 (
            .O(N__26299),
            .I(cmd_rdadcbuf_13));
    InMux I__3942 (
            .O(N__26294),
            .I(\ADC_VDC.n19434 ));
    CascadeMux I__3941 (
            .O(N__26291),
            .I(N__26285));
    CascadeMux I__3940 (
            .O(N__26290),
            .I(N__26281));
    InMux I__3939 (
            .O(N__26289),
            .I(N__26262));
    InMux I__3938 (
            .O(N__26288),
            .I(N__26262));
    InMux I__3937 (
            .O(N__26285),
            .I(N__26262));
    InMux I__3936 (
            .O(N__26284),
            .I(N__26262));
    InMux I__3935 (
            .O(N__26281),
            .I(N__26262));
    CascadeMux I__3934 (
            .O(N__26280),
            .I(N__26259));
    CascadeMux I__3933 (
            .O(N__26279),
            .I(N__26256));
    CascadeMux I__3932 (
            .O(N__26278),
            .I(N__26251));
    CascadeMux I__3931 (
            .O(N__26277),
            .I(N__26247));
    CascadeMux I__3930 (
            .O(N__26276),
            .I(N__26243));
    CascadeMux I__3929 (
            .O(N__26275),
            .I(N__26237));
    CascadeMux I__3928 (
            .O(N__26274),
            .I(N__26233));
    CascadeMux I__3927 (
            .O(N__26273),
            .I(N__26229));
    LocalMux I__3926 (
            .O(N__26262),
            .I(N__26226));
    InMux I__3925 (
            .O(N__26259),
            .I(N__26215));
    InMux I__3924 (
            .O(N__26256),
            .I(N__26215));
    InMux I__3923 (
            .O(N__26255),
            .I(N__26215));
    InMux I__3922 (
            .O(N__26254),
            .I(N__26215));
    InMux I__3921 (
            .O(N__26251),
            .I(N__26215));
    InMux I__3920 (
            .O(N__26250),
            .I(N__26202));
    InMux I__3919 (
            .O(N__26247),
            .I(N__26202));
    InMux I__3918 (
            .O(N__26246),
            .I(N__26202));
    InMux I__3917 (
            .O(N__26243),
            .I(N__26202));
    InMux I__3916 (
            .O(N__26242),
            .I(N__26202));
    InMux I__3915 (
            .O(N__26241),
            .I(N__26202));
    InMux I__3914 (
            .O(N__26240),
            .I(N__26189));
    InMux I__3913 (
            .O(N__26237),
            .I(N__26189));
    InMux I__3912 (
            .O(N__26236),
            .I(N__26189));
    InMux I__3911 (
            .O(N__26233),
            .I(N__26189));
    InMux I__3910 (
            .O(N__26232),
            .I(N__26189));
    InMux I__3909 (
            .O(N__26229),
            .I(N__26189));
    Odrv4 I__3908 (
            .O(N__26226),
            .I(n12875));
    LocalMux I__3907 (
            .O(N__26215),
            .I(n12875));
    LocalMux I__3906 (
            .O(N__26202),
            .I(n12875));
    LocalMux I__3905 (
            .O(N__26189),
            .I(n12875));
    CascadeMux I__3904 (
            .O(N__26180),
            .I(N__26176));
    CascadeMux I__3903 (
            .O(N__26179),
            .I(N__26172));
    InMux I__3902 (
            .O(N__26176),
            .I(N__26167));
    InMux I__3901 (
            .O(N__26175),
            .I(N__26167));
    InMux I__3900 (
            .O(N__26172),
            .I(N__26164));
    LocalMux I__3899 (
            .O(N__26167),
            .I(cmd_rdadctmp_0_adj_1479));
    LocalMux I__3898 (
            .O(N__26164),
            .I(cmd_rdadctmp_0_adj_1479));
    InMux I__3897 (
            .O(N__26159),
            .I(N__26156));
    LocalMux I__3896 (
            .O(N__26156),
            .I(\ADC_VDC.cmd_rdadcbuf_0 ));
    CascadeMux I__3895 (
            .O(N__26153),
            .I(N__26148));
    InMux I__3894 (
            .O(N__26152),
            .I(N__26145));
    InMux I__3893 (
            .O(N__26151),
            .I(N__26142));
    InMux I__3892 (
            .O(N__26148),
            .I(N__26139));
    LocalMux I__3891 (
            .O(N__26145),
            .I(cmd_rdadctmp_1_adj_1478));
    LocalMux I__3890 (
            .O(N__26142),
            .I(cmd_rdadctmp_1_adj_1478));
    LocalMux I__3889 (
            .O(N__26139),
            .I(cmd_rdadctmp_1_adj_1478));
    InMux I__3888 (
            .O(N__26132),
            .I(N__26129));
    LocalMux I__3887 (
            .O(N__26129),
            .I(\ADC_VDC.cmd_rdadcbuf_1 ));
    InMux I__3886 (
            .O(N__26126),
            .I(\ADC_VDC.n19422 ));
    CascadeMux I__3885 (
            .O(N__26123),
            .I(N__26118));
    InMux I__3884 (
            .O(N__26122),
            .I(N__26113));
    InMux I__3883 (
            .O(N__26121),
            .I(N__26113));
    InMux I__3882 (
            .O(N__26118),
            .I(N__26110));
    LocalMux I__3881 (
            .O(N__26113),
            .I(cmd_rdadctmp_2_adj_1477));
    LocalMux I__3880 (
            .O(N__26110),
            .I(cmd_rdadctmp_2_adj_1477));
    InMux I__3879 (
            .O(N__26105),
            .I(N__26102));
    LocalMux I__3878 (
            .O(N__26102),
            .I(\ADC_VDC.cmd_rdadcbuf_2 ));
    InMux I__3877 (
            .O(N__26099),
            .I(\ADC_VDC.n19423 ));
    CascadeMux I__3876 (
            .O(N__26096),
            .I(N__26092));
    CascadeMux I__3875 (
            .O(N__26095),
            .I(N__26088));
    InMux I__3874 (
            .O(N__26092),
            .I(N__26083));
    InMux I__3873 (
            .O(N__26091),
            .I(N__26083));
    InMux I__3872 (
            .O(N__26088),
            .I(N__26080));
    LocalMux I__3871 (
            .O(N__26083),
            .I(cmd_rdadctmp_3_adj_1476));
    LocalMux I__3870 (
            .O(N__26080),
            .I(cmd_rdadctmp_3_adj_1476));
    InMux I__3869 (
            .O(N__26075),
            .I(N__26072));
    LocalMux I__3868 (
            .O(N__26072),
            .I(\ADC_VDC.cmd_rdadcbuf_3 ));
    InMux I__3867 (
            .O(N__26069),
            .I(\ADC_VDC.n19424 ));
    CascadeMux I__3866 (
            .O(N__26066),
            .I(N__26061));
    InMux I__3865 (
            .O(N__26065),
            .I(N__26058));
    InMux I__3864 (
            .O(N__26064),
            .I(N__26055));
    InMux I__3863 (
            .O(N__26061),
            .I(N__26052));
    LocalMux I__3862 (
            .O(N__26058),
            .I(cmd_rdadctmp_4_adj_1475));
    LocalMux I__3861 (
            .O(N__26055),
            .I(cmd_rdadctmp_4_adj_1475));
    LocalMux I__3860 (
            .O(N__26052),
            .I(cmd_rdadctmp_4_adj_1475));
    InMux I__3859 (
            .O(N__26045),
            .I(N__26042));
    LocalMux I__3858 (
            .O(N__26042),
            .I(\ADC_VDC.cmd_rdadcbuf_4 ));
    InMux I__3857 (
            .O(N__26039),
            .I(\ADC_VDC.n19425 ));
    CascadeMux I__3856 (
            .O(N__26036),
            .I(N__26032));
    CascadeMux I__3855 (
            .O(N__26035),
            .I(N__26028));
    InMux I__3854 (
            .O(N__26032),
            .I(N__26025));
    InMux I__3853 (
            .O(N__26031),
            .I(N__26022));
    InMux I__3852 (
            .O(N__26028),
            .I(N__26019));
    LocalMux I__3851 (
            .O(N__26025),
            .I(cmd_rdadctmp_5_adj_1474));
    LocalMux I__3850 (
            .O(N__26022),
            .I(cmd_rdadctmp_5_adj_1474));
    LocalMux I__3849 (
            .O(N__26019),
            .I(cmd_rdadctmp_5_adj_1474));
    InMux I__3848 (
            .O(N__26012),
            .I(N__26009));
    LocalMux I__3847 (
            .O(N__26009),
            .I(\ADC_VDC.cmd_rdadcbuf_5 ));
    InMux I__3846 (
            .O(N__26006),
            .I(\ADC_VDC.n19426 ));
    CascadeMux I__3845 (
            .O(N__26003),
            .I(N__25998));
    InMux I__3844 (
            .O(N__26002),
            .I(N__25993));
    InMux I__3843 (
            .O(N__26001),
            .I(N__25993));
    InMux I__3842 (
            .O(N__25998),
            .I(N__25990));
    LocalMux I__3841 (
            .O(N__25993),
            .I(cmd_rdadctmp_6_adj_1473));
    LocalMux I__3840 (
            .O(N__25990),
            .I(cmd_rdadctmp_6_adj_1473));
    InMux I__3839 (
            .O(N__25985),
            .I(N__25982));
    LocalMux I__3838 (
            .O(N__25982),
            .I(\ADC_VDC.cmd_rdadcbuf_6 ));
    CascadeMux I__3837 (
            .O(N__25979),
            .I(N__25976));
    InMux I__3836 (
            .O(N__25976),
            .I(N__25973));
    LocalMux I__3835 (
            .O(N__25973),
            .I(N__25969));
    InMux I__3834 (
            .O(N__25972),
            .I(N__25965));
    Span4Mux_h I__3833 (
            .O(N__25969),
            .I(N__25962));
    InMux I__3832 (
            .O(N__25968),
            .I(N__25959));
    LocalMux I__3831 (
            .O(N__25965),
            .I(cmd_rdadctmp_12));
    Odrv4 I__3830 (
            .O(N__25962),
            .I(cmd_rdadctmp_12));
    LocalMux I__3829 (
            .O(N__25959),
            .I(cmd_rdadctmp_12));
    CascadeMux I__3828 (
            .O(N__25952),
            .I(N__25949));
    InMux I__3827 (
            .O(N__25949),
            .I(N__25945));
    CascadeMux I__3826 (
            .O(N__25948),
            .I(N__25941));
    LocalMux I__3825 (
            .O(N__25945),
            .I(N__25938));
    InMux I__3824 (
            .O(N__25944),
            .I(N__25935));
    InMux I__3823 (
            .O(N__25941),
            .I(N__25932));
    Span4Mux_h I__3822 (
            .O(N__25938),
            .I(N__25927));
    LocalMux I__3821 (
            .O(N__25935),
            .I(N__25927));
    LocalMux I__3820 (
            .O(N__25932),
            .I(cmd_rdadctmp_13));
    Odrv4 I__3819 (
            .O(N__25927),
            .I(cmd_rdadctmp_13));
    InMux I__3818 (
            .O(N__25922),
            .I(N__25918));
    CascadeMux I__3817 (
            .O(N__25921),
            .I(N__25915));
    LocalMux I__3816 (
            .O(N__25918),
            .I(N__25912));
    InMux I__3815 (
            .O(N__25915),
            .I(N__25909));
    Span4Mux_h I__3814 (
            .O(N__25912),
            .I(N__25906));
    LocalMux I__3813 (
            .O(N__25909),
            .I(cmd_rdadctmp_6));
    Odrv4 I__3812 (
            .O(N__25906),
            .I(cmd_rdadctmp_6));
    InMux I__3811 (
            .O(N__25901),
            .I(N__25897));
    InMux I__3810 (
            .O(N__25900),
            .I(N__25894));
    LocalMux I__3809 (
            .O(N__25897),
            .I(cmd_rdadctmp_7));
    LocalMux I__3808 (
            .O(N__25894),
            .I(cmd_rdadctmp_7));
    CascadeMux I__3807 (
            .O(N__25889),
            .I(N__25886));
    InMux I__3806 (
            .O(N__25886),
            .I(N__25882));
    CascadeMux I__3805 (
            .O(N__25885),
            .I(N__25879));
    LocalMux I__3804 (
            .O(N__25882),
            .I(N__25875));
    InMux I__3803 (
            .O(N__25879),
            .I(N__25870));
    InMux I__3802 (
            .O(N__25878),
            .I(N__25870));
    Odrv4 I__3801 (
            .O(N__25875),
            .I(cmd_rdadctmp_13_adj_1437));
    LocalMux I__3800 (
            .O(N__25870),
            .I(cmd_rdadctmp_13_adj_1437));
    InMux I__3799 (
            .O(N__25865),
            .I(N__25862));
    LocalMux I__3798 (
            .O(N__25862),
            .I(N__25857));
    InMux I__3797 (
            .O(N__25861),
            .I(N__25854));
    InMux I__3796 (
            .O(N__25860),
            .I(N__25851));
    Span4Mux_h I__3795 (
            .O(N__25857),
            .I(N__25846));
    LocalMux I__3794 (
            .O(N__25854),
            .I(N__25846));
    LocalMux I__3793 (
            .O(N__25851),
            .I(buf_adcdata_iac_5));
    Odrv4 I__3792 (
            .O(N__25846),
            .I(buf_adcdata_iac_5));
    InMux I__3791 (
            .O(N__25841),
            .I(N__25838));
    LocalMux I__3790 (
            .O(N__25838),
            .I(N__25835));
    Span4Mux_h I__3789 (
            .O(N__25835),
            .I(N__25832));
    Odrv4 I__3788 (
            .O(N__25832),
            .I(buf_data_iac_5));
    InMux I__3787 (
            .O(N__25829),
            .I(N__25826));
    LocalMux I__3786 (
            .O(N__25826),
            .I(N__25823));
    Odrv4 I__3785 (
            .O(N__25823),
            .I(n22_adj_1632));
    InMux I__3784 (
            .O(N__25820),
            .I(N__25817));
    LocalMux I__3783 (
            .O(N__25817),
            .I(N__25814));
    Span4Mux_v I__3782 (
            .O(N__25814),
            .I(N__25811));
    Span4Mux_h I__3781 (
            .O(N__25811),
            .I(N__25808));
    Odrv4 I__3780 (
            .O(N__25808),
            .I(\ADC_VDC.n21718 ));
    CascadeMux I__3779 (
            .O(N__25805),
            .I(n12383_cascade_));
    InMux I__3778 (
            .O(N__25802),
            .I(N__25799));
    LocalMux I__3777 (
            .O(N__25799),
            .I(N__25794));
    InMux I__3776 (
            .O(N__25798),
            .I(N__25791));
    InMux I__3775 (
            .O(N__25797),
            .I(N__25788));
    Odrv4 I__3774 (
            .O(N__25794),
            .I(buf_dds1_10));
    LocalMux I__3773 (
            .O(N__25791),
            .I(buf_dds1_10));
    LocalMux I__3772 (
            .O(N__25788),
            .I(buf_dds1_10));
    InMux I__3771 (
            .O(N__25781),
            .I(N__25777));
    InMux I__3770 (
            .O(N__25780),
            .I(N__25774));
    LocalMux I__3769 (
            .O(N__25777),
            .I(n20673));
    LocalMux I__3768 (
            .O(N__25774),
            .I(n20673));
    CascadeMux I__3767 (
            .O(N__25769),
            .I(n11412_cascade_));
    IoInMux I__3766 (
            .O(N__25766),
            .I(N__25763));
    LocalMux I__3765 (
            .O(N__25763),
            .I(N__25760));
    IoSpan4Mux I__3764 (
            .O(N__25760),
            .I(N__25757));
    IoSpan4Mux I__3763 (
            .O(N__25757),
            .I(N__25754));
    Span4Mux_s2_v I__3762 (
            .O(N__25754),
            .I(N__25751));
    Span4Mux_v I__3761 (
            .O(N__25751),
            .I(N__25748));
    Odrv4 I__3760 (
            .O(N__25748),
            .I(AC_ADC_SYNC));
    InMux I__3759 (
            .O(N__25745),
            .I(N__25741));
    InMux I__3758 (
            .O(N__25744),
            .I(N__25737));
    LocalMux I__3757 (
            .O(N__25741),
            .I(N__25734));
    InMux I__3756 (
            .O(N__25740),
            .I(N__25731));
    LocalMux I__3755 (
            .O(N__25737),
            .I(buf_dds1_4));
    Odrv4 I__3754 (
            .O(N__25734),
            .I(buf_dds1_4));
    LocalMux I__3753 (
            .O(N__25731),
            .I(buf_dds1_4));
    CascadeMux I__3752 (
            .O(N__25724),
            .I(n8_adj_1555_cascade_));
    CascadeMux I__3751 (
            .O(N__25721),
            .I(N__25718));
    CascadeBuf I__3750 (
            .O(N__25718),
            .I(N__25715));
    CascadeMux I__3749 (
            .O(N__25715),
            .I(N__25712));
    CascadeBuf I__3748 (
            .O(N__25712),
            .I(N__25709));
    CascadeMux I__3747 (
            .O(N__25709),
            .I(N__25706));
    CascadeBuf I__3746 (
            .O(N__25706),
            .I(N__25703));
    CascadeMux I__3745 (
            .O(N__25703),
            .I(N__25700));
    CascadeBuf I__3744 (
            .O(N__25700),
            .I(N__25697));
    CascadeMux I__3743 (
            .O(N__25697),
            .I(N__25694));
    CascadeBuf I__3742 (
            .O(N__25694),
            .I(N__25691));
    CascadeMux I__3741 (
            .O(N__25691),
            .I(N__25688));
    CascadeBuf I__3740 (
            .O(N__25688),
            .I(N__25685));
    CascadeMux I__3739 (
            .O(N__25685),
            .I(N__25682));
    CascadeBuf I__3738 (
            .O(N__25682),
            .I(N__25679));
    CascadeMux I__3737 (
            .O(N__25679),
            .I(N__25676));
    CascadeBuf I__3736 (
            .O(N__25676),
            .I(N__25672));
    CascadeMux I__3735 (
            .O(N__25675),
            .I(N__25669));
    CascadeMux I__3734 (
            .O(N__25672),
            .I(N__25666));
    CascadeBuf I__3733 (
            .O(N__25669),
            .I(N__25663));
    CascadeBuf I__3732 (
            .O(N__25666),
            .I(N__25660));
    CascadeMux I__3731 (
            .O(N__25663),
            .I(N__25657));
    CascadeMux I__3730 (
            .O(N__25660),
            .I(N__25654));
    InMux I__3729 (
            .O(N__25657),
            .I(N__25651));
    InMux I__3728 (
            .O(N__25654),
            .I(N__25648));
    LocalMux I__3727 (
            .O(N__25651),
            .I(N__25645));
    LocalMux I__3726 (
            .O(N__25648),
            .I(N__25642));
    Span12Mux_h I__3725 (
            .O(N__25645),
            .I(N__25639));
    Span12Mux_v I__3724 (
            .O(N__25642),
            .I(N__25636));
    Span12Mux_v I__3723 (
            .O(N__25639),
            .I(N__25633));
    Span12Mux_h I__3722 (
            .O(N__25636),
            .I(N__25630));
    Odrv12 I__3721 (
            .O(N__25633),
            .I(data_index_9_N_216_8));
    Odrv12 I__3720 (
            .O(N__25630),
            .I(data_index_9_N_216_8));
    InMux I__3719 (
            .O(N__25625),
            .I(N__25622));
    LocalMux I__3718 (
            .O(N__25622),
            .I(n8_adj_1555));
    InMux I__3717 (
            .O(N__25619),
            .I(N__25616));
    LocalMux I__3716 (
            .O(N__25616),
            .I(N__25613));
    Odrv4 I__3715 (
            .O(N__25613),
            .I(n22040));
    InMux I__3714 (
            .O(N__25610),
            .I(N__25605));
    InMux I__3713 (
            .O(N__25609),
            .I(N__25602));
    InMux I__3712 (
            .O(N__25608),
            .I(N__25599));
    LocalMux I__3711 (
            .O(N__25605),
            .I(buf_dds1_9));
    LocalMux I__3710 (
            .O(N__25602),
            .I(buf_dds1_9));
    LocalMux I__3709 (
            .O(N__25599),
            .I(buf_dds1_9));
    InMux I__3708 (
            .O(N__25592),
            .I(N__25588));
    InMux I__3707 (
            .O(N__25591),
            .I(N__25584));
    LocalMux I__3706 (
            .O(N__25588),
            .I(N__25581));
    InMux I__3705 (
            .O(N__25587),
            .I(N__25578));
    LocalMux I__3704 (
            .O(N__25584),
            .I(buf_dds1_8));
    Odrv4 I__3703 (
            .O(N__25581),
            .I(buf_dds1_8));
    LocalMux I__3702 (
            .O(N__25578),
            .I(buf_dds1_8));
    InMux I__3701 (
            .O(N__25571),
            .I(N__25568));
    LocalMux I__3700 (
            .O(N__25568),
            .I(n20849));
    CascadeMux I__3699 (
            .O(N__25565),
            .I(N__25562));
    InMux I__3698 (
            .O(N__25562),
            .I(N__25559));
    LocalMux I__3697 (
            .O(N__25559),
            .I(n22103));
    InMux I__3696 (
            .O(N__25556),
            .I(N__25553));
    LocalMux I__3695 (
            .O(N__25553),
            .I(N__25550));
    Span4Mux_v I__3694 (
            .O(N__25550),
            .I(N__25547));
    Sp12to4 I__3693 (
            .O(N__25547),
            .I(N__25542));
    CascadeMux I__3692 (
            .O(N__25546),
            .I(N__25539));
    InMux I__3691 (
            .O(N__25545),
            .I(N__25536));
    Span12Mux_h I__3690 (
            .O(N__25542),
            .I(N__25533));
    InMux I__3689 (
            .O(N__25539),
            .I(N__25530));
    LocalMux I__3688 (
            .O(N__25536),
            .I(buf_adcdata_iac_17));
    Odrv12 I__3687 (
            .O(N__25533),
            .I(buf_adcdata_iac_17));
    LocalMux I__3686 (
            .O(N__25530),
            .I(buf_adcdata_iac_17));
    InMux I__3685 (
            .O(N__25523),
            .I(N__25520));
    LocalMux I__3684 (
            .O(N__25520),
            .I(N__25517));
    Span12Mux_v I__3683 (
            .O(N__25517),
            .I(N__25514));
    Span12Mux_h I__3682 (
            .O(N__25514),
            .I(N__25511));
    Odrv12 I__3681 (
            .O(N__25511),
            .I(buf_data_iac_21));
    CascadeMux I__3680 (
            .O(N__25508),
            .I(n20876_cascade_));
    InMux I__3679 (
            .O(N__25505),
            .I(N__25502));
    LocalMux I__3678 (
            .O(N__25502),
            .I(n22106));
    InMux I__3677 (
            .O(N__25499),
            .I(N__25496));
    LocalMux I__3676 (
            .O(N__25496),
            .I(n20875));
    InMux I__3675 (
            .O(N__25493),
            .I(N__25490));
    LocalMux I__3674 (
            .O(N__25490),
            .I(n22022));
    InMux I__3673 (
            .O(N__25487),
            .I(N__25484));
    LocalMux I__3672 (
            .O(N__25484),
            .I(N__25480));
    InMux I__3671 (
            .O(N__25483),
            .I(N__25477));
    Span4Mux_v I__3670 (
            .O(N__25480),
            .I(N__25474));
    LocalMux I__3669 (
            .O(N__25477),
            .I(N__25471));
    Sp12to4 I__3668 (
            .O(N__25474),
            .I(N__25467));
    Span4Mux_v I__3667 (
            .O(N__25471),
            .I(N__25464));
    InMux I__3666 (
            .O(N__25470),
            .I(N__25461));
    Span12Mux_h I__3665 (
            .O(N__25467),
            .I(N__25458));
    Span4Mux_v I__3664 (
            .O(N__25464),
            .I(N__25455));
    LocalMux I__3663 (
            .O(N__25461),
            .I(buf_adcdata_vac_21));
    Odrv12 I__3662 (
            .O(N__25458),
            .I(buf_adcdata_vac_21));
    Odrv4 I__3661 (
            .O(N__25455),
            .I(buf_adcdata_vac_21));
    CascadeMux I__3660 (
            .O(N__25448),
            .I(N__25445));
    InMux I__3659 (
            .O(N__25445),
            .I(N__25442));
    LocalMux I__3658 (
            .O(N__25442),
            .I(N__25439));
    Span4Mux_v I__3657 (
            .O(N__25439),
            .I(N__25436));
    Span4Mux_v I__3656 (
            .O(N__25436),
            .I(N__25432));
    InMux I__3655 (
            .O(N__25435),
            .I(N__25429));
    Odrv4 I__3654 (
            .O(N__25432),
            .I(buf_adcdata_vdc_21));
    LocalMux I__3653 (
            .O(N__25429),
            .I(buf_adcdata_vdc_21));
    InMux I__3652 (
            .O(N__25424),
            .I(N__25421));
    LocalMux I__3651 (
            .O(N__25421),
            .I(n22184));
    CascadeMux I__3650 (
            .O(N__25418),
            .I(N__25415));
    InMux I__3649 (
            .O(N__25415),
            .I(N__25412));
    LocalMux I__3648 (
            .O(N__25412),
            .I(N__25409));
    Span4Mux_h I__3647 (
            .O(N__25409),
            .I(N__25405));
    InMux I__3646 (
            .O(N__25408),
            .I(N__25402));
    Odrv4 I__3645 (
            .O(N__25405),
            .I(buf_readRTD_12));
    LocalMux I__3644 (
            .O(N__25402),
            .I(buf_readRTD_12));
    InMux I__3643 (
            .O(N__25397),
            .I(N__25394));
    LocalMux I__3642 (
            .O(N__25394),
            .I(N__25391));
    Span4Mux_v I__3641 (
            .O(N__25391),
            .I(N__25388));
    Odrv4 I__3640 (
            .O(N__25388),
            .I(n22202));
    CascadeMux I__3639 (
            .O(N__25385),
            .I(N__25382));
    InMux I__3638 (
            .O(N__25382),
            .I(N__25379));
    LocalMux I__3637 (
            .O(N__25379),
            .I(N__25376));
    Span4Mux_h I__3636 (
            .O(N__25376),
            .I(N__25372));
    InMux I__3635 (
            .O(N__25375),
            .I(N__25369));
    Odrv4 I__3634 (
            .O(N__25372),
            .I(buf_readRTD_8));
    LocalMux I__3633 (
            .O(N__25369),
            .I(buf_readRTD_8));
    CascadeMux I__3632 (
            .O(N__25364),
            .I(N__25361));
    InMux I__3631 (
            .O(N__25361),
            .I(N__25356));
    InMux I__3630 (
            .O(N__25360),
            .I(N__25353));
    CascadeMux I__3629 (
            .O(N__25359),
            .I(N__25350));
    LocalMux I__3628 (
            .O(N__25356),
            .I(N__25347));
    LocalMux I__3627 (
            .O(N__25353),
            .I(N__25344));
    InMux I__3626 (
            .O(N__25350),
            .I(N__25341));
    Span4Mux_v I__3625 (
            .O(N__25347),
            .I(N__25333));
    Span4Mux_h I__3624 (
            .O(N__25344),
            .I(N__25333));
    LocalMux I__3623 (
            .O(N__25341),
            .I(N__25333));
    InMux I__3622 (
            .O(N__25340),
            .I(N__25329));
    Span4Mux_v I__3621 (
            .O(N__25333),
            .I(N__25326));
    InMux I__3620 (
            .O(N__25332),
            .I(N__25323));
    LocalMux I__3619 (
            .O(N__25329),
            .I(N__25320));
    Odrv4 I__3618 (
            .O(N__25326),
            .I(buf_cfgRTD_0));
    LocalMux I__3617 (
            .O(N__25323),
            .I(buf_cfgRTD_0));
    Odrv4 I__3616 (
            .O(N__25320),
            .I(buf_cfgRTD_0));
    CascadeMux I__3615 (
            .O(N__25313),
            .I(N__25310));
    InMux I__3614 (
            .O(N__25310),
            .I(N__25307));
    LocalMux I__3613 (
            .O(N__25307),
            .I(N__25304));
    Span4Mux_v I__3612 (
            .O(N__25304),
            .I(N__25301));
    Span4Mux_h I__3611 (
            .O(N__25301),
            .I(N__25298));
    Span4Mux_h I__3610 (
            .O(N__25298),
            .I(N__25293));
    InMux I__3609 (
            .O(N__25297),
            .I(N__25290));
    InMux I__3608 (
            .O(N__25296),
            .I(N__25287));
    Odrv4 I__3607 (
            .O(N__25293),
            .I(cmd_rdadctmp_27_adj_1423));
    LocalMux I__3606 (
            .O(N__25290),
            .I(cmd_rdadctmp_27_adj_1423));
    LocalMux I__3605 (
            .O(N__25287),
            .I(cmd_rdadctmp_27_adj_1423));
    InMux I__3604 (
            .O(N__25280),
            .I(N__25277));
    LocalMux I__3603 (
            .O(N__25277),
            .I(N__25272));
    InMux I__3602 (
            .O(N__25276),
            .I(N__25269));
    InMux I__3601 (
            .O(N__25275),
            .I(N__25266));
    Span4Mux_v I__3600 (
            .O(N__25272),
            .I(N__25261));
    LocalMux I__3599 (
            .O(N__25269),
            .I(N__25261));
    LocalMux I__3598 (
            .O(N__25266),
            .I(buf_dds1_15));
    Odrv4 I__3597 (
            .O(N__25261),
            .I(buf_dds1_15));
    CascadeMux I__3596 (
            .O(N__25256),
            .I(N__25252));
    CascadeMux I__3595 (
            .O(N__25255),
            .I(N__25249));
    InMux I__3594 (
            .O(N__25252),
            .I(N__25245));
    InMux I__3593 (
            .O(N__25249),
            .I(N__25242));
    CascadeMux I__3592 (
            .O(N__25248),
            .I(N__25239));
    LocalMux I__3591 (
            .O(N__25245),
            .I(N__25236));
    LocalMux I__3590 (
            .O(N__25242),
            .I(N__25233));
    InMux I__3589 (
            .O(N__25239),
            .I(N__25230));
    Span4Mux_h I__3588 (
            .O(N__25236),
            .I(N__25225));
    Span4Mux_v I__3587 (
            .O(N__25233),
            .I(N__25220));
    LocalMux I__3586 (
            .O(N__25230),
            .I(N__25220));
    InMux I__3585 (
            .O(N__25229),
            .I(N__25217));
    InMux I__3584 (
            .O(N__25228),
            .I(N__25214));
    Odrv4 I__3583 (
            .O(N__25225),
            .I(buf_cfgRTD_4));
    Odrv4 I__3582 (
            .O(N__25220),
            .I(buf_cfgRTD_4));
    LocalMux I__3581 (
            .O(N__25217),
            .I(buf_cfgRTD_4));
    LocalMux I__3580 (
            .O(N__25214),
            .I(buf_cfgRTD_4));
    InMux I__3579 (
            .O(N__25205),
            .I(N__25201));
    InMux I__3578 (
            .O(N__25204),
            .I(N__25198));
    LocalMux I__3577 (
            .O(N__25201),
            .I(N__25191));
    LocalMux I__3576 (
            .O(N__25198),
            .I(N__25191));
    InMux I__3575 (
            .O(N__25197),
            .I(N__25188));
    InMux I__3574 (
            .O(N__25196),
            .I(N__25184));
    Span4Mux_v I__3573 (
            .O(N__25191),
            .I(N__25181));
    LocalMux I__3572 (
            .O(N__25188),
            .I(N__25178));
    InMux I__3571 (
            .O(N__25187),
            .I(N__25175));
    LocalMux I__3570 (
            .O(N__25184),
            .I(N__25172));
    Odrv4 I__3569 (
            .O(N__25181),
            .I(buf_cfgRTD_3));
    Odrv4 I__3568 (
            .O(N__25178),
            .I(buf_cfgRTD_3));
    LocalMux I__3567 (
            .O(N__25175),
            .I(buf_cfgRTD_3));
    Odrv12 I__3566 (
            .O(N__25172),
            .I(buf_cfgRTD_3));
    InMux I__3565 (
            .O(N__25163),
            .I(N__25160));
    LocalMux I__3564 (
            .O(N__25160),
            .I(N__25156));
    CascadeMux I__3563 (
            .O(N__25159),
            .I(N__25153));
    Span4Mux_h I__3562 (
            .O(N__25156),
            .I(N__25150));
    InMux I__3561 (
            .O(N__25153),
            .I(N__25147));
    Odrv4 I__3560 (
            .O(N__25150),
            .I(cmd_rdadctmp_7_adj_1443));
    LocalMux I__3559 (
            .O(N__25147),
            .I(cmd_rdadctmp_7_adj_1443));
    CascadeMux I__3558 (
            .O(N__25142),
            .I(N__25139));
    InMux I__3557 (
            .O(N__25139),
            .I(N__25136));
    LocalMux I__3556 (
            .O(N__25136),
            .I(N__25133));
    Span4Mux_h I__3555 (
            .O(N__25133),
            .I(N__25129));
    InMux I__3554 (
            .O(N__25132),
            .I(N__25126));
    Odrv4 I__3553 (
            .O(N__25129),
            .I(buf_readRTD_13));
    LocalMux I__3552 (
            .O(N__25126),
            .I(buf_readRTD_13));
    InMux I__3551 (
            .O(N__25121),
            .I(N__25117));
    InMux I__3550 (
            .O(N__25120),
            .I(N__25114));
    LocalMux I__3549 (
            .O(N__25117),
            .I(N__25111));
    LocalMux I__3548 (
            .O(N__25114),
            .I(N__25108));
    Odrv4 I__3547 (
            .O(N__25111),
            .I(buf_readRTD_10));
    Odrv4 I__3546 (
            .O(N__25108),
            .I(buf_readRTD_10));
    InMux I__3545 (
            .O(N__25103),
            .I(N__25099));
    CascadeMux I__3544 (
            .O(N__25102),
            .I(N__25096));
    LocalMux I__3543 (
            .O(N__25099),
            .I(N__25092));
    InMux I__3542 (
            .O(N__25096),
            .I(N__25089));
    CascadeMux I__3541 (
            .O(N__25095),
            .I(N__25086));
    Span4Mux_v I__3540 (
            .O(N__25092),
            .I(N__25081));
    LocalMux I__3539 (
            .O(N__25089),
            .I(N__25078));
    InMux I__3538 (
            .O(N__25086),
            .I(N__25075));
    InMux I__3537 (
            .O(N__25085),
            .I(N__25072));
    InMux I__3536 (
            .O(N__25084),
            .I(N__25069));
    Odrv4 I__3535 (
            .O(N__25081),
            .I(buf_cfgRTD_2));
    Odrv4 I__3534 (
            .O(N__25078),
            .I(buf_cfgRTD_2));
    LocalMux I__3533 (
            .O(N__25075),
            .I(buf_cfgRTD_2));
    LocalMux I__3532 (
            .O(N__25072),
            .I(buf_cfgRTD_2));
    LocalMux I__3531 (
            .O(N__25069),
            .I(buf_cfgRTD_2));
    InMux I__3530 (
            .O(N__25058),
            .I(N__25055));
    LocalMux I__3529 (
            .O(N__25055),
            .I(N__25052));
    Odrv4 I__3528 (
            .O(N__25052),
            .I(n20834));
    CascadeMux I__3527 (
            .O(N__25049),
            .I(N__25044));
    CascadeMux I__3526 (
            .O(N__25048),
            .I(N__25041));
    InMux I__3525 (
            .O(N__25047),
            .I(N__25035));
    InMux I__3524 (
            .O(N__25044),
            .I(N__25027));
    InMux I__3523 (
            .O(N__25041),
            .I(N__25024));
    InMux I__3522 (
            .O(N__25040),
            .I(N__25021));
    InMux I__3521 (
            .O(N__25039),
            .I(N__25006));
    InMux I__3520 (
            .O(N__25038),
            .I(N__25003));
    LocalMux I__3519 (
            .O(N__25035),
            .I(N__25000));
    InMux I__3518 (
            .O(N__25034),
            .I(N__24989));
    InMux I__3517 (
            .O(N__25033),
            .I(N__24989));
    InMux I__3516 (
            .O(N__25032),
            .I(N__24989));
    InMux I__3515 (
            .O(N__25031),
            .I(N__24989));
    InMux I__3514 (
            .O(N__25030),
            .I(N__24989));
    LocalMux I__3513 (
            .O(N__25027),
            .I(N__24984));
    LocalMux I__3512 (
            .O(N__25024),
            .I(N__24984));
    LocalMux I__3511 (
            .O(N__25021),
            .I(N__24981));
    InMux I__3510 (
            .O(N__25020),
            .I(N__24976));
    InMux I__3509 (
            .O(N__25019),
            .I(N__24976));
    InMux I__3508 (
            .O(N__25018),
            .I(N__24969));
    InMux I__3507 (
            .O(N__25017),
            .I(N__24969));
    InMux I__3506 (
            .O(N__25016),
            .I(N__24969));
    InMux I__3505 (
            .O(N__25015),
            .I(N__24960));
    InMux I__3504 (
            .O(N__25014),
            .I(N__24960));
    InMux I__3503 (
            .O(N__25013),
            .I(N__24960));
    InMux I__3502 (
            .O(N__25012),
            .I(N__24960));
    InMux I__3501 (
            .O(N__25011),
            .I(N__24953));
    InMux I__3500 (
            .O(N__25010),
            .I(N__24953));
    InMux I__3499 (
            .O(N__25009),
            .I(N__24953));
    LocalMux I__3498 (
            .O(N__25006),
            .I(N__24944));
    LocalMux I__3497 (
            .O(N__25003),
            .I(N__24944));
    Span4Mux_h I__3496 (
            .O(N__25000),
            .I(N__24944));
    LocalMux I__3495 (
            .O(N__24989),
            .I(N__24944));
    Odrv4 I__3494 (
            .O(N__24984),
            .I(adc_state_1_adj_1483));
    Odrv4 I__3493 (
            .O(N__24981),
            .I(adc_state_1_adj_1483));
    LocalMux I__3492 (
            .O(N__24976),
            .I(adc_state_1_adj_1483));
    LocalMux I__3491 (
            .O(N__24969),
            .I(adc_state_1_adj_1483));
    LocalMux I__3490 (
            .O(N__24960),
            .I(adc_state_1_adj_1483));
    LocalMux I__3489 (
            .O(N__24953),
            .I(adc_state_1_adj_1483));
    Odrv4 I__3488 (
            .O(N__24944),
            .I(adc_state_1_adj_1483));
    InMux I__3487 (
            .O(N__24929),
            .I(N__24925));
    InMux I__3486 (
            .O(N__24928),
            .I(N__24922));
    LocalMux I__3485 (
            .O(N__24925),
            .I(\RTD.n20656 ));
    LocalMux I__3484 (
            .O(N__24922),
            .I(\RTD.n20656 ));
    CascadeMux I__3483 (
            .O(N__24917),
            .I(n12397_cascade_));
    InMux I__3482 (
            .O(N__24914),
            .I(N__24911));
    LocalMux I__3481 (
            .O(N__24911),
            .I(N__24908));
    Odrv4 I__3480 (
            .O(N__24908),
            .I(\RTD.n10 ));
    InMux I__3479 (
            .O(N__24905),
            .I(N__24901));
    InMux I__3478 (
            .O(N__24904),
            .I(N__24898));
    LocalMux I__3477 (
            .O(N__24901),
            .I(\RTD.cfg_buf_2 ));
    LocalMux I__3476 (
            .O(N__24898),
            .I(\RTD.cfg_buf_2 ));
    InMux I__3475 (
            .O(N__24893),
            .I(N__24889));
    InMux I__3474 (
            .O(N__24892),
            .I(N__24886));
    LocalMux I__3473 (
            .O(N__24889),
            .I(N__24882));
    LocalMux I__3472 (
            .O(N__24886),
            .I(N__24879));
    InMux I__3471 (
            .O(N__24885),
            .I(N__24876));
    Span4Mux_v I__3470 (
            .O(N__24882),
            .I(N__24871));
    Span4Mux_h I__3469 (
            .O(N__24879),
            .I(N__24871));
    LocalMux I__3468 (
            .O(N__24876),
            .I(read_buf_0));
    Odrv4 I__3467 (
            .O(N__24871),
            .I(read_buf_0));
    CascadeMux I__3466 (
            .O(N__24866),
            .I(N__24860));
    CascadeMux I__3465 (
            .O(N__24865),
            .I(N__24857));
    CascadeMux I__3464 (
            .O(N__24864),
            .I(N__24854));
    CascadeMux I__3463 (
            .O(N__24863),
            .I(N__24851));
    InMux I__3462 (
            .O(N__24860),
            .I(N__24826));
    InMux I__3461 (
            .O(N__24857),
            .I(N__24826));
    InMux I__3460 (
            .O(N__24854),
            .I(N__24826));
    InMux I__3459 (
            .O(N__24851),
            .I(N__24826));
    InMux I__3458 (
            .O(N__24850),
            .I(N__24826));
    InMux I__3457 (
            .O(N__24849),
            .I(N__24826));
    InMux I__3456 (
            .O(N__24848),
            .I(N__24823));
    InMux I__3455 (
            .O(N__24847),
            .I(N__24814));
    InMux I__3454 (
            .O(N__24846),
            .I(N__24814));
    InMux I__3453 (
            .O(N__24845),
            .I(N__24814));
    InMux I__3452 (
            .O(N__24844),
            .I(N__24814));
    InMux I__3451 (
            .O(N__24843),
            .I(N__24809));
    InMux I__3450 (
            .O(N__24842),
            .I(N__24809));
    InMux I__3449 (
            .O(N__24841),
            .I(N__24786));
    InMux I__3448 (
            .O(N__24840),
            .I(N__24786));
    InMux I__3447 (
            .O(N__24839),
            .I(N__24786));
    LocalMux I__3446 (
            .O(N__24826),
            .I(N__24781));
    LocalMux I__3445 (
            .O(N__24823),
            .I(N__24781));
    LocalMux I__3444 (
            .O(N__24814),
            .I(N__24776));
    LocalMux I__3443 (
            .O(N__24809),
            .I(N__24776));
    InMux I__3442 (
            .O(N__24808),
            .I(N__24773));
    CascadeMux I__3441 (
            .O(N__24807),
            .I(N__24770));
    CascadeMux I__3440 (
            .O(N__24806),
            .I(N__24766));
    InMux I__3439 (
            .O(N__24805),
            .I(N__24756));
    InMux I__3438 (
            .O(N__24804),
            .I(N__24756));
    InMux I__3437 (
            .O(N__24803),
            .I(N__24756));
    InMux I__3436 (
            .O(N__24802),
            .I(N__24756));
    InMux I__3435 (
            .O(N__24801),
            .I(N__24751));
    InMux I__3434 (
            .O(N__24800),
            .I(N__24751));
    InMux I__3433 (
            .O(N__24799),
            .I(N__24748));
    InMux I__3432 (
            .O(N__24798),
            .I(N__24745));
    InMux I__3431 (
            .O(N__24797),
            .I(N__24742));
    InMux I__3430 (
            .O(N__24796),
            .I(N__24739));
    InMux I__3429 (
            .O(N__24795),
            .I(N__24736));
    InMux I__3428 (
            .O(N__24794),
            .I(N__24731));
    InMux I__3427 (
            .O(N__24793),
            .I(N__24731));
    LocalMux I__3426 (
            .O(N__24786),
            .I(N__24724));
    Span4Mux_v I__3425 (
            .O(N__24781),
            .I(N__24724));
    Span4Mux_h I__3424 (
            .O(N__24776),
            .I(N__24724));
    LocalMux I__3423 (
            .O(N__24773),
            .I(N__24721));
    InMux I__3422 (
            .O(N__24770),
            .I(N__24716));
    InMux I__3421 (
            .O(N__24769),
            .I(N__24716));
    InMux I__3420 (
            .O(N__24766),
            .I(N__24711));
    InMux I__3419 (
            .O(N__24765),
            .I(N__24711));
    LocalMux I__3418 (
            .O(N__24756),
            .I(N__24708));
    LocalMux I__3417 (
            .O(N__24751),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3416 (
            .O(N__24748),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3415 (
            .O(N__24745),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3414 (
            .O(N__24742),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3413 (
            .O(N__24739),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3412 (
            .O(N__24736),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3411 (
            .O(N__24731),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3410 (
            .O(N__24724),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3409 (
            .O(N__24721),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3408 (
            .O(N__24716),
            .I(\RTD.adc_state_0 ));
    LocalMux I__3407 (
            .O(N__24711),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__3406 (
            .O(N__24708),
            .I(\RTD.adc_state_0 ));
    CascadeMux I__3405 (
            .O(N__24683),
            .I(N__24670));
    CascadeMux I__3404 (
            .O(N__24682),
            .I(N__24667));
    CascadeMux I__3403 (
            .O(N__24681),
            .I(N__24661));
    CascadeMux I__3402 (
            .O(N__24680),
            .I(N__24655));
    CascadeMux I__3401 (
            .O(N__24679),
            .I(N__24652));
    CascadeMux I__3400 (
            .O(N__24678),
            .I(N__24649));
    CascadeMux I__3399 (
            .O(N__24677),
            .I(N__24645));
    InMux I__3398 (
            .O(N__24676),
            .I(N__24640));
    CascadeMux I__3397 (
            .O(N__24675),
            .I(N__24637));
    InMux I__3396 (
            .O(N__24674),
            .I(N__24631));
    InMux I__3395 (
            .O(N__24673),
            .I(N__24628));
    InMux I__3394 (
            .O(N__24670),
            .I(N__24621));
    InMux I__3393 (
            .O(N__24667),
            .I(N__24621));
    InMux I__3392 (
            .O(N__24666),
            .I(N__24621));
    InMux I__3391 (
            .O(N__24665),
            .I(N__24616));
    InMux I__3390 (
            .O(N__24664),
            .I(N__24616));
    InMux I__3389 (
            .O(N__24661),
            .I(N__24609));
    InMux I__3388 (
            .O(N__24660),
            .I(N__24609));
    InMux I__3387 (
            .O(N__24659),
            .I(N__24609));
    InMux I__3386 (
            .O(N__24658),
            .I(N__24606));
    InMux I__3385 (
            .O(N__24655),
            .I(N__24603));
    InMux I__3384 (
            .O(N__24652),
            .I(N__24592));
    InMux I__3383 (
            .O(N__24649),
            .I(N__24592));
    InMux I__3382 (
            .O(N__24648),
            .I(N__24592));
    InMux I__3381 (
            .O(N__24645),
            .I(N__24592));
    InMux I__3380 (
            .O(N__24644),
            .I(N__24592));
    InMux I__3379 (
            .O(N__24643),
            .I(N__24588));
    LocalMux I__3378 (
            .O(N__24640),
            .I(N__24585));
    InMux I__3377 (
            .O(N__24637),
            .I(N__24579));
    InMux I__3376 (
            .O(N__24636),
            .I(N__24579));
    InMux I__3375 (
            .O(N__24635),
            .I(N__24574));
    InMux I__3374 (
            .O(N__24634),
            .I(N__24574));
    LocalMux I__3373 (
            .O(N__24631),
            .I(N__24571));
    LocalMux I__3372 (
            .O(N__24628),
            .I(N__24568));
    LocalMux I__3371 (
            .O(N__24621),
            .I(N__24561));
    LocalMux I__3370 (
            .O(N__24616),
            .I(N__24561));
    LocalMux I__3369 (
            .O(N__24609),
            .I(N__24561));
    LocalMux I__3368 (
            .O(N__24606),
            .I(N__24554));
    LocalMux I__3367 (
            .O(N__24603),
            .I(N__24554));
    LocalMux I__3366 (
            .O(N__24592),
            .I(N__24554));
    InMux I__3365 (
            .O(N__24591),
            .I(N__24551));
    LocalMux I__3364 (
            .O(N__24588),
            .I(N__24546));
    Span4Mux_v I__3363 (
            .O(N__24585),
            .I(N__24546));
    InMux I__3362 (
            .O(N__24584),
            .I(N__24543));
    LocalMux I__3361 (
            .O(N__24579),
            .I(N__24538));
    LocalMux I__3360 (
            .O(N__24574),
            .I(N__24538));
    Span4Mux_h I__3359 (
            .O(N__24571),
            .I(N__24529));
    Span4Mux_h I__3358 (
            .O(N__24568),
            .I(N__24529));
    Span4Mux_h I__3357 (
            .O(N__24561),
            .I(N__24529));
    Span4Mux_v I__3356 (
            .O(N__24554),
            .I(N__24529));
    LocalMux I__3355 (
            .O(N__24551),
            .I(adc_state_3_adj_1481));
    Odrv4 I__3354 (
            .O(N__24546),
            .I(adc_state_3_adj_1481));
    LocalMux I__3353 (
            .O(N__24543),
            .I(adc_state_3_adj_1481));
    Odrv12 I__3352 (
            .O(N__24538),
            .I(adc_state_3_adj_1481));
    Odrv4 I__3351 (
            .O(N__24529),
            .I(adc_state_3_adj_1481));
    SRMux I__3350 (
            .O(N__24518),
            .I(N__24515));
    LocalMux I__3349 (
            .O(N__24515),
            .I(N__24511));
    SRMux I__3348 (
            .O(N__24514),
            .I(N__24508));
    Span4Mux_h I__3347 (
            .O(N__24511),
            .I(N__24505));
    LocalMux I__3346 (
            .O(N__24508),
            .I(N__24502));
    Span4Mux_h I__3345 (
            .O(N__24505),
            .I(N__24499));
    Span4Mux_h I__3344 (
            .O(N__24502),
            .I(N__24496));
    Odrv4 I__3343 (
            .O(N__24499),
            .I(\RTD.n14717 ));
    Odrv4 I__3342 (
            .O(N__24496),
            .I(\RTD.n14717 ));
    InMux I__3341 (
            .O(N__24491),
            .I(N__24488));
    LocalMux I__3340 (
            .O(N__24488),
            .I(n16_adj_1524));
    InMux I__3339 (
            .O(N__24485),
            .I(N__24481));
    InMux I__3338 (
            .O(N__24484),
            .I(N__24478));
    LocalMux I__3337 (
            .O(N__24481),
            .I(\RTD.cfg_buf_4 ));
    LocalMux I__3336 (
            .O(N__24478),
            .I(\RTD.cfg_buf_4 ));
    InMux I__3335 (
            .O(N__24473),
            .I(N__24463));
    InMux I__3334 (
            .O(N__24472),
            .I(N__24456));
    InMux I__3333 (
            .O(N__24471),
            .I(N__24456));
    InMux I__3332 (
            .O(N__24470),
            .I(N__24456));
    InMux I__3331 (
            .O(N__24469),
            .I(N__24451));
    InMux I__3330 (
            .O(N__24468),
            .I(N__24451));
    CascadeMux I__3329 (
            .O(N__24467),
            .I(N__24428));
    InMux I__3328 (
            .O(N__24466),
            .I(N__24414));
    LocalMux I__3327 (
            .O(N__24463),
            .I(N__24406));
    LocalMux I__3326 (
            .O(N__24456),
            .I(N__24401));
    LocalMux I__3325 (
            .O(N__24451),
            .I(N__24401));
    InMux I__3324 (
            .O(N__24450),
            .I(N__24394));
    InMux I__3323 (
            .O(N__24449),
            .I(N__24394));
    InMux I__3322 (
            .O(N__24448),
            .I(N__24394));
    InMux I__3321 (
            .O(N__24447),
            .I(N__24383));
    InMux I__3320 (
            .O(N__24446),
            .I(N__24383));
    InMux I__3319 (
            .O(N__24445),
            .I(N__24383));
    InMux I__3318 (
            .O(N__24444),
            .I(N__24383));
    InMux I__3317 (
            .O(N__24443),
            .I(N__24383));
    InMux I__3316 (
            .O(N__24442),
            .I(N__24372));
    InMux I__3315 (
            .O(N__24441),
            .I(N__24372));
    InMux I__3314 (
            .O(N__24440),
            .I(N__24372));
    InMux I__3313 (
            .O(N__24439),
            .I(N__24372));
    InMux I__3312 (
            .O(N__24438),
            .I(N__24372));
    InMux I__3311 (
            .O(N__24437),
            .I(N__24362));
    InMux I__3310 (
            .O(N__24436),
            .I(N__24362));
    InMux I__3309 (
            .O(N__24435),
            .I(N__24362));
    InMux I__3308 (
            .O(N__24434),
            .I(N__24351));
    InMux I__3307 (
            .O(N__24433),
            .I(N__24351));
    InMux I__3306 (
            .O(N__24432),
            .I(N__24351));
    InMux I__3305 (
            .O(N__24431),
            .I(N__24351));
    InMux I__3304 (
            .O(N__24428),
            .I(N__24351));
    InMux I__3303 (
            .O(N__24427),
            .I(N__24334));
    InMux I__3302 (
            .O(N__24426),
            .I(N__24334));
    InMux I__3301 (
            .O(N__24425),
            .I(N__24334));
    InMux I__3300 (
            .O(N__24424),
            .I(N__24334));
    InMux I__3299 (
            .O(N__24423),
            .I(N__24334));
    InMux I__3298 (
            .O(N__24422),
            .I(N__24334));
    InMux I__3297 (
            .O(N__24421),
            .I(N__24334));
    InMux I__3296 (
            .O(N__24420),
            .I(N__24334));
    InMux I__3295 (
            .O(N__24419),
            .I(N__24329));
    InMux I__3294 (
            .O(N__24418),
            .I(N__24329));
    InMux I__3293 (
            .O(N__24417),
            .I(N__24326));
    LocalMux I__3292 (
            .O(N__24414),
            .I(N__24323));
    InMux I__3291 (
            .O(N__24413),
            .I(N__24316));
    InMux I__3290 (
            .O(N__24412),
            .I(N__24316));
    InMux I__3289 (
            .O(N__24411),
            .I(N__24316));
    InMux I__3288 (
            .O(N__24410),
            .I(N__24311));
    InMux I__3287 (
            .O(N__24409),
            .I(N__24311));
    Span4Mux_v I__3286 (
            .O(N__24406),
            .I(N__24302));
    Span4Mux_v I__3285 (
            .O(N__24401),
            .I(N__24302));
    LocalMux I__3284 (
            .O(N__24394),
            .I(N__24302));
    LocalMux I__3283 (
            .O(N__24383),
            .I(N__24302));
    LocalMux I__3282 (
            .O(N__24372),
            .I(N__24299));
    InMux I__3281 (
            .O(N__24371),
            .I(N__24292));
    InMux I__3280 (
            .O(N__24370),
            .I(N__24292));
    InMux I__3279 (
            .O(N__24369),
            .I(N__24292));
    LocalMux I__3278 (
            .O(N__24362),
            .I(N__24287));
    LocalMux I__3277 (
            .O(N__24351),
            .I(N__24287));
    LocalMux I__3276 (
            .O(N__24334),
            .I(adc_state_2_adj_1482));
    LocalMux I__3275 (
            .O(N__24329),
            .I(adc_state_2_adj_1482));
    LocalMux I__3274 (
            .O(N__24326),
            .I(adc_state_2_adj_1482));
    Odrv4 I__3273 (
            .O(N__24323),
            .I(adc_state_2_adj_1482));
    LocalMux I__3272 (
            .O(N__24316),
            .I(adc_state_2_adj_1482));
    LocalMux I__3271 (
            .O(N__24311),
            .I(adc_state_2_adj_1482));
    Odrv4 I__3270 (
            .O(N__24302),
            .I(adc_state_2_adj_1482));
    Odrv4 I__3269 (
            .O(N__24299),
            .I(adc_state_2_adj_1482));
    LocalMux I__3268 (
            .O(N__24292),
            .I(adc_state_2_adj_1482));
    Odrv4 I__3267 (
            .O(N__24287),
            .I(adc_state_2_adj_1482));
    CascadeMux I__3266 (
            .O(N__24266),
            .I(N__24263));
    InMux I__3265 (
            .O(N__24263),
            .I(N__24260));
    LocalMux I__3264 (
            .O(N__24260),
            .I(N__24255));
    CascadeMux I__3263 (
            .O(N__24259),
            .I(N__24252));
    CascadeMux I__3262 (
            .O(N__24258),
            .I(N__24249));
    Span4Mux_h I__3261 (
            .O(N__24255),
            .I(N__24246));
    InMux I__3260 (
            .O(N__24252),
            .I(N__24241));
    InMux I__3259 (
            .O(N__24249),
            .I(N__24241));
    Odrv4 I__3258 (
            .O(N__24246),
            .I(read_buf_6));
    LocalMux I__3257 (
            .O(N__24241),
            .I(read_buf_6));
    CascadeMux I__3256 (
            .O(N__24236),
            .I(N__24230));
    CascadeMux I__3255 (
            .O(N__24235),
            .I(N__24224));
    InMux I__3254 (
            .O(N__24234),
            .I(N__24213));
    InMux I__3253 (
            .O(N__24233),
            .I(N__24213));
    InMux I__3252 (
            .O(N__24230),
            .I(N__24208));
    InMux I__3251 (
            .O(N__24229),
            .I(N__24208));
    InMux I__3250 (
            .O(N__24228),
            .I(N__24203));
    InMux I__3249 (
            .O(N__24227),
            .I(N__24203));
    InMux I__3248 (
            .O(N__24224),
            .I(N__24194));
    InMux I__3247 (
            .O(N__24223),
            .I(N__24194));
    InMux I__3246 (
            .O(N__24222),
            .I(N__24194));
    InMux I__3245 (
            .O(N__24221),
            .I(N__24185));
    InMux I__3244 (
            .O(N__24220),
            .I(N__24185));
    InMux I__3243 (
            .O(N__24219),
            .I(N__24185));
    InMux I__3242 (
            .O(N__24218),
            .I(N__24185));
    LocalMux I__3241 (
            .O(N__24213),
            .I(N__24182));
    LocalMux I__3240 (
            .O(N__24208),
            .I(N__24179));
    LocalMux I__3239 (
            .O(N__24203),
            .I(N__24176));
    InMux I__3238 (
            .O(N__24202),
            .I(N__24173));
    InMux I__3237 (
            .O(N__24201),
            .I(N__24170));
    LocalMux I__3236 (
            .O(N__24194),
            .I(N__24167));
    LocalMux I__3235 (
            .O(N__24185),
            .I(N__24164));
    Span4Mux_h I__3234 (
            .O(N__24182),
            .I(N__24161));
    Span4Mux_v I__3233 (
            .O(N__24179),
            .I(N__24156));
    Span4Mux_h I__3232 (
            .O(N__24176),
            .I(N__24156));
    LocalMux I__3231 (
            .O(N__24173),
            .I(n11730));
    LocalMux I__3230 (
            .O(N__24170),
            .I(n11730));
    Odrv4 I__3229 (
            .O(N__24167),
            .I(n11730));
    Odrv12 I__3228 (
            .O(N__24164),
            .I(n11730));
    Odrv4 I__3227 (
            .O(N__24161),
            .I(n11730));
    Odrv4 I__3226 (
            .O(N__24156),
            .I(n11730));
    InMux I__3225 (
            .O(N__24143),
            .I(N__24128));
    InMux I__3224 (
            .O(N__24142),
            .I(N__24128));
    InMux I__3223 (
            .O(N__24141),
            .I(N__24128));
    InMux I__3222 (
            .O(N__24140),
            .I(N__24128));
    InMux I__3221 (
            .O(N__24139),
            .I(N__24128));
    LocalMux I__3220 (
            .O(N__24128),
            .I(N__24122));
    InMux I__3219 (
            .O(N__24127),
            .I(N__24115));
    InMux I__3218 (
            .O(N__24126),
            .I(N__24115));
    InMux I__3217 (
            .O(N__24125),
            .I(N__24115));
    Odrv4 I__3216 (
            .O(N__24122),
            .I(\RTD.n13192 ));
    LocalMux I__3215 (
            .O(N__24115),
            .I(\RTD.n13192 ));
    InMux I__3214 (
            .O(N__24110),
            .I(N__24091));
    InMux I__3213 (
            .O(N__24109),
            .I(N__24091));
    InMux I__3212 (
            .O(N__24108),
            .I(N__24091));
    InMux I__3211 (
            .O(N__24107),
            .I(N__24091));
    InMux I__3210 (
            .O(N__24106),
            .I(N__24091));
    InMux I__3209 (
            .O(N__24105),
            .I(N__24084));
    InMux I__3208 (
            .O(N__24104),
            .I(N__24084));
    InMux I__3207 (
            .O(N__24103),
            .I(N__24084));
    CascadeMux I__3206 (
            .O(N__24102),
            .I(N__24081));
    LocalMux I__3205 (
            .O(N__24091),
            .I(N__24078));
    LocalMux I__3204 (
            .O(N__24084),
            .I(N__24075));
    InMux I__3203 (
            .O(N__24081),
            .I(N__24072));
    Odrv4 I__3202 (
            .O(N__24078),
            .I(\RTD.n20631 ));
    Odrv4 I__3201 (
            .O(N__24075),
            .I(\RTD.n20631 ));
    LocalMux I__3200 (
            .O(N__24072),
            .I(\RTD.n20631 ));
    InMux I__3199 (
            .O(N__24065),
            .I(N__24059));
    InMux I__3198 (
            .O(N__24064),
            .I(N__24056));
    InMux I__3197 (
            .O(N__24063),
            .I(N__24051));
    InMux I__3196 (
            .O(N__24062),
            .I(N__24051));
    LocalMux I__3195 (
            .O(N__24059),
            .I(N__24048));
    LocalMux I__3194 (
            .O(N__24056),
            .I(N__24042));
    LocalMux I__3193 (
            .O(N__24051),
            .I(N__24042));
    Span12Mux_v I__3192 (
            .O(N__24048),
            .I(N__24039));
    InMux I__3191 (
            .O(N__24047),
            .I(N__24036));
    Span4Mux_v I__3190 (
            .O(N__24042),
            .I(N__24033));
    Odrv12 I__3189 (
            .O(N__24039),
            .I(buf_cfgRTD_7));
    LocalMux I__3188 (
            .O(N__24036),
            .I(buf_cfgRTD_7));
    Odrv4 I__3187 (
            .O(N__24033),
            .I(buf_cfgRTD_7));
    CascadeMux I__3186 (
            .O(N__24026),
            .I(N__24023));
    InMux I__3185 (
            .O(N__24023),
            .I(N__24019));
    InMux I__3184 (
            .O(N__24022),
            .I(N__24016));
    LocalMux I__3183 (
            .O(N__24019),
            .I(\RTD.cfg_buf_7 ));
    LocalMux I__3182 (
            .O(N__24016),
            .I(\RTD.cfg_buf_7 ));
    InMux I__3181 (
            .O(N__24011),
            .I(N__24008));
    LocalMux I__3180 (
            .O(N__24008),
            .I(N__24005));
    Odrv12 I__3179 (
            .O(N__24005),
            .I(\ADC_VDC.n18479 ));
    CascadeMux I__3178 (
            .O(N__24002),
            .I(\ADC_VDC.n21145_cascade_ ));
    CEMux I__3177 (
            .O(N__23999),
            .I(N__23996));
    LocalMux I__3176 (
            .O(N__23996),
            .I(N__23993));
    Odrv4 I__3175 (
            .O(N__23993),
            .I(\ADC_VDC.n13050 ));
    CascadeMux I__3174 (
            .O(N__23990),
            .I(N__23987));
    InMux I__3173 (
            .O(N__23987),
            .I(N__23984));
    LocalMux I__3172 (
            .O(N__23984),
            .I(N__23981));
    Span4Mux_v I__3171 (
            .O(N__23981),
            .I(N__23978));
    Span4Mux_h I__3170 (
            .O(N__23978),
            .I(N__23973));
    InMux I__3169 (
            .O(N__23977),
            .I(N__23968));
    InMux I__3168 (
            .O(N__23976),
            .I(N__23968));
    Odrv4 I__3167 (
            .O(N__23973),
            .I(read_buf_10));
    LocalMux I__3166 (
            .O(N__23968),
            .I(read_buf_10));
    InMux I__3165 (
            .O(N__23963),
            .I(N__23960));
    LocalMux I__3164 (
            .O(N__23960),
            .I(N__23957));
    Span4Mux_v I__3163 (
            .O(N__23957),
            .I(N__23953));
    CascadeMux I__3162 (
            .O(N__23956),
            .I(N__23950));
    Span4Mux_v I__3161 (
            .O(N__23953),
            .I(N__23947));
    InMux I__3160 (
            .O(N__23950),
            .I(N__23944));
    Odrv4 I__3159 (
            .O(N__23947),
            .I(buf_adcdata_vdc_18));
    LocalMux I__3158 (
            .O(N__23944),
            .I(buf_adcdata_vdc_18));
    CascadeMux I__3157 (
            .O(N__23939),
            .I(n20833_cascade_));
    CascadeMux I__3156 (
            .O(N__23936),
            .I(N__23933));
    InMux I__3155 (
            .O(N__23933),
            .I(N__23930));
    LocalMux I__3154 (
            .O(N__23930),
            .I(N__23927));
    Span4Mux_h I__3153 (
            .O(N__23927),
            .I(N__23922));
    InMux I__3152 (
            .O(N__23926),
            .I(N__23917));
    InMux I__3151 (
            .O(N__23925),
            .I(N__23917));
    Odrv4 I__3150 (
            .O(N__23922),
            .I(read_buf_14));
    LocalMux I__3149 (
            .O(N__23917),
            .I(read_buf_14));
    CascadeMux I__3148 (
            .O(N__23912),
            .I(N__23909));
    InMux I__3147 (
            .O(N__23909),
            .I(N__23906));
    LocalMux I__3146 (
            .O(N__23906),
            .I(N__23903));
    Span4Mux_v I__3145 (
            .O(N__23903),
            .I(N__23899));
    InMux I__3144 (
            .O(N__23902),
            .I(N__23896));
    Odrv4 I__3143 (
            .O(N__23899),
            .I(buf_readRTD_11));
    LocalMux I__3142 (
            .O(N__23896),
            .I(buf_readRTD_11));
    InMux I__3141 (
            .O(N__23891),
            .I(N__23888));
    LocalMux I__3140 (
            .O(N__23888),
            .I(N__23885));
    Odrv4 I__3139 (
            .O(N__23885),
            .I(n22214));
    CascadeMux I__3138 (
            .O(N__23882),
            .I(N__23879));
    InMux I__3137 (
            .O(N__23879),
            .I(N__23876));
    LocalMux I__3136 (
            .O(N__23876),
            .I(N__23872));
    CascadeMux I__3135 (
            .O(N__23875),
            .I(N__23869));
    Span4Mux_h I__3134 (
            .O(N__23872),
            .I(N__23866));
    InMux I__3133 (
            .O(N__23869),
            .I(N__23863));
    Odrv4 I__3132 (
            .O(N__23866),
            .I(buf_adcdata_vdc_19));
    LocalMux I__3131 (
            .O(N__23863),
            .I(buf_adcdata_vdc_19));
    InMux I__3130 (
            .O(N__23858),
            .I(N__23855));
    LocalMux I__3129 (
            .O(N__23855),
            .I(N__23851));
    InMux I__3128 (
            .O(N__23854),
            .I(N__23848));
    Span4Mux_v I__3127 (
            .O(N__23851),
            .I(N__23845));
    LocalMux I__3126 (
            .O(N__23848),
            .I(\ADC_VDC.avg_cnt_11 ));
    Odrv4 I__3125 (
            .O(N__23845),
            .I(\ADC_VDC.avg_cnt_11 ));
    InMux I__3124 (
            .O(N__23840),
            .I(N__23837));
    LocalMux I__3123 (
            .O(N__23837),
            .I(N__23833));
    InMux I__3122 (
            .O(N__23836),
            .I(N__23830));
    Span4Mux_h I__3121 (
            .O(N__23833),
            .I(N__23827));
    LocalMux I__3120 (
            .O(N__23830),
            .I(\ADC_VDC.avg_cnt_2 ));
    Odrv4 I__3119 (
            .O(N__23827),
            .I(\ADC_VDC.avg_cnt_2 ));
    CascadeMux I__3118 (
            .O(N__23822),
            .I(N__23819));
    InMux I__3117 (
            .O(N__23819),
            .I(N__23816));
    LocalMux I__3116 (
            .O(N__23816),
            .I(N__23812));
    InMux I__3115 (
            .O(N__23815),
            .I(N__23809));
    Span4Mux_v I__3114 (
            .O(N__23812),
            .I(N__23806));
    LocalMux I__3113 (
            .O(N__23809),
            .I(\ADC_VDC.avg_cnt_1 ));
    Odrv4 I__3112 (
            .O(N__23806),
            .I(\ADC_VDC.avg_cnt_1 ));
    InMux I__3111 (
            .O(N__23801),
            .I(N__23798));
    LocalMux I__3110 (
            .O(N__23798),
            .I(N__23794));
    InMux I__3109 (
            .O(N__23797),
            .I(N__23791));
    Span4Mux_h I__3108 (
            .O(N__23794),
            .I(N__23788));
    LocalMux I__3107 (
            .O(N__23791),
            .I(\ADC_VDC.avg_cnt_6 ));
    Odrv4 I__3106 (
            .O(N__23788),
            .I(\ADC_VDC.avg_cnt_6 ));
    InMux I__3105 (
            .O(N__23783),
            .I(N__23780));
    LocalMux I__3104 (
            .O(N__23780),
            .I(N__23777));
    Odrv12 I__3103 (
            .O(N__23777),
            .I(\ADC_VDC.n21 ));
    CascadeMux I__3102 (
            .O(N__23774),
            .I(n12875_cascade_));
    InMux I__3101 (
            .O(N__23771),
            .I(N__23768));
    LocalMux I__3100 (
            .O(N__23768),
            .I(N__23763));
    InMux I__3099 (
            .O(N__23767),
            .I(N__23758));
    InMux I__3098 (
            .O(N__23766),
            .I(N__23758));
    Span12Mux_s9_v I__3097 (
            .O(N__23763),
            .I(N__23755));
    LocalMux I__3096 (
            .O(N__23758),
            .I(buf_adcdata_iac_6));
    Odrv12 I__3095 (
            .O(N__23755),
            .I(buf_adcdata_iac_6));
    CascadeMux I__3094 (
            .O(N__23750),
            .I(n19_adj_1628_cascade_));
    InMux I__3093 (
            .O(N__23747),
            .I(N__23744));
    LocalMux I__3092 (
            .O(N__23744),
            .I(N__23741));
    Span12Mux_h I__3091 (
            .O(N__23741),
            .I(N__23738));
    Odrv12 I__3090 (
            .O(N__23738),
            .I(buf_data_iac_6));
    CascadeMux I__3089 (
            .O(N__23735),
            .I(n22_adj_1629_cascade_));
    CascadeMux I__3088 (
            .O(N__23732),
            .I(N__23728));
    InMux I__3087 (
            .O(N__23731),
            .I(N__23720));
    InMux I__3086 (
            .O(N__23728),
            .I(N__23720));
    InMux I__3085 (
            .O(N__23727),
            .I(N__23720));
    LocalMux I__3084 (
            .O(N__23720),
            .I(cmd_rdadctmp_14_adj_1436));
    CascadeMux I__3083 (
            .O(N__23717),
            .I(N__23713));
    CascadeMux I__3082 (
            .O(N__23716),
            .I(N__23710));
    InMux I__3081 (
            .O(N__23713),
            .I(N__23706));
    InMux I__3080 (
            .O(N__23710),
            .I(N__23701));
    InMux I__3079 (
            .O(N__23709),
            .I(N__23701));
    LocalMux I__3078 (
            .O(N__23706),
            .I(cmd_rdadctmp_15_adj_1435));
    LocalMux I__3077 (
            .O(N__23701),
            .I(cmd_rdadctmp_15_adj_1435));
    CascadeMux I__3076 (
            .O(N__23696),
            .I(N__23692));
    InMux I__3075 (
            .O(N__23695),
            .I(N__23687));
    InMux I__3074 (
            .O(N__23692),
            .I(N__23687));
    LocalMux I__3073 (
            .O(N__23687),
            .I(N__23683));
    InMux I__3072 (
            .O(N__23686),
            .I(N__23680));
    Odrv4 I__3071 (
            .O(N__23683),
            .I(cmd_rdadctmp_14));
    LocalMux I__3070 (
            .O(N__23680),
            .I(cmd_rdadctmp_14));
    InMux I__3069 (
            .O(N__23675),
            .I(N__23672));
    LocalMux I__3068 (
            .O(N__23672),
            .I(N__23668));
    CascadeMux I__3067 (
            .O(N__23671),
            .I(N__23665));
    Span4Mux_h I__3066 (
            .O(N__23668),
            .I(N__23662));
    InMux I__3065 (
            .O(N__23665),
            .I(N__23659));
    Odrv4 I__3064 (
            .O(N__23662),
            .I(buf_adcdata_vdc_7));
    LocalMux I__3063 (
            .O(N__23659),
            .I(buf_adcdata_vdc_7));
    InMux I__3062 (
            .O(N__23654),
            .I(N__23651));
    LocalMux I__3061 (
            .O(N__23651),
            .I(N__23647));
    InMux I__3060 (
            .O(N__23650),
            .I(N__23643));
    Span4Mux_h I__3059 (
            .O(N__23647),
            .I(N__23640));
    InMux I__3058 (
            .O(N__23646),
            .I(N__23637));
    LocalMux I__3057 (
            .O(N__23643),
            .I(buf_adcdata_vac_7));
    Odrv4 I__3056 (
            .O(N__23640),
            .I(buf_adcdata_vac_7));
    LocalMux I__3055 (
            .O(N__23637),
            .I(buf_adcdata_vac_7));
    InMux I__3054 (
            .O(N__23630),
            .I(N__23627));
    LocalMux I__3053 (
            .O(N__23627),
            .I(N__23624));
    Span12Mux_s8_v I__3052 (
            .O(N__23624),
            .I(N__23619));
    InMux I__3051 (
            .O(N__23623),
            .I(N__23614));
    InMux I__3050 (
            .O(N__23622),
            .I(N__23614));
    Odrv12 I__3049 (
            .O(N__23619),
            .I(buf_adcdata_iac_7));
    LocalMux I__3048 (
            .O(N__23614),
            .I(buf_adcdata_iac_7));
    CascadeMux I__3047 (
            .O(N__23609),
            .I(n19_adj_1625_cascade_));
    InMux I__3046 (
            .O(N__23606),
            .I(N__23603));
    LocalMux I__3045 (
            .O(N__23603),
            .I(N__23600));
    Span12Mux_h I__3044 (
            .O(N__23600),
            .I(N__23597));
    Odrv12 I__3043 (
            .O(N__23597),
            .I(buf_data_iac_7));
    CascadeMux I__3042 (
            .O(N__23594),
            .I(n22_adj_1626_cascade_));
    InMux I__3041 (
            .O(N__23591),
            .I(N__23587));
    CascadeMux I__3040 (
            .O(N__23590),
            .I(N__23584));
    LocalMux I__3039 (
            .O(N__23587),
            .I(N__23580));
    InMux I__3038 (
            .O(N__23584),
            .I(N__23577));
    InMux I__3037 (
            .O(N__23583),
            .I(N__23574));
    Span4Mux_h I__3036 (
            .O(N__23580),
            .I(N__23571));
    LocalMux I__3035 (
            .O(N__23577),
            .I(buf_adcdata_vac_6));
    LocalMux I__3034 (
            .O(N__23574),
            .I(buf_adcdata_vac_6));
    Odrv4 I__3033 (
            .O(N__23571),
            .I(buf_adcdata_vac_6));
    InMux I__3032 (
            .O(N__23564),
            .I(N__23561));
    LocalMux I__3031 (
            .O(N__23561),
            .I(N__23558));
    Span4Mux_v I__3030 (
            .O(N__23558),
            .I(N__23554));
    InMux I__3029 (
            .O(N__23557),
            .I(N__23551));
    Odrv4 I__3028 (
            .O(N__23554),
            .I(buf_adcdata_vdc_6));
    LocalMux I__3027 (
            .O(N__23551),
            .I(buf_adcdata_vdc_6));
    CascadeMux I__3026 (
            .O(N__23546),
            .I(N__23543));
    InMux I__3025 (
            .O(N__23543),
            .I(N__23540));
    LocalMux I__3024 (
            .O(N__23540),
            .I(\CLK_DDS.tmp_buf_14 ));
    CascadeMux I__3023 (
            .O(N__23537),
            .I(N__23534));
    InMux I__3022 (
            .O(N__23534),
            .I(N__23530));
    InMux I__3021 (
            .O(N__23533),
            .I(N__23527));
    LocalMux I__3020 (
            .O(N__23530),
            .I(N__23524));
    LocalMux I__3019 (
            .O(N__23527),
            .I(N__23519));
    Span4Mux_h I__3018 (
            .O(N__23524),
            .I(N__23519));
    Span4Mux_v I__3017 (
            .O(N__23519),
            .I(N__23516));
    Odrv4 I__3016 (
            .O(N__23516),
            .I(tmp_buf_15_adj_1455));
    CascadeMux I__3015 (
            .O(N__23513),
            .I(N__23500));
    CascadeMux I__3014 (
            .O(N__23512),
            .I(N__23491));
    InMux I__3013 (
            .O(N__23511),
            .I(N__23485));
    InMux I__3012 (
            .O(N__23510),
            .I(N__23480));
    InMux I__3011 (
            .O(N__23509),
            .I(N__23465));
    InMux I__3010 (
            .O(N__23508),
            .I(N__23465));
    InMux I__3009 (
            .O(N__23507),
            .I(N__23465));
    InMux I__3008 (
            .O(N__23506),
            .I(N__23465));
    InMux I__3007 (
            .O(N__23505),
            .I(N__23465));
    InMux I__3006 (
            .O(N__23504),
            .I(N__23465));
    InMux I__3005 (
            .O(N__23503),
            .I(N__23465));
    InMux I__3004 (
            .O(N__23500),
            .I(N__23460));
    InMux I__3003 (
            .O(N__23499),
            .I(N__23460));
    InMux I__3002 (
            .O(N__23498),
            .I(N__23451));
    InMux I__3001 (
            .O(N__23497),
            .I(N__23451));
    InMux I__3000 (
            .O(N__23496),
            .I(N__23451));
    InMux I__2999 (
            .O(N__23495),
            .I(N__23451));
    InMux I__2998 (
            .O(N__23494),
            .I(N__23444));
    InMux I__2997 (
            .O(N__23491),
            .I(N__23444));
    InMux I__2996 (
            .O(N__23490),
            .I(N__23444));
    InMux I__2995 (
            .O(N__23489),
            .I(N__23441));
    InMux I__2994 (
            .O(N__23488),
            .I(N__23437));
    LocalMux I__2993 (
            .O(N__23485),
            .I(N__23434));
    InMux I__2992 (
            .O(N__23484),
            .I(N__23431));
    InMux I__2991 (
            .O(N__23483),
            .I(N__23428));
    LocalMux I__2990 (
            .O(N__23480),
            .I(N__23425));
    LocalMux I__2989 (
            .O(N__23465),
            .I(N__23422));
    LocalMux I__2988 (
            .O(N__23460),
            .I(N__23412));
    LocalMux I__2987 (
            .O(N__23451),
            .I(N__23412));
    LocalMux I__2986 (
            .O(N__23444),
            .I(N__23412));
    LocalMux I__2985 (
            .O(N__23441),
            .I(N__23412));
    InMux I__2984 (
            .O(N__23440),
            .I(N__23409));
    LocalMux I__2983 (
            .O(N__23437),
            .I(N__23406));
    Span4Mux_h I__2982 (
            .O(N__23434),
            .I(N__23403));
    LocalMux I__2981 (
            .O(N__23431),
            .I(N__23394));
    LocalMux I__2980 (
            .O(N__23428),
            .I(N__23394));
    Span4Mux_v I__2979 (
            .O(N__23425),
            .I(N__23394));
    Span4Mux_h I__2978 (
            .O(N__23422),
            .I(N__23394));
    InMux I__2977 (
            .O(N__23421),
            .I(N__23389));
    Span4Mux_v I__2976 (
            .O(N__23412),
            .I(N__23386));
    LocalMux I__2975 (
            .O(N__23409),
            .I(N__23377));
    Span4Mux_v I__2974 (
            .O(N__23406),
            .I(N__23377));
    Span4Mux_v I__2973 (
            .O(N__23403),
            .I(N__23377));
    Span4Mux_v I__2972 (
            .O(N__23394),
            .I(N__23377));
    InMux I__2971 (
            .O(N__23393),
            .I(N__23372));
    InMux I__2970 (
            .O(N__23392),
            .I(N__23372));
    LocalMux I__2969 (
            .O(N__23389),
            .I(N__23367));
    Span4Mux_h I__2968 (
            .O(N__23386),
            .I(N__23367));
    Odrv4 I__2967 (
            .O(N__23377),
            .I(dds_state_2_adj_1452));
    LocalMux I__2966 (
            .O(N__23372),
            .I(dds_state_2_adj_1452));
    Odrv4 I__2965 (
            .O(N__23367),
            .I(dds_state_2_adj_1452));
    CascadeMux I__2964 (
            .O(N__23360),
            .I(N__23354));
    SRMux I__2963 (
            .O(N__23359),
            .I(N__23349));
    InMux I__2962 (
            .O(N__23358),
            .I(N__23346));
    CEMux I__2961 (
            .O(N__23357),
            .I(N__23343));
    InMux I__2960 (
            .O(N__23354),
            .I(N__23328));
    CascadeMux I__2959 (
            .O(N__23353),
            .I(N__23320));
    InMux I__2958 (
            .O(N__23352),
            .I(N__23313));
    LocalMux I__2957 (
            .O(N__23349),
            .I(N__23310));
    LocalMux I__2956 (
            .O(N__23346),
            .I(N__23305));
    LocalMux I__2955 (
            .O(N__23343),
            .I(N__23305));
    InMux I__2954 (
            .O(N__23342),
            .I(N__23302));
    InMux I__2953 (
            .O(N__23341),
            .I(N__23287));
    InMux I__2952 (
            .O(N__23340),
            .I(N__23287));
    InMux I__2951 (
            .O(N__23339),
            .I(N__23287));
    InMux I__2950 (
            .O(N__23338),
            .I(N__23287));
    InMux I__2949 (
            .O(N__23337),
            .I(N__23287));
    InMux I__2948 (
            .O(N__23336),
            .I(N__23287));
    InMux I__2947 (
            .O(N__23335),
            .I(N__23287));
    InMux I__2946 (
            .O(N__23334),
            .I(N__23278));
    InMux I__2945 (
            .O(N__23333),
            .I(N__23278));
    InMux I__2944 (
            .O(N__23332),
            .I(N__23278));
    InMux I__2943 (
            .O(N__23331),
            .I(N__23278));
    LocalMux I__2942 (
            .O(N__23328),
            .I(N__23275));
    InMux I__2941 (
            .O(N__23327),
            .I(N__23264));
    InMux I__2940 (
            .O(N__23326),
            .I(N__23264));
    InMux I__2939 (
            .O(N__23325),
            .I(N__23264));
    InMux I__2938 (
            .O(N__23324),
            .I(N__23264));
    InMux I__2937 (
            .O(N__23323),
            .I(N__23264));
    InMux I__2936 (
            .O(N__23320),
            .I(N__23261));
    InMux I__2935 (
            .O(N__23319),
            .I(N__23258));
    InMux I__2934 (
            .O(N__23318),
            .I(N__23255));
    InMux I__2933 (
            .O(N__23317),
            .I(N__23252));
    InMux I__2932 (
            .O(N__23316),
            .I(N__23249));
    LocalMux I__2931 (
            .O(N__23313),
            .I(N__23246));
    Span4Mux_h I__2930 (
            .O(N__23310),
            .I(N__23243));
    Span4Mux_v I__2929 (
            .O(N__23305),
            .I(N__23240));
    LocalMux I__2928 (
            .O(N__23302),
            .I(N__23229));
    LocalMux I__2927 (
            .O(N__23287),
            .I(N__23229));
    LocalMux I__2926 (
            .O(N__23278),
            .I(N__23229));
    Span4Mux_v I__2925 (
            .O(N__23275),
            .I(N__23229));
    LocalMux I__2924 (
            .O(N__23264),
            .I(N__23229));
    LocalMux I__2923 (
            .O(N__23261),
            .I(N__23217));
    LocalMux I__2922 (
            .O(N__23258),
            .I(N__23217));
    LocalMux I__2921 (
            .O(N__23255),
            .I(N__23217));
    LocalMux I__2920 (
            .O(N__23252),
            .I(N__23217));
    LocalMux I__2919 (
            .O(N__23249),
            .I(N__23217));
    Span4Mux_h I__2918 (
            .O(N__23246),
            .I(N__23214));
    Span4Mux_h I__2917 (
            .O(N__23243),
            .I(N__23207));
    Span4Mux_v I__2916 (
            .O(N__23240),
            .I(N__23207));
    Span4Mux_v I__2915 (
            .O(N__23229),
            .I(N__23207));
    InMux I__2914 (
            .O(N__23228),
            .I(N__23204));
    Odrv12 I__2913 (
            .O(N__23217),
            .I(dds_state_1_adj_1453));
    Odrv4 I__2912 (
            .O(N__23214),
            .I(dds_state_1_adj_1453));
    Odrv4 I__2911 (
            .O(N__23207),
            .I(dds_state_1_adj_1453));
    LocalMux I__2910 (
            .O(N__23204),
            .I(dds_state_1_adj_1453));
    CascadeMux I__2909 (
            .O(N__23195),
            .I(N__23192));
    InMux I__2908 (
            .O(N__23192),
            .I(N__23189));
    LocalMux I__2907 (
            .O(N__23189),
            .I(\CLK_DDS.tmp_buf_8 ));
    CascadeMux I__2906 (
            .O(N__23186),
            .I(N__23183));
    InMux I__2905 (
            .O(N__23183),
            .I(N__23180));
    LocalMux I__2904 (
            .O(N__23180),
            .I(\CLK_DDS.tmp_buf_9 ));
    CEMux I__2903 (
            .O(N__23177),
            .I(N__23174));
    LocalMux I__2902 (
            .O(N__23174),
            .I(N__23171));
    Span4Mux_h I__2901 (
            .O(N__23171),
            .I(N__23166));
    CEMux I__2900 (
            .O(N__23170),
            .I(N__23163));
    CEMux I__2899 (
            .O(N__23169),
            .I(N__23160));
    Span4Mux_v I__2898 (
            .O(N__23166),
            .I(N__23155));
    LocalMux I__2897 (
            .O(N__23163),
            .I(N__23155));
    LocalMux I__2896 (
            .O(N__23160),
            .I(N__23152));
    Span4Mux_h I__2895 (
            .O(N__23155),
            .I(N__23149));
    Span4Mux_h I__2894 (
            .O(N__23152),
            .I(N__23146));
    Span4Mux_v I__2893 (
            .O(N__23149),
            .I(N__23139));
    Span4Mux_h I__2892 (
            .O(N__23146),
            .I(N__23139));
    CEMux I__2891 (
            .O(N__23145),
            .I(N__23136));
    CEMux I__2890 (
            .O(N__23144),
            .I(N__23133));
    Odrv4 I__2889 (
            .O(N__23139),
            .I(\CLK_DDS.n12800 ));
    LocalMux I__2888 (
            .O(N__23136),
            .I(\CLK_DDS.n12800 ));
    LocalMux I__2887 (
            .O(N__23133),
            .I(\CLK_DDS.n12800 ));
    CascadeMux I__2886 (
            .O(N__23126),
            .I(N__23122));
    CascadeMux I__2885 (
            .O(N__23125),
            .I(N__23118));
    InMux I__2884 (
            .O(N__23122),
            .I(N__23115));
    CascadeMux I__2883 (
            .O(N__23121),
            .I(N__23111));
    InMux I__2882 (
            .O(N__23118),
            .I(N__23108));
    LocalMux I__2881 (
            .O(N__23115),
            .I(N__23105));
    InMux I__2880 (
            .O(N__23114),
            .I(N__23100));
    InMux I__2879 (
            .O(N__23111),
            .I(N__23100));
    LocalMux I__2878 (
            .O(N__23108),
            .I(trig_dds1));
    Odrv4 I__2877 (
            .O(N__23105),
            .I(trig_dds1));
    LocalMux I__2876 (
            .O(N__23100),
            .I(trig_dds1));
    InMux I__2875 (
            .O(N__23093),
            .I(N__23090));
    LocalMux I__2874 (
            .O(N__23090),
            .I(N__23087));
    Span4Mux_v I__2873 (
            .O(N__23087),
            .I(N__23084));
    Sp12to4 I__2872 (
            .O(N__23084),
            .I(N__23081));
    Span12Mux_h I__2871 (
            .O(N__23081),
            .I(N__23078));
    Odrv12 I__2870 (
            .O(N__23078),
            .I(ICE_GPMO_1));
    IoInMux I__2869 (
            .O(N__23075),
            .I(N__23072));
    LocalMux I__2868 (
            .O(N__23072),
            .I(N__23069));
    IoSpan4Mux I__2867 (
            .O(N__23069),
            .I(N__23065));
    IoInMux I__2866 (
            .O(N__23068),
            .I(N__23062));
    IoSpan4Mux I__2865 (
            .O(N__23065),
            .I(N__23059));
    LocalMux I__2864 (
            .O(N__23062),
            .I(N__23056));
    Span4Mux_s2_v I__2863 (
            .O(N__23059),
            .I(N__23053));
    IoSpan4Mux I__2862 (
            .O(N__23056),
            .I(N__23050));
    Span4Mux_v I__2861 (
            .O(N__23053),
            .I(N__23047));
    Sp12to4 I__2860 (
            .O(N__23050),
            .I(N__23044));
    Sp12to4 I__2859 (
            .O(N__23047),
            .I(N__23039));
    Span12Mux_h I__2858 (
            .O(N__23044),
            .I(N__23039));
    Span12Mux_v I__2857 (
            .O(N__23039),
            .I(N__23036));
    Odrv12 I__2856 (
            .O(N__23036),
            .I(IAC_CLK));
    CascadeMux I__2855 (
            .O(N__23033),
            .I(N__23030));
    InMux I__2854 (
            .O(N__23030),
            .I(N__23027));
    LocalMux I__2853 (
            .O(N__23027),
            .I(n22100));
    IoInMux I__2852 (
            .O(N__23024),
            .I(N__23021));
    LocalMux I__2851 (
            .O(N__23021),
            .I(N__23018));
    IoSpan4Mux I__2850 (
            .O(N__23018),
            .I(N__23015));
    Span4Mux_s0_v I__2849 (
            .O(N__23015),
            .I(N__23012));
    Sp12to4 I__2848 (
            .O(N__23012),
            .I(N__23008));
    InMux I__2847 (
            .O(N__23011),
            .I(N__23004));
    Span12Mux_v I__2846 (
            .O(N__23008),
            .I(N__23001));
    InMux I__2845 (
            .O(N__23007),
            .I(N__22998));
    LocalMux I__2844 (
            .O(N__23004),
            .I(N__22995));
    Odrv12 I__2843 (
            .O(N__23001),
            .I(SELIRNG0));
    LocalMux I__2842 (
            .O(N__22998),
            .I(SELIRNG0));
    Odrv4 I__2841 (
            .O(N__22995),
            .I(SELIRNG0));
    CascadeMux I__2840 (
            .O(N__22988),
            .I(N__22985));
    InMux I__2839 (
            .O(N__22985),
            .I(N__22982));
    LocalMux I__2838 (
            .O(N__22982),
            .I(\CLK_DDS.tmp_buf_10 ));
    CascadeMux I__2837 (
            .O(N__22979),
            .I(N__22976));
    InMux I__2836 (
            .O(N__22976),
            .I(N__22973));
    LocalMux I__2835 (
            .O(N__22973),
            .I(\CLK_DDS.tmp_buf_11 ));
    CascadeMux I__2834 (
            .O(N__22970),
            .I(N__22967));
    InMux I__2833 (
            .O(N__22967),
            .I(N__22964));
    LocalMux I__2832 (
            .O(N__22964),
            .I(\CLK_DDS.tmp_buf_12 ));
    InMux I__2831 (
            .O(N__22961),
            .I(N__22958));
    LocalMux I__2830 (
            .O(N__22958),
            .I(\CLK_DDS.tmp_buf_13 ));
    CascadeMux I__2829 (
            .O(N__22955),
            .I(N__22951));
    CascadeMux I__2828 (
            .O(N__22954),
            .I(N__22947));
    InMux I__2827 (
            .O(N__22951),
            .I(N__22944));
    InMux I__2826 (
            .O(N__22950),
            .I(N__22941));
    InMux I__2825 (
            .O(N__22947),
            .I(N__22938));
    LocalMux I__2824 (
            .O(N__22944),
            .I(cmd_rdadctmp_25_adj_1425));
    LocalMux I__2823 (
            .O(N__22941),
            .I(cmd_rdadctmp_25_adj_1425));
    LocalMux I__2822 (
            .O(N__22938),
            .I(cmd_rdadctmp_25_adj_1425));
    CascadeMux I__2821 (
            .O(N__22931),
            .I(N__22927));
    CascadeMux I__2820 (
            .O(N__22930),
            .I(N__22924));
    InMux I__2819 (
            .O(N__22927),
            .I(N__22921));
    InMux I__2818 (
            .O(N__22924),
            .I(N__22918));
    LocalMux I__2817 (
            .O(N__22921),
            .I(cmd_rdadctmp_31_adj_1419));
    LocalMux I__2816 (
            .O(N__22918),
            .I(cmd_rdadctmp_31_adj_1419));
    IoInMux I__2815 (
            .O(N__22913),
            .I(N__22910));
    LocalMux I__2814 (
            .O(N__22910),
            .I(N__22907));
    Span12Mux_s11_h I__2813 (
            .O(N__22907),
            .I(N__22902));
    InMux I__2812 (
            .O(N__22906),
            .I(N__22897));
    InMux I__2811 (
            .O(N__22905),
            .I(N__22897));
    Odrv12 I__2810 (
            .O(N__22902),
            .I(VAC_OSR1));
    LocalMux I__2809 (
            .O(N__22897),
            .I(VAC_OSR1));
    InMux I__2808 (
            .O(N__22892),
            .I(N__22889));
    LocalMux I__2807 (
            .O(N__22889),
            .I(N__22886));
    Span4Mux_v I__2806 (
            .O(N__22886),
            .I(N__22883));
    Sp12to4 I__2805 (
            .O(N__22883),
            .I(N__22878));
    CascadeMux I__2804 (
            .O(N__22882),
            .I(N__22875));
    InMux I__2803 (
            .O(N__22881),
            .I(N__22872));
    Span12Mux_h I__2802 (
            .O(N__22878),
            .I(N__22869));
    InMux I__2801 (
            .O(N__22875),
            .I(N__22866));
    LocalMux I__2800 (
            .O(N__22872),
            .I(buf_adcdata_iac_21));
    Odrv12 I__2799 (
            .O(N__22869),
            .I(buf_adcdata_iac_21));
    LocalMux I__2798 (
            .O(N__22866),
            .I(buf_adcdata_iac_21));
    InMux I__2797 (
            .O(N__22859),
            .I(N__22856));
    LocalMux I__2796 (
            .O(N__22856),
            .I(N__22853));
    Span12Mux_h I__2795 (
            .O(N__22853),
            .I(N__22850));
    Span12Mux_v I__2794 (
            .O(N__22850),
            .I(N__22845));
    InMux I__2793 (
            .O(N__22849),
            .I(N__22840));
    InMux I__2792 (
            .O(N__22848),
            .I(N__22840));
    Odrv12 I__2791 (
            .O(N__22845),
            .I(buf_adcdata_iac_23));
    LocalMux I__2790 (
            .O(N__22840),
            .I(buf_adcdata_iac_23));
    IoInMux I__2789 (
            .O(N__22835),
            .I(N__22832));
    LocalMux I__2788 (
            .O(N__22832),
            .I(N__22829));
    IoSpan4Mux I__2787 (
            .O(N__22829),
            .I(N__22826));
    Span4Mux_s0_h I__2786 (
            .O(N__22826),
            .I(N__22823));
    Sp12to4 I__2785 (
            .O(N__22823),
            .I(N__22820));
    Span12Mux_s11_h I__2784 (
            .O(N__22820),
            .I(N__22815));
    InMux I__2783 (
            .O(N__22819),
            .I(N__22810));
    InMux I__2782 (
            .O(N__22818),
            .I(N__22810));
    Odrv12 I__2781 (
            .O(N__22815),
            .I(VAC_FLT1));
    LocalMux I__2780 (
            .O(N__22810),
            .I(VAC_FLT1));
    InMux I__2779 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__2778 (
            .O(N__22802),
            .I(N__22799));
    Span4Mux_v I__2777 (
            .O(N__22799),
            .I(N__22796));
    Odrv4 I__2776 (
            .O(N__22796),
            .I(n17_adj_1525));
    InMux I__2775 (
            .O(N__22793),
            .I(N__22790));
    LocalMux I__2774 (
            .O(N__22790),
            .I(N__22787));
    Span4Mux_v I__2773 (
            .O(N__22787),
            .I(N__22784));
    Sp12to4 I__2772 (
            .O(N__22784),
            .I(N__22779));
    CascadeMux I__2771 (
            .O(N__22783),
            .I(N__22776));
    InMux I__2770 (
            .O(N__22782),
            .I(N__22773));
    Span12Mux_h I__2769 (
            .O(N__22779),
            .I(N__22770));
    InMux I__2768 (
            .O(N__22776),
            .I(N__22767));
    LocalMux I__2767 (
            .O(N__22773),
            .I(buf_adcdata_iac_16));
    Odrv12 I__2766 (
            .O(N__22770),
            .I(buf_adcdata_iac_16));
    LocalMux I__2765 (
            .O(N__22767),
            .I(buf_adcdata_iac_16));
    IoInMux I__2764 (
            .O(N__22760),
            .I(N__22757));
    LocalMux I__2763 (
            .O(N__22757),
            .I(N__22754));
    Span4Mux_s2_v I__2762 (
            .O(N__22754),
            .I(N__22751));
    Span4Mux_h I__2761 (
            .O(N__22751),
            .I(N__22748));
    Span4Mux_h I__2760 (
            .O(N__22748),
            .I(N__22745));
    Sp12to4 I__2759 (
            .O(N__22745),
            .I(N__22740));
    InMux I__2758 (
            .O(N__22744),
            .I(N__22735));
    InMux I__2757 (
            .O(N__22743),
            .I(N__22735));
    Odrv12 I__2756 (
            .O(N__22740),
            .I(IAC_OSR0));
    LocalMux I__2755 (
            .O(N__22735),
            .I(IAC_OSR0));
    CascadeMux I__2754 (
            .O(N__22730),
            .I(\RTD.n21276_cascade_ ));
    InMux I__2753 (
            .O(N__22727),
            .I(N__22724));
    LocalMux I__2752 (
            .O(N__22724),
            .I(\RTD.n21275 ));
    InMux I__2751 (
            .O(N__22721),
            .I(N__22717));
    InMux I__2750 (
            .O(N__22720),
            .I(N__22714));
    LocalMux I__2749 (
            .O(N__22717),
            .I(\RTD.adc_state_3_N_1368_1 ));
    LocalMux I__2748 (
            .O(N__22714),
            .I(\RTD.adc_state_3_N_1368_1 ));
    CascadeMux I__2747 (
            .O(N__22709),
            .I(\RTD.adc_state_3_N_1368_1_cascade_ ));
    InMux I__2746 (
            .O(N__22706),
            .I(N__22703));
    LocalMux I__2745 (
            .O(N__22703),
            .I(\RTD.n7 ));
    CascadeMux I__2744 (
            .O(N__22700),
            .I(N__22697));
    InMux I__2743 (
            .O(N__22697),
            .I(N__22694));
    LocalMux I__2742 (
            .O(N__22694),
            .I(N__22691));
    Span4Mux_h I__2741 (
            .O(N__22691),
            .I(N__22688));
    Odrv4 I__2740 (
            .O(N__22688),
            .I(\RTD.n20762 ));
    CEMux I__2739 (
            .O(N__22685),
            .I(N__22680));
    CEMux I__2738 (
            .O(N__22684),
            .I(N__22677));
    CEMux I__2737 (
            .O(N__22683),
            .I(N__22674));
    LocalMux I__2736 (
            .O(N__22680),
            .I(N__22671));
    LocalMux I__2735 (
            .O(N__22677),
            .I(N__22668));
    LocalMux I__2734 (
            .O(N__22674),
            .I(N__22665));
    Odrv4 I__2733 (
            .O(N__22671),
            .I(\RTD.n11742 ));
    Odrv4 I__2732 (
            .O(N__22668),
            .I(\RTD.n11742 ));
    Odrv4 I__2731 (
            .O(N__22665),
            .I(\RTD.n11742 ));
    CascadeMux I__2730 (
            .O(N__22658),
            .I(n16_adj_1512_cascade_));
    CascadeMux I__2729 (
            .O(N__22655),
            .I(\RTD.n21323_cascade_ ));
    InMux I__2728 (
            .O(N__22652),
            .I(N__22649));
    LocalMux I__2727 (
            .O(N__22649),
            .I(\RTD.n26 ));
    CascadeMux I__2726 (
            .O(N__22646),
            .I(\RTD.n21325_cascade_ ));
    InMux I__2725 (
            .O(N__22643),
            .I(N__22640));
    LocalMux I__2724 (
            .O(N__22640),
            .I(\RTD.n4 ));
    InMux I__2723 (
            .O(N__22637),
            .I(N__22634));
    LocalMux I__2722 (
            .O(N__22634),
            .I(N__22629));
    InMux I__2721 (
            .O(N__22633),
            .I(N__22624));
    InMux I__2720 (
            .O(N__22632),
            .I(N__22624));
    Odrv4 I__2719 (
            .O(N__22629),
            .I(\RTD.n1 ));
    LocalMux I__2718 (
            .O(N__22624),
            .I(\RTD.n1 ));
    CascadeMux I__2717 (
            .O(N__22619),
            .I(\RTD.n1_cascade_ ));
    InMux I__2716 (
            .O(N__22616),
            .I(N__22612));
    InMux I__2715 (
            .O(N__22615),
            .I(N__22609));
    LocalMux I__2714 (
            .O(N__22612),
            .I(\RTD.n20587 ));
    LocalMux I__2713 (
            .O(N__22609),
            .I(\RTD.n20587 ));
    InMux I__2712 (
            .O(N__22604),
            .I(N__22601));
    LocalMux I__2711 (
            .O(N__22601),
            .I(N__22598));
    Odrv12 I__2710 (
            .O(N__22598),
            .I(n8_adj_1608));
    InMux I__2709 (
            .O(N__22595),
            .I(N__22592));
    LocalMux I__2708 (
            .O(N__22592),
            .I(N__22589));
    Span4Mux_v I__2707 (
            .O(N__22589),
            .I(N__22586));
    Odrv4 I__2706 (
            .O(N__22586),
            .I(n21227));
    InMux I__2705 (
            .O(N__22583),
            .I(N__22577));
    InMux I__2704 (
            .O(N__22582),
            .I(N__22570));
    InMux I__2703 (
            .O(N__22581),
            .I(N__22567));
    InMux I__2702 (
            .O(N__22580),
            .I(N__22564));
    LocalMux I__2701 (
            .O(N__22577),
            .I(N__22561));
    InMux I__2700 (
            .O(N__22576),
            .I(N__22556));
    InMux I__2699 (
            .O(N__22575),
            .I(N__22556));
    InMux I__2698 (
            .O(N__22574),
            .I(N__22553));
    InMux I__2697 (
            .O(N__22573),
            .I(N__22550));
    LocalMux I__2696 (
            .O(N__22570),
            .I(N__22547));
    LocalMux I__2695 (
            .O(N__22567),
            .I(N__22544));
    LocalMux I__2694 (
            .O(N__22564),
            .I(N__22540));
    Span4Mux_v I__2693 (
            .O(N__22561),
            .I(N__22533));
    LocalMux I__2692 (
            .O(N__22556),
            .I(N__22533));
    LocalMux I__2691 (
            .O(N__22553),
            .I(N__22533));
    LocalMux I__2690 (
            .O(N__22550),
            .I(N__22529));
    Span4Mux_h I__2689 (
            .O(N__22547),
            .I(N__22524));
    Span4Mux_h I__2688 (
            .O(N__22544),
            .I(N__22524));
    InMux I__2687 (
            .O(N__22543),
            .I(N__22521));
    Span4Mux_h I__2686 (
            .O(N__22540),
            .I(N__22516));
    Span4Mux_h I__2685 (
            .O(N__22533),
            .I(N__22516));
    InMux I__2684 (
            .O(N__22532),
            .I(N__22513));
    Span4Mux_h I__2683 (
            .O(N__22529),
            .I(N__22508));
    Span4Mux_v I__2682 (
            .O(N__22524),
            .I(N__22508));
    LocalMux I__2681 (
            .O(N__22521),
            .I(N__22505));
    Span4Mux_v I__2680 (
            .O(N__22516),
            .I(N__22502));
    LocalMux I__2679 (
            .O(N__22513),
            .I(dds_state_0_adj_1454));
    Odrv4 I__2678 (
            .O(N__22508),
            .I(dds_state_0_adj_1454));
    Odrv12 I__2677 (
            .O(N__22505),
            .I(dds_state_0_adj_1454));
    Odrv4 I__2676 (
            .O(N__22502),
            .I(dds_state_0_adj_1454));
    CEMux I__2675 (
            .O(N__22493),
            .I(N__22489));
    CEMux I__2674 (
            .O(N__22492),
            .I(N__22486));
    LocalMux I__2673 (
            .O(N__22489),
            .I(N__22483));
    LocalMux I__2672 (
            .O(N__22486),
            .I(N__22480));
    Span4Mux_v I__2671 (
            .O(N__22483),
            .I(N__22477));
    Span4Mux_h I__2670 (
            .O(N__22480),
            .I(N__22474));
    Odrv4 I__2669 (
            .O(N__22477),
            .I(\CLK_DDS.n9 ));
    Odrv4 I__2668 (
            .O(N__22474),
            .I(\CLK_DDS.n9 ));
    CascadeMux I__2667 (
            .O(N__22469),
            .I(N__22465));
    CascadeMux I__2666 (
            .O(N__22468),
            .I(N__22462));
    InMux I__2665 (
            .O(N__22465),
            .I(N__22458));
    InMux I__2664 (
            .O(N__22462),
            .I(N__22455));
    CascadeMux I__2663 (
            .O(N__22461),
            .I(N__22451));
    LocalMux I__2662 (
            .O(N__22458),
            .I(N__22448));
    LocalMux I__2661 (
            .O(N__22455),
            .I(N__22445));
    InMux I__2660 (
            .O(N__22454),
            .I(N__22440));
    InMux I__2659 (
            .O(N__22451),
            .I(N__22440));
    Span4Mux_h I__2658 (
            .O(N__22448),
            .I(N__22437));
    Odrv4 I__2657 (
            .O(N__22445),
            .I(\RTD.mode ));
    LocalMux I__2656 (
            .O(N__22440),
            .I(\RTD.mode ));
    Odrv4 I__2655 (
            .O(N__22437),
            .I(\RTD.mode ));
    InMux I__2654 (
            .O(N__22430),
            .I(N__22427));
    LocalMux I__2653 (
            .O(N__22427),
            .I(N__22422));
    InMux I__2652 (
            .O(N__22426),
            .I(N__22417));
    InMux I__2651 (
            .O(N__22425),
            .I(N__22417));
    Span4Mux_v I__2650 (
            .O(N__22422),
            .I(N__22412));
    LocalMux I__2649 (
            .O(N__22417),
            .I(N__22412));
    Span4Mux_h I__2648 (
            .O(N__22412),
            .I(N__22409));
    Span4Mux_h I__2647 (
            .O(N__22409),
            .I(N__22406));
    Sp12to4 I__2646 (
            .O(N__22406),
            .I(N__22403));
    Span12Mux_v I__2645 (
            .O(N__22403),
            .I(N__22400));
    Odrv12 I__2644 (
            .O(N__22400),
            .I(RTD_DRDY));
    InMux I__2643 (
            .O(N__22397),
            .I(N__22394));
    LocalMux I__2642 (
            .O(N__22394),
            .I(N__22391));
    Span4Mux_h I__2641 (
            .O(N__22391),
            .I(N__22384));
    InMux I__2640 (
            .O(N__22390),
            .I(N__22379));
    InMux I__2639 (
            .O(N__22389),
            .I(N__22379));
    InMux I__2638 (
            .O(N__22388),
            .I(N__22376));
    InMux I__2637 (
            .O(N__22387),
            .I(N__22373));
    Odrv4 I__2636 (
            .O(N__22384),
            .I(\RTD.adress_7_N_1340_7 ));
    LocalMux I__2635 (
            .O(N__22379),
            .I(\RTD.adress_7_N_1340_7 ));
    LocalMux I__2634 (
            .O(N__22376),
            .I(\RTD.adress_7_N_1340_7 ));
    LocalMux I__2633 (
            .O(N__22373),
            .I(\RTD.adress_7_N_1340_7 ));
    InMux I__2632 (
            .O(N__22364),
            .I(N__22361));
    LocalMux I__2631 (
            .O(N__22361),
            .I(\RTD.n16669 ));
    CascadeMux I__2630 (
            .O(N__22358),
            .I(\RTD.n16669_cascade_ ));
    IoInMux I__2629 (
            .O(N__22355),
            .I(N__22352));
    LocalMux I__2628 (
            .O(N__22352),
            .I(N__22349));
    IoSpan4Mux I__2627 (
            .O(N__22349),
            .I(N__22346));
    Span4Mux_s0_h I__2626 (
            .O(N__22346),
            .I(N__22343));
    Sp12to4 I__2625 (
            .O(N__22343),
            .I(N__22340));
    Span12Mux_s11_h I__2624 (
            .O(N__22340),
            .I(N__22337));
    Odrv12 I__2623 (
            .O(N__22337),
            .I(RTD_CS));
    CEMux I__2622 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__2621 (
            .O(N__22331),
            .I(N__22328));
    Span4Mux_h I__2620 (
            .O(N__22328),
            .I(N__22325));
    Span4Mux_h I__2619 (
            .O(N__22325),
            .I(N__22322));
    Span4Mux_v I__2618 (
            .O(N__22322),
            .I(N__22319));
    Odrv4 I__2617 (
            .O(N__22319),
            .I(\RTD.n11703 ));
    InMux I__2616 (
            .O(N__22316),
            .I(N__22312));
    InMux I__2615 (
            .O(N__22315),
            .I(N__22309));
    LocalMux I__2614 (
            .O(N__22312),
            .I(\RTD.cfg_buf_1 ));
    LocalMux I__2613 (
            .O(N__22309),
            .I(\RTD.cfg_buf_1 ));
    InMux I__2612 (
            .O(N__22304),
            .I(N__22301));
    LocalMux I__2611 (
            .O(N__22301),
            .I(\RTD.n12_adj_1397 ));
    InMux I__2610 (
            .O(N__22298),
            .I(N__22295));
    LocalMux I__2609 (
            .O(N__22295),
            .I(N__22291));
    CascadeMux I__2608 (
            .O(N__22294),
            .I(N__22288));
    Span4Mux_h I__2607 (
            .O(N__22291),
            .I(N__22285));
    InMux I__2606 (
            .O(N__22288),
            .I(N__22282));
    Odrv4 I__2605 (
            .O(N__22285),
            .I(buf_adcdata_vdc_23));
    LocalMux I__2604 (
            .O(N__22282),
            .I(buf_adcdata_vdc_23));
    InMux I__2603 (
            .O(N__22277),
            .I(N__22274));
    LocalMux I__2602 (
            .O(N__22274),
            .I(N__22271));
    Span4Mux_v I__2601 (
            .O(N__22271),
            .I(N__22268));
    Span4Mux_h I__2600 (
            .O(N__22268),
            .I(N__22265));
    Sp12to4 I__2599 (
            .O(N__22265),
            .I(N__22260));
    InMux I__2598 (
            .O(N__22264),
            .I(N__22257));
    InMux I__2597 (
            .O(N__22263),
            .I(N__22254));
    Span12Mux_h I__2596 (
            .O(N__22260),
            .I(N__22249));
    LocalMux I__2595 (
            .O(N__22257),
            .I(N__22249));
    LocalMux I__2594 (
            .O(N__22254),
            .I(buf_adcdata_vac_23));
    Odrv12 I__2593 (
            .O(N__22249),
            .I(buf_adcdata_vac_23));
    CascadeMux I__2592 (
            .O(N__22244),
            .I(n19_adj_1526_cascade_));
    CascadeMux I__2591 (
            .O(N__22241),
            .I(n22076_cascade_));
    InMux I__2590 (
            .O(N__22238),
            .I(N__22235));
    LocalMux I__2589 (
            .O(N__22235),
            .I(N__22232));
    Span4Mux_v I__2588 (
            .O(N__22232),
            .I(N__22228));
    InMux I__2587 (
            .O(N__22231),
            .I(N__22225));
    Odrv4 I__2586 (
            .O(N__22228),
            .I(buf_readRTD_15));
    LocalMux I__2585 (
            .O(N__22225),
            .I(buf_readRTD_15));
    InMux I__2584 (
            .O(N__22220),
            .I(N__22217));
    LocalMux I__2583 (
            .O(N__22217),
            .I(n20));
    InMux I__2582 (
            .O(N__22214),
            .I(N__22211));
    LocalMux I__2581 (
            .O(N__22211),
            .I(N__22208));
    Odrv4 I__2580 (
            .O(N__22208),
            .I(\RTD.n22370 ));
    IoInMux I__2579 (
            .O(N__22205),
            .I(N__22202));
    LocalMux I__2578 (
            .O(N__22202),
            .I(N__22199));
    IoSpan4Mux I__2577 (
            .O(N__22199),
            .I(N__22196));
    Span4Mux_s3_h I__2576 (
            .O(N__22196),
            .I(N__22193));
    Span4Mux_h I__2575 (
            .O(N__22193),
            .I(N__22190));
    Span4Mux_h I__2574 (
            .O(N__22190),
            .I(N__22187));
    Sp12to4 I__2573 (
            .O(N__22187),
            .I(N__22184));
    Odrv12 I__2572 (
            .O(N__22184),
            .I(RTD_SCLK));
    CEMux I__2571 (
            .O(N__22181),
            .I(N__22178));
    LocalMux I__2570 (
            .O(N__22178),
            .I(N__22175));
    Span4Mux_h I__2569 (
            .O(N__22175),
            .I(N__22172));
    Odrv4 I__2568 (
            .O(N__22172),
            .I(\RTD.n8 ));
    InMux I__2567 (
            .O(N__22169),
            .I(N__22147));
    InMux I__2566 (
            .O(N__22168),
            .I(N__22147));
    InMux I__2565 (
            .O(N__22167),
            .I(N__22147));
    InMux I__2564 (
            .O(N__22166),
            .I(N__22140));
    InMux I__2563 (
            .O(N__22165),
            .I(N__22140));
    InMux I__2562 (
            .O(N__22164),
            .I(N__22140));
    InMux I__2561 (
            .O(N__22163),
            .I(N__22133));
    InMux I__2560 (
            .O(N__22162),
            .I(N__22133));
    InMux I__2559 (
            .O(N__22161),
            .I(N__22133));
    InMux I__2558 (
            .O(N__22160),
            .I(N__22118));
    InMux I__2557 (
            .O(N__22159),
            .I(N__22118));
    InMux I__2556 (
            .O(N__22158),
            .I(N__22118));
    InMux I__2555 (
            .O(N__22157),
            .I(N__22118));
    InMux I__2554 (
            .O(N__22156),
            .I(N__22118));
    InMux I__2553 (
            .O(N__22155),
            .I(N__22118));
    InMux I__2552 (
            .O(N__22154),
            .I(N__22118));
    LocalMux I__2551 (
            .O(N__22147),
            .I(N__22115));
    LocalMux I__2550 (
            .O(N__22140),
            .I(N__22112));
    LocalMux I__2549 (
            .O(N__22133),
            .I(N__22109));
    LocalMux I__2548 (
            .O(N__22118),
            .I(N__22106));
    Span4Mux_v I__2547 (
            .O(N__22115),
            .I(N__22103));
    Span4Mux_v I__2546 (
            .O(N__22112),
            .I(N__22098));
    Span4Mux_h I__2545 (
            .O(N__22109),
            .I(N__22098));
    Span4Mux_h I__2544 (
            .O(N__22106),
            .I(N__22095));
    Odrv4 I__2543 (
            .O(N__22103),
            .I(n13309));
    Odrv4 I__2542 (
            .O(N__22098),
            .I(n13309));
    Odrv4 I__2541 (
            .O(N__22095),
            .I(n13309));
    CascadeMux I__2540 (
            .O(N__22088),
            .I(N__22083));
    InMux I__2539 (
            .O(N__22087),
            .I(N__22076));
    InMux I__2538 (
            .O(N__22086),
            .I(N__22076));
    InMux I__2537 (
            .O(N__22083),
            .I(N__22076));
    LocalMux I__2536 (
            .O(N__22076),
            .I(cmd_rdadctmp_30));
    CascadeMux I__2535 (
            .O(N__22073),
            .I(N__22069));
    CascadeMux I__2534 (
            .O(N__22072),
            .I(N__22066));
    InMux I__2533 (
            .O(N__22069),
            .I(N__22061));
    InMux I__2532 (
            .O(N__22066),
            .I(N__22061));
    LocalMux I__2531 (
            .O(N__22061),
            .I(cmd_rdadctmp_31));
    InMux I__2530 (
            .O(N__22058),
            .I(N__22055));
    LocalMux I__2529 (
            .O(N__22055),
            .I(N__22051));
    InMux I__2528 (
            .O(N__22054),
            .I(N__22048));
    Odrv4 I__2527 (
            .O(N__22051),
            .I(buf_adcdata_vdc_5));
    LocalMux I__2526 (
            .O(N__22048),
            .I(buf_adcdata_vdc_5));
    InMux I__2525 (
            .O(N__22043),
            .I(N__22040));
    LocalMux I__2524 (
            .O(N__22040),
            .I(N__22036));
    InMux I__2523 (
            .O(N__22039),
            .I(N__22033));
    Odrv12 I__2522 (
            .O(N__22036),
            .I(buf_adcdata_vdc_4));
    LocalMux I__2521 (
            .O(N__22033),
            .I(buf_adcdata_vdc_4));
    CascadeMux I__2520 (
            .O(N__22028),
            .I(N__22025));
    InMux I__2519 (
            .O(N__22025),
            .I(N__22022));
    LocalMux I__2518 (
            .O(N__22022),
            .I(N__22018));
    InMux I__2517 (
            .O(N__22021),
            .I(N__22015));
    Odrv4 I__2516 (
            .O(N__22018),
            .I(buf_adcdata_vdc_20));
    LocalMux I__2515 (
            .O(N__22015),
            .I(buf_adcdata_vdc_20));
    CEMux I__2514 (
            .O(N__22010),
            .I(N__22007));
    LocalMux I__2513 (
            .O(N__22007),
            .I(N__22004));
    Span4Mux_h I__2512 (
            .O(N__22004),
            .I(N__22001));
    Odrv4 I__2511 (
            .O(N__22001),
            .I(\ADC_VDC.n47 ));
    CascadeMux I__2510 (
            .O(N__21998),
            .I(N__21995));
    InMux I__2509 (
            .O(N__21995),
            .I(N__21986));
    InMux I__2508 (
            .O(N__21994),
            .I(N__21986));
    InMux I__2507 (
            .O(N__21993),
            .I(N__21986));
    LocalMux I__2506 (
            .O(N__21986),
            .I(cmd_rdadctmp_15));
    InMux I__2505 (
            .O(N__21983),
            .I(N__21980));
    LocalMux I__2504 (
            .O(N__21980),
            .I(n19_adj_1631));
    InMux I__2503 (
            .O(N__21977),
            .I(N__21974));
    LocalMux I__2502 (
            .O(N__21974),
            .I(N__21970));
    InMux I__2501 (
            .O(N__21973),
            .I(N__21966));
    Span12Mux_s10_v I__2500 (
            .O(N__21970),
            .I(N__21963));
    InMux I__2499 (
            .O(N__21969),
            .I(N__21960));
    LocalMux I__2498 (
            .O(N__21966),
            .I(buf_adcdata_vac_5));
    Odrv12 I__2497 (
            .O(N__21963),
            .I(buf_adcdata_vac_5));
    LocalMux I__2496 (
            .O(N__21960),
            .I(buf_adcdata_vac_5));
    InMux I__2495 (
            .O(N__21953),
            .I(N__21950));
    LocalMux I__2494 (
            .O(N__21950),
            .I(N__21947));
    Span4Mux_v I__2493 (
            .O(N__21947),
            .I(N__21944));
    Sp12to4 I__2492 (
            .O(N__21944),
            .I(N__21939));
    InMux I__2491 (
            .O(N__21943),
            .I(N__21936));
    InMux I__2490 (
            .O(N__21942),
            .I(N__21933));
    Span12Mux_h I__2489 (
            .O(N__21939),
            .I(N__21928));
    LocalMux I__2488 (
            .O(N__21936),
            .I(N__21928));
    LocalMux I__2487 (
            .O(N__21933),
            .I(buf_adcdata_vac_20));
    Odrv12 I__2486 (
            .O(N__21928),
            .I(buf_adcdata_vac_20));
    CascadeMux I__2485 (
            .O(N__21923),
            .I(N__21919));
    InMux I__2484 (
            .O(N__21922),
            .I(N__21916));
    InMux I__2483 (
            .O(N__21919),
            .I(N__21913));
    LocalMux I__2482 (
            .O(N__21916),
            .I(N__21910));
    LocalMux I__2481 (
            .O(N__21913),
            .I(N__21906));
    Span4Mux_h I__2480 (
            .O(N__21910),
            .I(N__21903));
    InMux I__2479 (
            .O(N__21909),
            .I(N__21900));
    Odrv12 I__2478 (
            .O(N__21906),
            .I(cmd_rdadctmp_29));
    Odrv4 I__2477 (
            .O(N__21903),
            .I(cmd_rdadctmp_29));
    LocalMux I__2476 (
            .O(N__21900),
            .I(cmd_rdadctmp_29));
    InMux I__2475 (
            .O(N__21893),
            .I(N__21890));
    LocalMux I__2474 (
            .O(N__21890),
            .I(N__21887));
    Span4Mux_h I__2473 (
            .O(N__21887),
            .I(N__21882));
    InMux I__2472 (
            .O(N__21886),
            .I(N__21877));
    InMux I__2471 (
            .O(N__21885),
            .I(N__21877));
    Odrv4 I__2470 (
            .O(N__21882),
            .I(buf_adcdata_vac_4));
    LocalMux I__2469 (
            .O(N__21877),
            .I(buf_adcdata_vac_4));
    CascadeMux I__2468 (
            .O(N__21872),
            .I(n19_adj_1636_cascade_));
    InMux I__2467 (
            .O(N__21869),
            .I(N__21866));
    LocalMux I__2466 (
            .O(N__21866),
            .I(N__21863));
    Span4Mux_h I__2465 (
            .O(N__21863),
            .I(N__21858));
    InMux I__2464 (
            .O(N__21862),
            .I(N__21853));
    InMux I__2463 (
            .O(N__21861),
            .I(N__21853));
    Odrv4 I__2462 (
            .O(N__21858),
            .I(buf_adcdata_iac_4));
    LocalMux I__2461 (
            .O(N__21853),
            .I(buf_adcdata_iac_4));
    InMux I__2460 (
            .O(N__21848),
            .I(N__21845));
    LocalMux I__2459 (
            .O(N__21845),
            .I(N__21842));
    Span4Mux_h I__2458 (
            .O(N__21842),
            .I(N__21839));
    Odrv4 I__2457 (
            .O(N__21839),
            .I(buf_data_iac_4));
    CascadeMux I__2456 (
            .O(N__21836),
            .I(n22_adj_1637_cascade_));
    InMux I__2455 (
            .O(N__21833),
            .I(N__21830));
    LocalMux I__2454 (
            .O(N__21830),
            .I(N__21827));
    Span12Mux_v I__2453 (
            .O(N__21827),
            .I(N__21823));
    InMux I__2452 (
            .O(N__21826),
            .I(N__21820));
    Odrv12 I__2451 (
            .O(N__21823),
            .I(cmd_rdadctmp_4));
    LocalMux I__2450 (
            .O(N__21820),
            .I(cmd_rdadctmp_4));
    CascadeMux I__2449 (
            .O(N__21815),
            .I(N__21811));
    InMux I__2448 (
            .O(N__21814),
            .I(N__21806));
    InMux I__2447 (
            .O(N__21811),
            .I(N__21806));
    LocalMux I__2446 (
            .O(N__21806),
            .I(cmd_rdadctmp_5));
    CascadeMux I__2445 (
            .O(N__21803),
            .I(N__21800));
    InMux I__2444 (
            .O(N__21800),
            .I(N__21797));
    LocalMux I__2443 (
            .O(N__21797),
            .I(\CLK_DDS.tmp_buf_2 ));
    CascadeMux I__2442 (
            .O(N__21794),
            .I(N__21791));
    InMux I__2441 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__2440 (
            .O(N__21788),
            .I(\CLK_DDS.tmp_buf_3 ));
    CascadeMux I__2439 (
            .O(N__21785),
            .I(N__21782));
    InMux I__2438 (
            .O(N__21782),
            .I(N__21779));
    LocalMux I__2437 (
            .O(N__21779),
            .I(\CLK_DDS.tmp_buf_4 ));
    InMux I__2436 (
            .O(N__21776),
            .I(N__21773));
    LocalMux I__2435 (
            .O(N__21773),
            .I(\CLK_DDS.tmp_buf_5 ));
    CascadeMux I__2434 (
            .O(N__21770),
            .I(N__21767));
    InMux I__2433 (
            .O(N__21767),
            .I(N__21764));
    LocalMux I__2432 (
            .O(N__21764),
            .I(\CLK_DDS.tmp_buf_6 ));
    InMux I__2431 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__2430 (
            .O(N__21758),
            .I(\CLK_DDS.tmp_buf_7 ));
    CEMux I__2429 (
            .O(N__21755),
            .I(N__21752));
    LocalMux I__2428 (
            .O(N__21752),
            .I(N__21749));
    Span4Mux_h I__2427 (
            .O(N__21749),
            .I(N__21746));
    Span4Mux_v I__2426 (
            .O(N__21746),
            .I(N__21743));
    Odrv4 I__2425 (
            .O(N__21743),
            .I(\CLK_DDS.n9_adj_1395 ));
    CascadeMux I__2424 (
            .O(N__21740),
            .I(N__21737));
    InMux I__2423 (
            .O(N__21737),
            .I(N__21730));
    InMux I__2422 (
            .O(N__21736),
            .I(N__21730));
    InMux I__2421 (
            .O(N__21735),
            .I(N__21727));
    LocalMux I__2420 (
            .O(N__21730),
            .I(cmd_rdadctmp_30_adj_1420));
    LocalMux I__2419 (
            .O(N__21727),
            .I(cmd_rdadctmp_30_adj_1420));
    IoInMux I__2418 (
            .O(N__21722),
            .I(N__21719));
    LocalMux I__2417 (
            .O(N__21719),
            .I(N__21716));
    Span12Mux_s9_v I__2416 (
            .O(N__21716),
            .I(N__21712));
    InMux I__2415 (
            .O(N__21715),
            .I(N__21709));
    Odrv12 I__2414 (
            .O(N__21712),
            .I(DDS_MOSI1));
    LocalMux I__2413 (
            .O(N__21709),
            .I(DDS_MOSI1));
    CascadeMux I__2412 (
            .O(N__21704),
            .I(N__21701));
    InMux I__2411 (
            .O(N__21701),
            .I(N__21696));
    InMux I__2410 (
            .O(N__21700),
            .I(N__21691));
    InMux I__2409 (
            .O(N__21699),
            .I(N__21691));
    LocalMux I__2408 (
            .O(N__21696),
            .I(cmd_rdadctmp_23_adj_1427));
    LocalMux I__2407 (
            .O(N__21691),
            .I(cmd_rdadctmp_23_adj_1427));
    CascadeMux I__2406 (
            .O(N__21686),
            .I(N__21682));
    CascadeMux I__2405 (
            .O(N__21685),
            .I(N__21678));
    InMux I__2404 (
            .O(N__21682),
            .I(N__21671));
    InMux I__2403 (
            .O(N__21681),
            .I(N__21671));
    InMux I__2402 (
            .O(N__21678),
            .I(N__21671));
    LocalMux I__2401 (
            .O(N__21671),
            .I(cmd_rdadctmp_24_adj_1426));
    CascadeMux I__2400 (
            .O(N__21668),
            .I(N__21663));
    CascadeMux I__2399 (
            .O(N__21667),
            .I(N__21660));
    InMux I__2398 (
            .O(N__21666),
            .I(N__21655));
    InMux I__2397 (
            .O(N__21663),
            .I(N__21655));
    InMux I__2396 (
            .O(N__21660),
            .I(N__21652));
    LocalMux I__2395 (
            .O(N__21655),
            .I(cmd_rdadctmp_26_adj_1424));
    LocalMux I__2394 (
            .O(N__21652),
            .I(cmd_rdadctmp_26_adj_1424));
    CascadeMux I__2393 (
            .O(N__21647),
            .I(N__21644));
    InMux I__2392 (
            .O(N__21644),
            .I(N__21641));
    LocalMux I__2391 (
            .O(N__21641),
            .I(N__21638));
    Span4Mux_v I__2390 (
            .O(N__21638),
            .I(N__21635));
    Span4Mux_v I__2389 (
            .O(N__21635),
            .I(N__21632));
    Odrv4 I__2388 (
            .O(N__21632),
            .I(\CLK_DDS.tmp_buf_1 ));
    CascadeMux I__2387 (
            .O(N__21629),
            .I(N__21625));
    CascadeMux I__2386 (
            .O(N__21628),
            .I(N__21622));
    InMux I__2385 (
            .O(N__21625),
            .I(N__21618));
    InMux I__2384 (
            .O(N__21622),
            .I(N__21613));
    InMux I__2383 (
            .O(N__21621),
            .I(N__21613));
    LocalMux I__2382 (
            .O(N__21618),
            .I(read_buf_7));
    LocalMux I__2381 (
            .O(N__21613),
            .I(read_buf_7));
    CascadeMux I__2380 (
            .O(N__21608),
            .I(N__21603));
    CascadeMux I__2379 (
            .O(N__21607),
            .I(N__21600));
    InMux I__2378 (
            .O(N__21606),
            .I(N__21595));
    InMux I__2377 (
            .O(N__21603),
            .I(N__21595));
    InMux I__2376 (
            .O(N__21600),
            .I(N__21592));
    LocalMux I__2375 (
            .O(N__21595),
            .I(read_buf_2));
    LocalMux I__2374 (
            .O(N__21592),
            .I(read_buf_2));
    CascadeMux I__2373 (
            .O(N__21587),
            .I(N__21582));
    CascadeMux I__2372 (
            .O(N__21586),
            .I(N__21579));
    CascadeMux I__2371 (
            .O(N__21585),
            .I(N__21576));
    InMux I__2370 (
            .O(N__21582),
            .I(N__21573));
    InMux I__2369 (
            .O(N__21579),
            .I(N__21568));
    InMux I__2368 (
            .O(N__21576),
            .I(N__21568));
    LocalMux I__2367 (
            .O(N__21573),
            .I(read_buf_3));
    LocalMux I__2366 (
            .O(N__21568),
            .I(read_buf_3));
    CascadeMux I__2365 (
            .O(N__21563),
            .I(N__21556));
    CascadeMux I__2364 (
            .O(N__21562),
            .I(N__21553));
    CascadeMux I__2363 (
            .O(N__21561),
            .I(N__21550));
    CascadeMux I__2362 (
            .O(N__21560),
            .I(N__21547));
    CascadeMux I__2361 (
            .O(N__21559),
            .I(N__21542));
    InMux I__2360 (
            .O(N__21556),
            .I(N__21529));
    InMux I__2359 (
            .O(N__21553),
            .I(N__21529));
    InMux I__2358 (
            .O(N__21550),
            .I(N__21529));
    InMux I__2357 (
            .O(N__21547),
            .I(N__21529));
    InMux I__2356 (
            .O(N__21546),
            .I(N__21529));
    InMux I__2355 (
            .O(N__21545),
            .I(N__21529));
    InMux I__2354 (
            .O(N__21542),
            .I(N__21526));
    LocalMux I__2353 (
            .O(N__21529),
            .I(N__21513));
    LocalMux I__2352 (
            .O(N__21526),
            .I(N__21513));
    InMux I__2351 (
            .O(N__21525),
            .I(N__21510));
    InMux I__2350 (
            .O(N__21524),
            .I(N__21505));
    InMux I__2349 (
            .O(N__21523),
            .I(N__21505));
    InMux I__2348 (
            .O(N__21522),
            .I(N__21498));
    InMux I__2347 (
            .O(N__21521),
            .I(N__21498));
    InMux I__2346 (
            .O(N__21520),
            .I(N__21498));
    InMux I__2345 (
            .O(N__21519),
            .I(N__21493));
    InMux I__2344 (
            .O(N__21518),
            .I(N__21493));
    Span4Mux_h I__2343 (
            .O(N__21513),
            .I(N__21490));
    LocalMux I__2342 (
            .O(N__21510),
            .I(n1_adj_1601));
    LocalMux I__2341 (
            .O(N__21505),
            .I(n1_adj_1601));
    LocalMux I__2340 (
            .O(N__21498),
            .I(n1_adj_1601));
    LocalMux I__2339 (
            .O(N__21493),
            .I(n1_adj_1601));
    Odrv4 I__2338 (
            .O(N__21490),
            .I(n1_adj_1601));
    InMux I__2337 (
            .O(N__21479),
            .I(N__21470));
    InMux I__2336 (
            .O(N__21478),
            .I(N__21470));
    InMux I__2335 (
            .O(N__21477),
            .I(N__21470));
    LocalMux I__2334 (
            .O(N__21470),
            .I(read_buf_4));
    CascadeMux I__2333 (
            .O(N__21467),
            .I(n1_adj_1601_cascade_));
    InMux I__2332 (
            .O(N__21464),
            .I(N__21459));
    InMux I__2331 (
            .O(N__21463),
            .I(N__21454));
    InMux I__2330 (
            .O(N__21462),
            .I(N__21454));
    LocalMux I__2329 (
            .O(N__21459),
            .I(read_buf_5));
    LocalMux I__2328 (
            .O(N__21454),
            .I(read_buf_5));
    CascadeMux I__2327 (
            .O(N__21449),
            .I(N__21445));
    CascadeMux I__2326 (
            .O(N__21448),
            .I(N__21441));
    InMux I__2325 (
            .O(N__21445),
            .I(N__21438));
    InMux I__2324 (
            .O(N__21444),
            .I(N__21433));
    InMux I__2323 (
            .O(N__21441),
            .I(N__21433));
    LocalMux I__2322 (
            .O(N__21438),
            .I(cmd_rdadctmp_29_adj_1421));
    LocalMux I__2321 (
            .O(N__21433),
            .I(cmd_rdadctmp_29_adj_1421));
    InMux I__2320 (
            .O(N__21428),
            .I(N__21425));
    LocalMux I__2319 (
            .O(N__21425),
            .I(\RTD.cfg_tmp_2 ));
    InMux I__2318 (
            .O(N__21422),
            .I(N__21419));
    LocalMux I__2317 (
            .O(N__21419),
            .I(\RTD.cfg_tmp_3 ));
    InMux I__2316 (
            .O(N__21416),
            .I(N__21413));
    LocalMux I__2315 (
            .O(N__21413),
            .I(\RTD.cfg_tmp_4 ));
    InMux I__2314 (
            .O(N__21410),
            .I(N__21407));
    LocalMux I__2313 (
            .O(N__21407),
            .I(\RTD.cfg_tmp_5 ));
    InMux I__2312 (
            .O(N__21404),
            .I(N__21401));
    LocalMux I__2311 (
            .O(N__21401),
            .I(\RTD.cfg_tmp_6 ));
    CascadeMux I__2310 (
            .O(N__21398),
            .I(N__21395));
    InMux I__2309 (
            .O(N__21395),
            .I(N__21391));
    InMux I__2308 (
            .O(N__21394),
            .I(N__21388));
    LocalMux I__2307 (
            .O(N__21391),
            .I(\RTD.cfg_tmp_7 ));
    LocalMux I__2306 (
            .O(N__21388),
            .I(\RTD.cfg_tmp_7 ));
    InMux I__2305 (
            .O(N__21383),
            .I(N__21380));
    LocalMux I__2304 (
            .O(N__21380),
            .I(\RTD.cfg_tmp_0 ));
    CEMux I__2303 (
            .O(N__21377),
            .I(N__21373));
    InMux I__2302 (
            .O(N__21376),
            .I(N__21370));
    LocalMux I__2301 (
            .O(N__21373),
            .I(\RTD.n13228 ));
    LocalMux I__2300 (
            .O(N__21370),
            .I(\RTD.n13228 ));
    SRMux I__2299 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__2298 (
            .O(N__21362),
            .I(N__21359));
    Span4Mux_v I__2297 (
            .O(N__21359),
            .I(N__21356));
    Odrv4 I__2296 (
            .O(N__21356),
            .I(\RTD.n15015 ));
    CascadeMux I__2295 (
            .O(N__21353),
            .I(\RTD.n7333_cascade_ ));
    CascadeMux I__2294 (
            .O(N__21350),
            .I(\RTD.n13_cascade_ ));
    CEMux I__2293 (
            .O(N__21347),
            .I(N__21344));
    LocalMux I__2292 (
            .O(N__21344),
            .I(N__21341));
    Odrv4 I__2291 (
            .O(N__21341),
            .I(\RTD.n11734 ));
    InMux I__2290 (
            .O(N__21338),
            .I(N__21335));
    LocalMux I__2289 (
            .O(N__21335),
            .I(N__21330));
    InMux I__2288 (
            .O(N__21334),
            .I(N__21327));
    InMux I__2287 (
            .O(N__21333),
            .I(N__21324));
    Odrv4 I__2286 (
            .O(N__21330),
            .I(\RTD.n7333 ));
    LocalMux I__2285 (
            .O(N__21327),
            .I(\RTD.n7333 ));
    LocalMux I__2284 (
            .O(N__21324),
            .I(\RTD.n7333 ));
    InMux I__2283 (
            .O(N__21317),
            .I(N__21314));
    LocalMux I__2282 (
            .O(N__21314),
            .I(\RTD.cfg_tmp_1 ));
    InMux I__2281 (
            .O(N__21311),
            .I(N__21308));
    LocalMux I__2280 (
            .O(N__21308),
            .I(N__21305));
    Span4Mux_h I__2279 (
            .O(N__21305),
            .I(N__21301));
    CascadeMux I__2278 (
            .O(N__21304),
            .I(N__21298));
    Span4Mux_h I__2277 (
            .O(N__21301),
            .I(N__21295));
    InMux I__2276 (
            .O(N__21298),
            .I(N__21292));
    Odrv4 I__2275 (
            .O(N__21295),
            .I(read_buf_15));
    LocalMux I__2274 (
            .O(N__21292),
            .I(read_buf_15));
    CascadeMux I__2273 (
            .O(N__21287),
            .I(n11730_cascade_));
    InMux I__2272 (
            .O(N__21284),
            .I(N__21280));
    InMux I__2271 (
            .O(N__21283),
            .I(N__21277));
    LocalMux I__2270 (
            .O(N__21280),
            .I(adress_6));
    LocalMux I__2269 (
            .O(N__21277),
            .I(adress_6));
    InMux I__2268 (
            .O(N__21272),
            .I(N__21268));
    InMux I__2267 (
            .O(N__21271),
            .I(N__21265));
    LocalMux I__2266 (
            .O(N__21268),
            .I(\RTD.cfg_buf_6 ));
    LocalMux I__2265 (
            .O(N__21265),
            .I(\RTD.cfg_buf_6 ));
    InMux I__2264 (
            .O(N__21260),
            .I(N__21256));
    InMux I__2263 (
            .O(N__21259),
            .I(N__21253));
    LocalMux I__2262 (
            .O(N__21256),
            .I(\RTD.cfg_buf_0 ));
    LocalMux I__2261 (
            .O(N__21253),
            .I(\RTD.cfg_buf_0 ));
    CascadeMux I__2260 (
            .O(N__21248),
            .I(\RTD.n9_cascade_ ));
    CascadeMux I__2259 (
            .O(N__21245),
            .I(\RTD.adress_7_N_1340_7_cascade_ ));
    CascadeMux I__2258 (
            .O(N__21242),
            .I(N__21239));
    InMux I__2257 (
            .O(N__21239),
            .I(N__21235));
    InMux I__2256 (
            .O(N__21238),
            .I(N__21232));
    LocalMux I__2255 (
            .O(N__21235),
            .I(\RTD.adress_7 ));
    LocalMux I__2254 (
            .O(N__21232),
            .I(\RTD.adress_7 ));
    CascadeMux I__2253 (
            .O(N__21227),
            .I(N__21224));
    InMux I__2252 (
            .O(N__21224),
            .I(N__21221));
    LocalMux I__2251 (
            .O(N__21221),
            .I(N__21218));
    Odrv4 I__2250 (
            .O(N__21218),
            .I(adress_0));
    CEMux I__2249 (
            .O(N__21215),
            .I(N__21212));
    LocalMux I__2248 (
            .O(N__21212),
            .I(N__21203));
    InMux I__2247 (
            .O(N__21211),
            .I(N__21192));
    InMux I__2246 (
            .O(N__21210),
            .I(N__21192));
    InMux I__2245 (
            .O(N__21209),
            .I(N__21192));
    InMux I__2244 (
            .O(N__21208),
            .I(N__21192));
    InMux I__2243 (
            .O(N__21207),
            .I(N__21192));
    InMux I__2242 (
            .O(N__21206),
            .I(N__21189));
    Odrv4 I__2241 (
            .O(N__21203),
            .I(n13181));
    LocalMux I__2240 (
            .O(N__21192),
            .I(n13181));
    LocalMux I__2239 (
            .O(N__21189),
            .I(n13181));
    InMux I__2238 (
            .O(N__21182),
            .I(N__21178));
    InMux I__2237 (
            .O(N__21181),
            .I(N__21175));
    LocalMux I__2236 (
            .O(N__21178),
            .I(\RTD.cfg_buf_5 ));
    LocalMux I__2235 (
            .O(N__21175),
            .I(\RTD.cfg_buf_5 ));
    CascadeMux I__2234 (
            .O(N__21170),
            .I(N__21167));
    InMux I__2233 (
            .O(N__21167),
            .I(N__21163));
    InMux I__2232 (
            .O(N__21166),
            .I(N__21160));
    LocalMux I__2231 (
            .O(N__21163),
            .I(\RTD.cfg_buf_3 ));
    LocalMux I__2230 (
            .O(N__21160),
            .I(\RTD.cfg_buf_3 ));
    InMux I__2229 (
            .O(N__21155),
            .I(N__21152));
    LocalMux I__2228 (
            .O(N__21152),
            .I(\RTD.n11 ));
    CascadeMux I__2227 (
            .O(N__21149),
            .I(\ADC_VDC.n13038_cascade_ ));
    InMux I__2226 (
            .O(N__21146),
            .I(N__21143));
    LocalMux I__2225 (
            .O(N__21143),
            .I(N__21140));
    Odrv4 I__2224 (
            .O(N__21140),
            .I(\ADC_VDC.n20659 ));
    CascadeMux I__2223 (
            .O(N__21137),
            .I(\ADC_VDC.n17432_cascade_ ));
    SRMux I__2222 (
            .O(N__21134),
            .I(N__21131));
    LocalMux I__2221 (
            .O(N__21131),
            .I(N__21128));
    Span4Mux_h I__2220 (
            .O(N__21128),
            .I(N__21125));
    Odrv4 I__2219 (
            .O(N__21125),
            .I(\ADC_VDC.n18466 ));
    CascadeMux I__2218 (
            .O(N__21122),
            .I(N__21119));
    InMux I__2217 (
            .O(N__21119),
            .I(N__21116));
    LocalMux I__2216 (
            .O(N__21116),
            .I(N__21112));
    CascadeMux I__2215 (
            .O(N__21115),
            .I(N__21108));
    Span4Mux_h I__2214 (
            .O(N__21112),
            .I(N__21105));
    InMux I__2213 (
            .O(N__21111),
            .I(N__21100));
    InMux I__2212 (
            .O(N__21108),
            .I(N__21100));
    Odrv4 I__2211 (
            .O(N__21105),
            .I(read_buf_11));
    LocalMux I__2210 (
            .O(N__21100),
            .I(read_buf_11));
    CascadeMux I__2209 (
            .O(N__21095),
            .I(\ADC_VDC.n11692_cascade_ ));
    IoInMux I__2208 (
            .O(N__21092),
            .I(N__21089));
    LocalMux I__2207 (
            .O(N__21089),
            .I(N__21085));
    InMux I__2206 (
            .O(N__21088),
            .I(N__21082));
    Span12Mux_s5_h I__2205 (
            .O(N__21085),
            .I(N__21079));
    LocalMux I__2204 (
            .O(N__21082),
            .I(N__21076));
    Odrv12 I__2203 (
            .O(N__21079),
            .I(VDC_SCLK));
    Odrv4 I__2202 (
            .O(N__21076),
            .I(VDC_SCLK));
    CascadeMux I__2201 (
            .O(N__21071),
            .I(N__21064));
    InMux I__2200 (
            .O(N__21070),
            .I(N__21061));
    InMux I__2199 (
            .O(N__21069),
            .I(N__21058));
    InMux I__2198 (
            .O(N__21068),
            .I(N__21053));
    InMux I__2197 (
            .O(N__21067),
            .I(N__21053));
    InMux I__2196 (
            .O(N__21064),
            .I(N__21050));
    LocalMux I__2195 (
            .O(N__21061),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__2194 (
            .O(N__21058),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__2193 (
            .O(N__21053),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__2192 (
            .O(N__21050),
            .I(\ADC_VDC.bit_cnt_1 ));
    InMux I__2191 (
            .O(N__21041),
            .I(N__21037));
    InMux I__2190 (
            .O(N__21040),
            .I(N__21034));
    LocalMux I__2189 (
            .O(N__21037),
            .I(\ADC_VDC.n20534 ));
    LocalMux I__2188 (
            .O(N__21034),
            .I(\ADC_VDC.n20534 ));
    CascadeMux I__2187 (
            .O(N__21029),
            .I(N__21024));
    CascadeMux I__2186 (
            .O(N__21028),
            .I(N__21021));
    CascadeMux I__2185 (
            .O(N__21027),
            .I(N__21017));
    InMux I__2184 (
            .O(N__21024),
            .I(N__21011));
    InMux I__2183 (
            .O(N__21021),
            .I(N__21011));
    InMux I__2182 (
            .O(N__21020),
            .I(N__21008));
    InMux I__2181 (
            .O(N__21017),
            .I(N__21005));
    InMux I__2180 (
            .O(N__21016),
            .I(N__21002));
    LocalMux I__2179 (
            .O(N__21011),
            .I(N__20999));
    LocalMux I__2178 (
            .O(N__21008),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__2177 (
            .O(N__21005),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__2176 (
            .O(N__21002),
            .I(\ADC_VDC.bit_cnt_4 ));
    Odrv4 I__2175 (
            .O(N__20999),
            .I(\ADC_VDC.bit_cnt_4 ));
    InMux I__2174 (
            .O(N__20990),
            .I(N__20987));
    LocalMux I__2173 (
            .O(N__20987),
            .I(N__20984));
    Span4Mux_h I__2172 (
            .O(N__20984),
            .I(N__20981));
    Odrv4 I__2171 (
            .O(N__20981),
            .I(\ADC_VDC.n6_adj_1410 ));
    CascadeMux I__2170 (
            .O(N__20978),
            .I(\ADC_VDC.n11281_cascade_ ));
    InMux I__2169 (
            .O(N__20975),
            .I(N__20968));
    InMux I__2168 (
            .O(N__20974),
            .I(N__20965));
    InMux I__2167 (
            .O(N__20973),
            .I(N__20960));
    InMux I__2166 (
            .O(N__20972),
            .I(N__20960));
    InMux I__2165 (
            .O(N__20971),
            .I(N__20957));
    LocalMux I__2164 (
            .O(N__20968),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__2163 (
            .O(N__20965),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__2162 (
            .O(N__20960),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__2161 (
            .O(N__20957),
            .I(\ADC_VDC.bit_cnt_0 ));
    InMux I__2160 (
            .O(N__20948),
            .I(N__20942));
    InMux I__2159 (
            .O(N__20947),
            .I(N__20942));
    LocalMux I__2158 (
            .O(N__20942),
            .I(\ADC_VDC.n15 ));
    CascadeMux I__2157 (
            .O(N__20939),
            .I(\ADC_VDC.n15_cascade_ ));
    CascadeMux I__2156 (
            .O(N__20936),
            .I(\ADC_VDC.n20746_cascade_ ));
    InMux I__2155 (
            .O(N__20933),
            .I(N__20930));
    LocalMux I__2154 (
            .O(N__20930),
            .I(\ADC_VDC.n72 ));
    CEMux I__2153 (
            .O(N__20927),
            .I(N__20924));
    LocalMux I__2152 (
            .O(N__20924),
            .I(N__20921));
    Odrv4 I__2151 (
            .O(N__20921),
            .I(\ADC_VDC.n12823 ));
    CascadeMux I__2150 (
            .O(N__20918),
            .I(\ADC_VDC.n19_adj_1413_cascade_ ));
    CEMux I__2149 (
            .O(N__20915),
            .I(N__20912));
    LocalMux I__2148 (
            .O(N__20912),
            .I(\ADC_VDC.n17 ));
    SRMux I__2147 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__2146 (
            .O(N__20906),
            .I(N__20903));
    Span4Mux_h I__2145 (
            .O(N__20903),
            .I(N__20900));
    Odrv4 I__2144 (
            .O(N__20900),
            .I(\ADC_VDC.n4 ));
    CascadeMux I__2143 (
            .O(N__20897),
            .I(\ADC_VDC.n10132_cascade_ ));
    InMux I__2142 (
            .O(N__20894),
            .I(N__20888));
    InMux I__2141 (
            .O(N__20893),
            .I(N__20888));
    LocalMux I__2140 (
            .O(N__20888),
            .I(\ADC_VDC.n7_adj_1411 ));
    InMux I__2139 (
            .O(N__20885),
            .I(N__20879));
    InMux I__2138 (
            .O(N__20884),
            .I(N__20879));
    LocalMux I__2137 (
            .O(N__20879),
            .I(\ADC_VDC.n20750 ));
    InMux I__2136 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2135 (
            .O(N__20873),
            .I(\ADC_VDC.n12 ));
    CascadeMux I__2134 (
            .O(N__20870),
            .I(\ADC_VDC.n20750_cascade_ ));
    InMux I__2133 (
            .O(N__20867),
            .I(N__20863));
    InMux I__2132 (
            .O(N__20866),
            .I(N__20860));
    LocalMux I__2131 (
            .O(N__20863),
            .I(\ADC_IAC.bit_cnt_4 ));
    LocalMux I__2130 (
            .O(N__20860),
            .I(\ADC_IAC.bit_cnt_4 ));
    InMux I__2129 (
            .O(N__20855),
            .I(\ADC_IAC.n19418 ));
    InMux I__2128 (
            .O(N__20852),
            .I(N__20848));
    InMux I__2127 (
            .O(N__20851),
            .I(N__20845));
    LocalMux I__2126 (
            .O(N__20848),
            .I(\ADC_IAC.bit_cnt_5 ));
    LocalMux I__2125 (
            .O(N__20845),
            .I(\ADC_IAC.bit_cnt_5 ));
    InMux I__2124 (
            .O(N__20840),
            .I(\ADC_IAC.n19419 ));
    InMux I__2123 (
            .O(N__20837),
            .I(N__20833));
    InMux I__2122 (
            .O(N__20836),
            .I(N__20830));
    LocalMux I__2121 (
            .O(N__20833),
            .I(\ADC_IAC.bit_cnt_6 ));
    LocalMux I__2120 (
            .O(N__20830),
            .I(\ADC_IAC.bit_cnt_6 ));
    InMux I__2119 (
            .O(N__20825),
            .I(\ADC_IAC.n19420 ));
    InMux I__2118 (
            .O(N__20822),
            .I(\ADC_IAC.n19421 ));
    InMux I__2117 (
            .O(N__20819),
            .I(N__20815));
    InMux I__2116 (
            .O(N__20818),
            .I(N__20812));
    LocalMux I__2115 (
            .O(N__20815),
            .I(\ADC_IAC.bit_cnt_7 ));
    LocalMux I__2114 (
            .O(N__20812),
            .I(\ADC_IAC.bit_cnt_7 ));
    CEMux I__2113 (
            .O(N__20807),
            .I(N__20804));
    LocalMux I__2112 (
            .O(N__20804),
            .I(N__20801));
    Span4Mux_v I__2111 (
            .O(N__20801),
            .I(N__20798));
    Span4Mux_h I__2110 (
            .O(N__20798),
            .I(N__20794));
    InMux I__2109 (
            .O(N__20797),
            .I(N__20791));
    Odrv4 I__2108 (
            .O(N__20794),
            .I(\ADC_IAC.n12586 ));
    LocalMux I__2107 (
            .O(N__20791),
            .I(\ADC_IAC.n12586 ));
    SRMux I__2106 (
            .O(N__20786),
            .I(N__20783));
    LocalMux I__2105 (
            .O(N__20783),
            .I(N__20780));
    Span4Mux_h I__2104 (
            .O(N__20780),
            .I(N__20777));
    Odrv4 I__2103 (
            .O(N__20777),
            .I(\ADC_IAC.n14860 ));
    CascadeMux I__2102 (
            .O(N__20774),
            .I(N__20770));
    InMux I__2101 (
            .O(N__20773),
            .I(N__20767));
    InMux I__2100 (
            .O(N__20770),
            .I(N__20764));
    LocalMux I__2099 (
            .O(N__20767),
            .I(cmd_rdadctmp_1_adj_1449));
    LocalMux I__2098 (
            .O(N__20764),
            .I(cmd_rdadctmp_1_adj_1449));
    CascadeMux I__2097 (
            .O(N__20759),
            .I(N__20756));
    InMux I__2096 (
            .O(N__20756),
            .I(N__20752));
    CascadeMux I__2095 (
            .O(N__20755),
            .I(N__20749));
    LocalMux I__2094 (
            .O(N__20752),
            .I(N__20746));
    InMux I__2093 (
            .O(N__20749),
            .I(N__20743));
    Odrv12 I__2092 (
            .O(N__20746),
            .I(cmd_rdadctmp_2_adj_1448));
    LocalMux I__2091 (
            .O(N__20743),
            .I(cmd_rdadctmp_2_adj_1448));
    IoInMux I__2090 (
            .O(N__20738),
            .I(N__20735));
    LocalMux I__2089 (
            .O(N__20735),
            .I(N__20732));
    Span4Mux_s2_v I__2088 (
            .O(N__20732),
            .I(N__20729));
    Span4Mux_v I__2087 (
            .O(N__20729),
            .I(N__20726));
    Span4Mux_h I__2086 (
            .O(N__20726),
            .I(N__20723));
    Odrv4 I__2085 (
            .O(N__20723),
            .I(DDS_MCLK1));
    CascadeMux I__2084 (
            .O(N__20720),
            .I(N__20717));
    InMux I__2083 (
            .O(N__20717),
            .I(N__20714));
    LocalMux I__2082 (
            .O(N__20714),
            .I(N__20711));
    Span4Mux_v I__2081 (
            .O(N__20711),
            .I(N__20707));
    CascadeMux I__2080 (
            .O(N__20710),
            .I(N__20703));
    Span4Mux_v I__2079 (
            .O(N__20707),
            .I(N__20700));
    InMux I__2078 (
            .O(N__20706),
            .I(N__20697));
    InMux I__2077 (
            .O(N__20703),
            .I(N__20694));
    Odrv4 I__2076 (
            .O(N__20700),
            .I(cmd_rdadctmp_28_adj_1422));
    LocalMux I__2075 (
            .O(N__20697),
            .I(cmd_rdadctmp_28_adj_1422));
    LocalMux I__2074 (
            .O(N__20694),
            .I(cmd_rdadctmp_28_adj_1422));
    CascadeMux I__2073 (
            .O(N__20687),
            .I(N__20684));
    InMux I__2072 (
            .O(N__20684),
            .I(N__20678));
    InMux I__2071 (
            .O(N__20683),
            .I(N__20678));
    LocalMux I__2070 (
            .O(N__20678),
            .I(cmd_rdadctmp_3_adj_1447));
    CascadeMux I__2069 (
            .O(N__20675),
            .I(N__20672));
    InMux I__2068 (
            .O(N__20672),
            .I(N__20666));
    InMux I__2067 (
            .O(N__20671),
            .I(N__20663));
    InMux I__2066 (
            .O(N__20670),
            .I(N__20658));
    InMux I__2065 (
            .O(N__20669),
            .I(N__20658));
    LocalMux I__2064 (
            .O(N__20666),
            .I(N__20650));
    LocalMux I__2063 (
            .O(N__20663),
            .I(N__20650));
    LocalMux I__2062 (
            .O(N__20658),
            .I(N__20650));
    CascadeMux I__2061 (
            .O(N__20657),
            .I(N__20647));
    Span4Mux_v I__2060 (
            .O(N__20650),
            .I(N__20644));
    InMux I__2059 (
            .O(N__20647),
            .I(N__20641));
    Sp12to4 I__2058 (
            .O(N__20644),
            .I(N__20636));
    LocalMux I__2057 (
            .O(N__20641),
            .I(N__20636));
    Span12Mux_h I__2056 (
            .O(N__20636),
            .I(N__20633));
    Odrv12 I__2055 (
            .O(N__20633),
            .I(IAC_DRDY));
    InMux I__2054 (
            .O(N__20630),
            .I(N__20627));
    LocalMux I__2053 (
            .O(N__20627),
            .I(n20612));
    CascadeMux I__2052 (
            .O(N__20624),
            .I(n14_adj_1604_cascade_));
    IoInMux I__2051 (
            .O(N__20621),
            .I(N__20618));
    LocalMux I__2050 (
            .O(N__20618),
            .I(N__20615));
    IoSpan4Mux I__2049 (
            .O(N__20615),
            .I(N__20612));
    Sp12to4 I__2048 (
            .O(N__20612),
            .I(N__20608));
    CascadeMux I__2047 (
            .O(N__20611),
            .I(N__20605));
    Span12Mux_v I__2046 (
            .O(N__20608),
            .I(N__20602));
    InMux I__2045 (
            .O(N__20605),
            .I(N__20599));
    Odrv12 I__2044 (
            .O(N__20602),
            .I(IAC_CS));
    LocalMux I__2043 (
            .O(N__20599),
            .I(IAC_CS));
    InMux I__2042 (
            .O(N__20594),
            .I(N__20590));
    InMux I__2041 (
            .O(N__20593),
            .I(N__20587));
    LocalMux I__2040 (
            .O(N__20590),
            .I(\ADC_IAC.bit_cnt_0 ));
    LocalMux I__2039 (
            .O(N__20587),
            .I(\ADC_IAC.bit_cnt_0 ));
    InMux I__2038 (
            .O(N__20582),
            .I(bfn_6_15_0_));
    CascadeMux I__2037 (
            .O(N__20579),
            .I(N__20575));
    InMux I__2036 (
            .O(N__20578),
            .I(N__20572));
    InMux I__2035 (
            .O(N__20575),
            .I(N__20569));
    LocalMux I__2034 (
            .O(N__20572),
            .I(\ADC_IAC.bit_cnt_1 ));
    LocalMux I__2033 (
            .O(N__20569),
            .I(\ADC_IAC.bit_cnt_1 ));
    InMux I__2032 (
            .O(N__20564),
            .I(\ADC_IAC.n19415 ));
    InMux I__2031 (
            .O(N__20561),
            .I(N__20557));
    InMux I__2030 (
            .O(N__20560),
            .I(N__20554));
    LocalMux I__2029 (
            .O(N__20557),
            .I(\ADC_IAC.bit_cnt_2 ));
    LocalMux I__2028 (
            .O(N__20554),
            .I(\ADC_IAC.bit_cnt_2 ));
    InMux I__2027 (
            .O(N__20549),
            .I(\ADC_IAC.n19416 ));
    InMux I__2026 (
            .O(N__20546),
            .I(N__20542));
    InMux I__2025 (
            .O(N__20545),
            .I(N__20539));
    LocalMux I__2024 (
            .O(N__20542),
            .I(\ADC_IAC.bit_cnt_3 ));
    LocalMux I__2023 (
            .O(N__20539),
            .I(\ADC_IAC.bit_cnt_3 ));
    InMux I__2022 (
            .O(N__20534),
            .I(\ADC_IAC.n19417 ));
    CascadeMux I__2021 (
            .O(N__20531),
            .I(N__20528));
    InMux I__2020 (
            .O(N__20528),
            .I(N__20525));
    LocalMux I__2019 (
            .O(N__20525),
            .I(N__20520));
    InMux I__2018 (
            .O(N__20524),
            .I(N__20515));
    InMux I__2017 (
            .O(N__20523),
            .I(N__20515));
    Odrv4 I__2016 (
            .O(N__20520),
            .I(read_buf_13));
    LocalMux I__2015 (
            .O(N__20515),
            .I(read_buf_13));
    InMux I__2014 (
            .O(N__20510),
            .I(N__20507));
    LocalMux I__2013 (
            .O(N__20507),
            .I(N__20502));
    InMux I__2012 (
            .O(N__20506),
            .I(N__20497));
    InMux I__2011 (
            .O(N__20505),
            .I(N__20497));
    Odrv4 I__2010 (
            .O(N__20502),
            .I(read_buf_8));
    LocalMux I__2009 (
            .O(N__20497),
            .I(read_buf_8));
    CascadeMux I__2008 (
            .O(N__20492),
            .I(N__20487));
    CascadeMux I__2007 (
            .O(N__20491),
            .I(N__20483));
    InMux I__2006 (
            .O(N__20490),
            .I(N__20471));
    InMux I__2005 (
            .O(N__20487),
            .I(N__20471));
    InMux I__2004 (
            .O(N__20486),
            .I(N__20471));
    InMux I__2003 (
            .O(N__20483),
            .I(N__20471));
    InMux I__2002 (
            .O(N__20482),
            .I(N__20471));
    LocalMux I__2001 (
            .O(N__20471),
            .I(N__20467));
    InMux I__2000 (
            .O(N__20470),
            .I(N__20464));
    Odrv12 I__1999 (
            .O(N__20467),
            .I(n20754));
    LocalMux I__1998 (
            .O(N__20464),
            .I(n20754));
    InMux I__1997 (
            .O(N__20459),
            .I(N__20455));
    InMux I__1996 (
            .O(N__20458),
            .I(N__20452));
    LocalMux I__1995 (
            .O(N__20455),
            .I(cmd_rdadctmp_5_adj_1445));
    LocalMux I__1994 (
            .O(N__20452),
            .I(cmd_rdadctmp_5_adj_1445));
    CascadeMux I__1993 (
            .O(N__20447),
            .I(N__20444));
    InMux I__1992 (
            .O(N__20444),
            .I(N__20438));
    InMux I__1991 (
            .O(N__20443),
            .I(N__20438));
    LocalMux I__1990 (
            .O(N__20438),
            .I(cmd_rdadctmp_4_adj_1446));
    CascadeMux I__1989 (
            .O(N__20435),
            .I(\RTD.n19_cascade_ ));
    CascadeMux I__1988 (
            .O(N__20432),
            .I(N__20427));
    InMux I__1987 (
            .O(N__20431),
            .I(N__20424));
    InMux I__1986 (
            .O(N__20430),
            .I(N__20419));
    InMux I__1985 (
            .O(N__20427),
            .I(N__20419));
    LocalMux I__1984 (
            .O(N__20424),
            .I(read_buf_9));
    LocalMux I__1983 (
            .O(N__20419),
            .I(read_buf_9));
    CascadeMux I__1982 (
            .O(N__20414),
            .I(N__20411));
    InMux I__1981 (
            .O(N__20411),
            .I(N__20408));
    LocalMux I__1980 (
            .O(N__20408),
            .I(N__20404));
    InMux I__1979 (
            .O(N__20407),
            .I(N__20401));
    Odrv4 I__1978 (
            .O(N__20404),
            .I(adress_1));
    LocalMux I__1977 (
            .O(N__20401),
            .I(adress_1));
    CascadeMux I__1976 (
            .O(N__20396),
            .I(N__20391));
    CascadeMux I__1975 (
            .O(N__20395),
            .I(N__20388));
    InMux I__1974 (
            .O(N__20394),
            .I(N__20381));
    InMux I__1973 (
            .O(N__20391),
            .I(N__20381));
    InMux I__1972 (
            .O(N__20388),
            .I(N__20381));
    LocalMux I__1971 (
            .O(N__20381),
            .I(read_buf_1));
    InMux I__1970 (
            .O(N__20378),
            .I(N__20372));
    InMux I__1969 (
            .O(N__20377),
            .I(N__20372));
    LocalMux I__1968 (
            .O(N__20372),
            .I(adress_2));
    InMux I__1967 (
            .O(N__20369),
            .I(N__20363));
    InMux I__1966 (
            .O(N__20368),
            .I(N__20363));
    LocalMux I__1965 (
            .O(N__20363),
            .I(adress_4));
    CascadeMux I__1964 (
            .O(N__20360),
            .I(N__20357));
    InMux I__1963 (
            .O(N__20357),
            .I(N__20351));
    InMux I__1962 (
            .O(N__20356),
            .I(N__20351));
    LocalMux I__1961 (
            .O(N__20351),
            .I(adress_5));
    IoInMux I__1960 (
            .O(N__20348),
            .I(N__20345));
    LocalMux I__1959 (
            .O(N__20345),
            .I(N__20342));
    Span4Mux_s1_h I__1958 (
            .O(N__20342),
            .I(N__20339));
    Span4Mux_v I__1957 (
            .O(N__20339),
            .I(N__20336));
    Span4Mux_v I__1956 (
            .O(N__20336),
            .I(N__20333));
    Span4Mux_h I__1955 (
            .O(N__20333),
            .I(N__20330));
    Span4Mux_h I__1954 (
            .O(N__20330),
            .I(N__20327));
    Odrv4 I__1953 (
            .O(N__20327),
            .I(RTD_SDI));
    CascadeMux I__1952 (
            .O(N__20324),
            .I(\RTD.n21309_cascade_ ));
    InMux I__1951 (
            .O(N__20321),
            .I(N__20318));
    LocalMux I__1950 (
            .O(N__20318),
            .I(\RTD.n12 ));
    InMux I__1949 (
            .O(N__20315),
            .I(N__20311));
    InMux I__1948 (
            .O(N__20314),
            .I(N__20305));
    LocalMux I__1947 (
            .O(N__20311),
            .I(N__20302));
    InMux I__1946 (
            .O(N__20310),
            .I(N__20299));
    InMux I__1945 (
            .O(N__20309),
            .I(N__20294));
    InMux I__1944 (
            .O(N__20308),
            .I(N__20294));
    LocalMux I__1943 (
            .O(N__20305),
            .I(\ADC_VDC.bit_cnt_2 ));
    Odrv4 I__1942 (
            .O(N__20302),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__1941 (
            .O(N__20299),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__1940 (
            .O(N__20294),
            .I(\ADC_VDC.bit_cnt_2 ));
    InMux I__1939 (
            .O(N__20285),
            .I(N__20282));
    LocalMux I__1938 (
            .O(N__20282),
            .I(\ADC_VDC.n6 ));
    CascadeMux I__1937 (
            .O(N__20279),
            .I(\ADC_VDC.n10552_cascade_ ));
    InMux I__1936 (
            .O(N__20276),
            .I(N__20273));
    LocalMux I__1935 (
            .O(N__20273),
            .I(\ADC_VDC.n21974 ));
    InMux I__1934 (
            .O(N__20270),
            .I(N__20262));
    InMux I__1933 (
            .O(N__20269),
            .I(N__20262));
    CascadeMux I__1932 (
            .O(N__20268),
            .I(N__20259));
    InMux I__1931 (
            .O(N__20267),
            .I(N__20255));
    LocalMux I__1930 (
            .O(N__20262),
            .I(N__20252));
    InMux I__1929 (
            .O(N__20259),
            .I(N__20249));
    InMux I__1928 (
            .O(N__20258),
            .I(N__20246));
    LocalMux I__1927 (
            .O(N__20255),
            .I(\ADC_VDC.bit_cnt_3 ));
    Odrv4 I__1926 (
            .O(N__20252),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__1925 (
            .O(N__20249),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__1924 (
            .O(N__20246),
            .I(\ADC_VDC.bit_cnt_3 ));
    InMux I__1923 (
            .O(N__20237),
            .I(N__20234));
    LocalMux I__1922 (
            .O(N__20234),
            .I(N__20231));
    Odrv4 I__1921 (
            .O(N__20231),
            .I(\ADC_VDC.n20562 ));
    CascadeMux I__1920 (
            .O(N__20228),
            .I(\ADC_VDC.n21224_cascade_ ));
    InMux I__1919 (
            .O(N__20225),
            .I(N__20222));
    LocalMux I__1918 (
            .O(N__20222),
            .I(N__20219));
    Odrv4 I__1917 (
            .O(N__20219),
            .I(\ADC_VDC.n20748 ));
    CascadeMux I__1916 (
            .O(N__20216),
            .I(\ADC_VDC.n31_cascade_ ));
    CEMux I__1915 (
            .O(N__20213),
            .I(N__20210));
    LocalMux I__1914 (
            .O(N__20210),
            .I(N__20207));
    Span4Mux_v I__1913 (
            .O(N__20207),
            .I(N__20204));
    Odrv4 I__1912 (
            .O(N__20204),
            .I(\ADC_VDC.n20555 ));
    CascadeMux I__1911 (
            .O(N__20201),
            .I(N__20198));
    InMux I__1910 (
            .O(N__20198),
            .I(N__20193));
    InMux I__1909 (
            .O(N__20197),
            .I(N__20188));
    InMux I__1908 (
            .O(N__20196),
            .I(N__20188));
    LocalMux I__1907 (
            .O(N__20193),
            .I(read_buf_12));
    LocalMux I__1906 (
            .O(N__20188),
            .I(read_buf_12));
    CascadeMux I__1905 (
            .O(N__20183),
            .I(N__20180));
    InMux I__1904 (
            .O(N__20180),
            .I(N__20174));
    InMux I__1903 (
            .O(N__20179),
            .I(N__20174));
    LocalMux I__1902 (
            .O(N__20174),
            .I(adress_3));
    InMux I__1901 (
            .O(N__20171),
            .I(N__20166));
    InMux I__1900 (
            .O(N__20170),
            .I(N__20163));
    InMux I__1899 (
            .O(N__20169),
            .I(N__20160));
    LocalMux I__1898 (
            .O(N__20166),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__1897 (
            .O(N__20163),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__1896 (
            .O(N__20160),
            .I(\ADC_VDC.bit_cnt_5 ));
    CascadeMux I__1895 (
            .O(N__20153),
            .I(\ADC_VDC.n20534_cascade_ ));
    InMux I__1894 (
            .O(N__20150),
            .I(N__20147));
    LocalMux I__1893 (
            .O(N__20147),
            .I(\ADC_VDC.n10 ));
    InMux I__1892 (
            .O(N__20144),
            .I(N__20139));
    InMux I__1891 (
            .O(N__20143),
            .I(N__20134));
    InMux I__1890 (
            .O(N__20142),
            .I(N__20134));
    LocalMux I__1889 (
            .O(N__20139),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__1888 (
            .O(N__20134),
            .I(\ADC_VDC.bit_cnt_7 ));
    InMux I__1887 (
            .O(N__20129),
            .I(N__20124));
    InMux I__1886 (
            .O(N__20128),
            .I(N__20119));
    InMux I__1885 (
            .O(N__20127),
            .I(N__20119));
    LocalMux I__1884 (
            .O(N__20124),
            .I(\ADC_VDC.bit_cnt_6 ));
    LocalMux I__1883 (
            .O(N__20119),
            .I(\ADC_VDC.bit_cnt_6 ));
    InMux I__1882 (
            .O(N__20114),
            .I(N__20111));
    LocalMux I__1881 (
            .O(N__20111),
            .I(\ADC_VDC.n21082 ));
    CascadeMux I__1880 (
            .O(N__20108),
            .I(N__20105));
    InMux I__1879 (
            .O(N__20105),
            .I(N__20102));
    LocalMux I__1878 (
            .O(N__20102),
            .I(N__20099));
    Odrv4 I__1877 (
            .O(N__20099),
            .I(\ADC_VDC.n21079 ));
    CascadeMux I__1876 (
            .O(N__20096),
            .I(\ADC_VDC.n21977_cascade_ ));
    InMux I__1875 (
            .O(N__20093),
            .I(N__20090));
    LocalMux I__1874 (
            .O(N__20090),
            .I(\ADC_VDC.n18482 ));
    InMux I__1873 (
            .O(N__20087),
            .I(bfn_6_6_0_));
    InMux I__1872 (
            .O(N__20084),
            .I(\ADC_VDC.n19531 ));
    InMux I__1871 (
            .O(N__20081),
            .I(\ADC_VDC.n19532 ));
    InMux I__1870 (
            .O(N__20078),
            .I(\ADC_VDC.n19533 ));
    InMux I__1869 (
            .O(N__20075),
            .I(\ADC_VDC.n19534 ));
    InMux I__1868 (
            .O(N__20072),
            .I(\ADC_VDC.n19535 ));
    InMux I__1867 (
            .O(N__20069),
            .I(\ADC_VDC.n19536 ));
    InMux I__1866 (
            .O(N__20066),
            .I(\ADC_VDC.n19537 ));
    CascadeMux I__1865 (
            .O(N__20063),
            .I(\ADC_IAC.n21068_cascade_ ));
    CEMux I__1864 (
            .O(N__20060),
            .I(N__20057));
    LocalMux I__1863 (
            .O(N__20057),
            .I(N__20054));
    Odrv4 I__1862 (
            .O(N__20054),
            .I(\ADC_IAC.n20714 ));
    CascadeMux I__1861 (
            .O(N__20051),
            .I(N__20048));
    InMux I__1860 (
            .O(N__20048),
            .I(N__20045));
    LocalMux I__1859 (
            .O(N__20045),
            .I(N__20042));
    Span4Mux_v I__1858 (
            .O(N__20042),
            .I(N__20039));
    Span4Mux_v I__1857 (
            .O(N__20039),
            .I(N__20036));
    IoSpan4Mux I__1856 (
            .O(N__20036),
            .I(N__20033));
    Odrv4 I__1855 (
            .O(N__20033),
            .I(IAC_MISO));
    InMux I__1854 (
            .O(N__20030),
            .I(N__20024));
    InMux I__1853 (
            .O(N__20029),
            .I(N__20024));
    LocalMux I__1852 (
            .O(N__20024),
            .I(cmd_rdadctmp_0_adj_1450));
    IoInMux I__1851 (
            .O(N__20021),
            .I(N__20018));
    LocalMux I__1850 (
            .O(N__20018),
            .I(N__20015));
    Span4Mux_s2_v I__1849 (
            .O(N__20015),
            .I(N__20012));
    Span4Mux_v I__1848 (
            .O(N__20012),
            .I(N__20008));
    CascadeMux I__1847 (
            .O(N__20011),
            .I(N__20005));
    Span4Mux_v I__1846 (
            .O(N__20008),
            .I(N__20002));
    InMux I__1845 (
            .O(N__20005),
            .I(N__19999));
    Odrv4 I__1844 (
            .O(N__20002),
            .I(IAC_SCLK));
    LocalMux I__1843 (
            .O(N__19999),
            .I(IAC_SCLK));
    CascadeMux I__1842 (
            .O(N__19994),
            .I(N__19989));
    CascadeMux I__1841 (
            .O(N__19993),
            .I(N__19986));
    CascadeMux I__1840 (
            .O(N__19992),
            .I(N__19983));
    InMux I__1839 (
            .O(N__19989),
            .I(N__19980));
    InMux I__1838 (
            .O(N__19986),
            .I(N__19975));
    InMux I__1837 (
            .O(N__19983),
            .I(N__19975));
    LocalMux I__1836 (
            .O(N__19980),
            .I(cmd_rdadctmp_28));
    LocalMux I__1835 (
            .O(N__19975),
            .I(cmd_rdadctmp_28));
    CEMux I__1834 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__1833 (
            .O(N__19967),
            .I(N__19964));
    Span4Mux_v I__1832 (
            .O(N__19964),
            .I(N__19961));
    Span4Mux_h I__1831 (
            .O(N__19961),
            .I(N__19958));
    Odrv4 I__1830 (
            .O(N__19958),
            .I(\ADC_IAC.n12 ));
    CascadeMux I__1829 (
            .O(N__19955),
            .I(n20612_cascade_));
    InMux I__1828 (
            .O(N__19952),
            .I(N__19949));
    LocalMux I__1827 (
            .O(N__19949),
            .I(\ADC_IAC.n20713 ));
    CascadeMux I__1826 (
            .O(N__19946),
            .I(\ADC_IAC.n20783_cascade_ ));
    CascadeMux I__1825 (
            .O(N__19943),
            .I(\ADC_IAC.n20795_cascade_ ));
    CascadeMux I__1824 (
            .O(N__19940),
            .I(N__19937));
    InMux I__1823 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__1822 (
            .O(N__19934),
            .I(N__19931));
    Odrv12 I__1821 (
            .O(N__19931),
            .I(\CLK_DDS.tmp_buf_0 ));
    CascadeMux I__1820 (
            .O(N__19928),
            .I(N__19924));
    InMux I__1819 (
            .O(N__19927),
            .I(N__19921));
    InMux I__1818 (
            .O(N__19924),
            .I(N__19918));
    LocalMux I__1817 (
            .O(N__19921),
            .I(N__19915));
    LocalMux I__1816 (
            .O(N__19918),
            .I(bit_cnt_3));
    Odrv4 I__1815 (
            .O(N__19915),
            .I(bit_cnt_3));
    InMux I__1814 (
            .O(N__19910),
            .I(N__19901));
    InMux I__1813 (
            .O(N__19909),
            .I(N__19901));
    InMux I__1812 (
            .O(N__19908),
            .I(N__19901));
    LocalMux I__1811 (
            .O(N__19901),
            .I(N__19896));
    InMux I__1810 (
            .O(N__19900),
            .I(N__19891));
    InMux I__1809 (
            .O(N__19899),
            .I(N__19891));
    Odrv4 I__1808 (
            .O(N__19896),
            .I(bit_cnt_0_adj_1456));
    LocalMux I__1807 (
            .O(N__19891),
            .I(bit_cnt_0_adj_1456));
    CascadeMux I__1806 (
            .O(N__19886),
            .I(\ADC_IAC.n17_cascade_ ));
    IoInMux I__1805 (
            .O(N__19883),
            .I(N__19880));
    LocalMux I__1804 (
            .O(N__19880),
            .I(N__19877));
    IoSpan4Mux I__1803 (
            .O(N__19877),
            .I(N__19874));
    Span4Mux_s2_v I__1802 (
            .O(N__19874),
            .I(N__19871));
    Sp12to4 I__1801 (
            .O(N__19871),
            .I(N__19867));
    CascadeMux I__1800 (
            .O(N__19870),
            .I(N__19864));
    Span12Mux_s11_v I__1799 (
            .O(N__19867),
            .I(N__19861));
    InMux I__1798 (
            .O(N__19864),
            .I(N__19858));
    Odrv12 I__1797 (
            .O(N__19861),
            .I(DDS_SCK1));
    LocalMux I__1796 (
            .O(N__19858),
            .I(DDS_SCK1));
    CascadeMux I__1795 (
            .O(N__19853),
            .I(N__19849));
    InMux I__1794 (
            .O(N__19852),
            .I(N__19844));
    InMux I__1793 (
            .O(N__19849),
            .I(N__19844));
    LocalMux I__1792 (
            .O(N__19844),
            .I(cmd_rdadctmp_6_adj_1444));
    IoInMux I__1791 (
            .O(N__19841),
            .I(N__19838));
    LocalMux I__1790 (
            .O(N__19838),
            .I(N__19835));
    Span4Mux_s2_v I__1789 (
            .O(N__19835),
            .I(N__19832));
    Span4Mux_v I__1788 (
            .O(N__19832),
            .I(N__19829));
    Span4Mux_v I__1787 (
            .O(N__19829),
            .I(N__19826));
    Span4Mux_v I__1786 (
            .O(N__19826),
            .I(N__19823));
    Odrv4 I__1785 (
            .O(N__19823),
            .I(DDS_CS1));
    InMux I__1784 (
            .O(N__19820),
            .I(N__19817));
    LocalMux I__1783 (
            .O(N__19817),
            .I(N__19814));
    Span12Mux_h I__1782 (
            .O(N__19814),
            .I(N__19811));
    Span12Mux_v I__1781 (
            .O(N__19811),
            .I(N__19808));
    Odrv12 I__1780 (
            .O(N__19808),
            .I(RTD_SDO));
    InMux I__1779 (
            .O(N__19805),
            .I(\ADC_VDC.n19466 ));
    InMux I__1778 (
            .O(N__19802),
            .I(\ADC_VDC.n19467 ));
    InMux I__1777 (
            .O(N__19799),
            .I(N__19795));
    InMux I__1776 (
            .O(N__19798),
            .I(N__19792));
    LocalMux I__1775 (
            .O(N__19795),
            .I(N__19789));
    LocalMux I__1774 (
            .O(N__19792),
            .I(\ADC_VDC.avg_cnt_4 ));
    Odrv4 I__1773 (
            .O(N__19789),
            .I(\ADC_VDC.avg_cnt_4 ));
    InMux I__1772 (
            .O(N__19784),
            .I(N__19780));
    InMux I__1771 (
            .O(N__19783),
            .I(N__19777));
    LocalMux I__1770 (
            .O(N__19780),
            .I(N__19774));
    LocalMux I__1769 (
            .O(N__19777),
            .I(\ADC_VDC.avg_cnt_7 ));
    Odrv4 I__1768 (
            .O(N__19774),
            .I(\ADC_VDC.avg_cnt_7 ));
    CascadeMux I__1767 (
            .O(N__19769),
            .I(N__19766));
    InMux I__1766 (
            .O(N__19766),
            .I(N__19762));
    InMux I__1765 (
            .O(N__19765),
            .I(N__19759));
    LocalMux I__1764 (
            .O(N__19762),
            .I(N__19756));
    LocalMux I__1763 (
            .O(N__19759),
            .I(\ADC_VDC.avg_cnt_3 ));
    Odrv4 I__1762 (
            .O(N__19756),
            .I(\ADC_VDC.avg_cnt_3 ));
    InMux I__1761 (
            .O(N__19751),
            .I(N__19747));
    InMux I__1760 (
            .O(N__19750),
            .I(N__19744));
    LocalMux I__1759 (
            .O(N__19747),
            .I(N__19741));
    LocalMux I__1758 (
            .O(N__19744),
            .I(\ADC_VDC.avg_cnt_5 ));
    Odrv4 I__1757 (
            .O(N__19741),
            .I(\ADC_VDC.avg_cnt_5 ));
    InMux I__1756 (
            .O(N__19736),
            .I(N__19732));
    InMux I__1755 (
            .O(N__19735),
            .I(N__19729));
    LocalMux I__1754 (
            .O(N__19732),
            .I(N__19726));
    LocalMux I__1753 (
            .O(N__19729),
            .I(\ADC_VDC.avg_cnt_9 ));
    Odrv12 I__1752 (
            .O(N__19726),
            .I(\ADC_VDC.avg_cnt_9 ));
    InMux I__1751 (
            .O(N__19721),
            .I(N__19717));
    InMux I__1750 (
            .O(N__19720),
            .I(N__19714));
    LocalMux I__1749 (
            .O(N__19717),
            .I(N__19711));
    LocalMux I__1748 (
            .O(N__19714),
            .I(\ADC_VDC.avg_cnt_0 ));
    Odrv12 I__1747 (
            .O(N__19711),
            .I(\ADC_VDC.avg_cnt_0 ));
    CascadeMux I__1746 (
            .O(N__19706),
            .I(N__19703));
    InMux I__1745 (
            .O(N__19703),
            .I(N__19699));
    InMux I__1744 (
            .O(N__19702),
            .I(N__19696));
    LocalMux I__1743 (
            .O(N__19699),
            .I(N__19693));
    LocalMux I__1742 (
            .O(N__19696),
            .I(\ADC_VDC.avg_cnt_8 ));
    Odrv4 I__1741 (
            .O(N__19693),
            .I(\ADC_VDC.avg_cnt_8 ));
    InMux I__1740 (
            .O(N__19688),
            .I(N__19684));
    InMux I__1739 (
            .O(N__19687),
            .I(N__19681));
    LocalMux I__1738 (
            .O(N__19684),
            .I(N__19678));
    LocalMux I__1737 (
            .O(N__19681),
            .I(\ADC_VDC.avg_cnt_10 ));
    Odrv4 I__1736 (
            .O(N__19678),
            .I(\ADC_VDC.avg_cnt_10 ));
    InMux I__1735 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__1734 (
            .O(N__19670),
            .I(\ADC_VDC.n20 ));
    CascadeMux I__1733 (
            .O(N__19667),
            .I(\ADC_VDC.n19_adj_1412_cascade_ ));
    CascadeMux I__1732 (
            .O(N__19664),
            .I(\ADC_VDC.n18479_cascade_ ));
    InMux I__1731 (
            .O(N__19661),
            .I(\ADC_VDC.n19457 ));
    InMux I__1730 (
            .O(N__19658),
            .I(\ADC_VDC.n19458 ));
    InMux I__1729 (
            .O(N__19655),
            .I(\ADC_VDC.n19459 ));
    InMux I__1728 (
            .O(N__19652),
            .I(\ADC_VDC.n19460 ));
    InMux I__1727 (
            .O(N__19649),
            .I(\ADC_VDC.n19461 ));
    InMux I__1726 (
            .O(N__19646),
            .I(\ADC_VDC.n19462 ));
    InMux I__1725 (
            .O(N__19643),
            .I(\ADC_VDC.n19463 ));
    InMux I__1724 (
            .O(N__19640),
            .I(bfn_5_6_0_));
    InMux I__1723 (
            .O(N__19637),
            .I(\ADC_VDC.n19465 ));
    InMux I__1722 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__1721 (
            .O(N__19631),
            .I(n20615));
    CascadeMux I__1720 (
            .O(N__19628),
            .I(N__19623));
    CascadeMux I__1719 (
            .O(N__19627),
            .I(N__19620));
    CascadeMux I__1718 (
            .O(N__19626),
            .I(N__19617));
    InMux I__1717 (
            .O(N__19623),
            .I(N__19610));
    InMux I__1716 (
            .O(N__19620),
            .I(N__19610));
    InMux I__1715 (
            .O(N__19617),
            .I(N__19610));
    LocalMux I__1714 (
            .O(N__19610),
            .I(N__19605));
    InMux I__1713 (
            .O(N__19609),
            .I(N__19600));
    InMux I__1712 (
            .O(N__19608),
            .I(N__19600));
    Span4Mux_v I__1711 (
            .O(N__19605),
            .I(N__19595));
    LocalMux I__1710 (
            .O(N__19600),
            .I(N__19595));
    Span4Mux_v I__1709 (
            .O(N__19595),
            .I(N__19592));
    Span4Mux_h I__1708 (
            .O(N__19592),
            .I(N__19589));
    Odrv4 I__1707 (
            .O(N__19589),
            .I(VAC_DRDY));
    CascadeMux I__1706 (
            .O(N__19586),
            .I(n20615_cascade_));
    InMux I__1705 (
            .O(N__19583),
            .I(N__19576));
    InMux I__1704 (
            .O(N__19582),
            .I(N__19576));
    InMux I__1703 (
            .O(N__19581),
            .I(N__19573));
    LocalMux I__1702 (
            .O(N__19576),
            .I(bit_cnt_2));
    LocalMux I__1701 (
            .O(N__19573),
            .I(bit_cnt_2));
    CascadeMux I__1700 (
            .O(N__19568),
            .I(N__19563));
    CascadeMux I__1699 (
            .O(N__19567),
            .I(N__19559));
    InMux I__1698 (
            .O(N__19566),
            .I(N__19552));
    InMux I__1697 (
            .O(N__19563),
            .I(N__19552));
    InMux I__1696 (
            .O(N__19562),
            .I(N__19552));
    InMux I__1695 (
            .O(N__19559),
            .I(N__19549));
    LocalMux I__1694 (
            .O(N__19552),
            .I(bit_cnt_1));
    LocalMux I__1693 (
            .O(N__19549),
            .I(bit_cnt_1));
    SRMux I__1692 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__1691 (
            .O(N__19541),
            .I(N__19538));
    Span4Mux_h I__1690 (
            .O(N__19538),
            .I(N__19535));
    Odrv4 I__1689 (
            .O(N__19535),
            .I(\CLK_DDS.n16766 ));
    InMux I__1688 (
            .O(N__19532),
            .I(bfn_5_5_0_));
    CascadeMux I__1687 (
            .O(N__19529),
            .I(\ADC_VAC.n20715_cascade_ ));
    InMux I__1686 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__1685 (
            .O(N__19523),
            .I(\ADC_VAC.n21053 ));
    CEMux I__1684 (
            .O(N__19520),
            .I(N__19517));
    LocalMux I__1683 (
            .O(N__19517),
            .I(\ADC_VAC.n20716 ));
    CascadeMux I__1682 (
            .O(N__19514),
            .I(\ADC_VAC.n17_cascade_ ));
    CEMux I__1681 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__1680 (
            .O(N__19508),
            .I(N__19505));
    Span4Mux_h I__1679 (
            .O(N__19505),
            .I(N__19502));
    Odrv4 I__1678 (
            .O(N__19502),
            .I(\ADC_VAC.n12 ));
    CEMux I__1677 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__1676 (
            .O(N__19496),
            .I(N__19492));
    InMux I__1675 (
            .O(N__19495),
            .I(N__19489));
    Span4Mux_h I__1674 (
            .O(N__19492),
            .I(N__19486));
    LocalMux I__1673 (
            .O(N__19489),
            .I(N__19483));
    Odrv4 I__1672 (
            .O(N__19486),
            .I(\ADC_VAC.n12489 ));
    Odrv4 I__1671 (
            .O(N__19483),
            .I(\ADC_VAC.n12489 ));
    IoInMux I__1670 (
            .O(N__19478),
            .I(N__19475));
    LocalMux I__1669 (
            .O(N__19475),
            .I(N__19472));
    IoSpan4Mux I__1668 (
            .O(N__19472),
            .I(N__19469));
    Span4Mux_s2_h I__1667 (
            .O(N__19469),
            .I(N__19465));
    CascadeMux I__1666 (
            .O(N__19468),
            .I(N__19462));
    Span4Mux_h I__1665 (
            .O(N__19465),
            .I(N__19459));
    InMux I__1664 (
            .O(N__19462),
            .I(N__19456));
    Odrv4 I__1663 (
            .O(N__19459),
            .I(VAC_SCLK));
    LocalMux I__1662 (
            .O(N__19456),
            .I(VAC_SCLK));
    CascadeMux I__1661 (
            .O(N__19451),
            .I(n14_adj_1606_cascade_));
    IoInMux I__1660 (
            .O(N__19448),
            .I(N__19445));
    LocalMux I__1659 (
            .O(N__19445),
            .I(N__19442));
    Span4Mux_s2_h I__1658 (
            .O(N__19442),
            .I(N__19439));
    Span4Mux_h I__1657 (
            .O(N__19439),
            .I(N__19435));
    CascadeMux I__1656 (
            .O(N__19438),
            .I(N__19432));
    Sp12to4 I__1655 (
            .O(N__19435),
            .I(N__19429));
    InMux I__1654 (
            .O(N__19432),
            .I(N__19426));
    Odrv12 I__1653 (
            .O(N__19429),
            .I(VAC_CS));
    LocalMux I__1652 (
            .O(N__19426),
            .I(VAC_CS));
    InMux I__1651 (
            .O(N__19421),
            .I(N__19417));
    InMux I__1650 (
            .O(N__19420),
            .I(N__19414));
    LocalMux I__1649 (
            .O(N__19417),
            .I(\ADC_VAC.bit_cnt_7 ));
    LocalMux I__1648 (
            .O(N__19414),
            .I(\ADC_VAC.bit_cnt_7 ));
    InMux I__1647 (
            .O(N__19409),
            .I(N__19405));
    InMux I__1646 (
            .O(N__19408),
            .I(N__19402));
    LocalMux I__1645 (
            .O(N__19405),
            .I(\ADC_VAC.bit_cnt_1 ));
    LocalMux I__1644 (
            .O(N__19402),
            .I(\ADC_VAC.bit_cnt_1 ));
    CascadeMux I__1643 (
            .O(N__19397),
            .I(\ADC_VAC.n21054_cascade_ ));
    InMux I__1642 (
            .O(N__19394),
            .I(N__19391));
    LocalMux I__1641 (
            .O(N__19391),
            .I(\ADC_VAC.n16 ));
    CascadeMux I__1640 (
            .O(N__19388),
            .I(N__19385));
    InMux I__1639 (
            .O(N__19385),
            .I(N__19382));
    LocalMux I__1638 (
            .O(N__19382),
            .I(N__19379));
    Span4Mux_h I__1637 (
            .O(N__19379),
            .I(N__19376));
    Span4Mux_v I__1636 (
            .O(N__19376),
            .I(N__19373));
    Span4Mux_v I__1635 (
            .O(N__19373),
            .I(N__19370));
    Odrv4 I__1634 (
            .O(N__19370),
            .I(VAC_MISO));
    InMux I__1633 (
            .O(N__19367),
            .I(N__19361));
    InMux I__1632 (
            .O(N__19366),
            .I(N__19361));
    LocalMux I__1631 (
            .O(N__19361),
            .I(cmd_rdadctmp_0));
    CascadeMux I__1630 (
            .O(N__19358),
            .I(N__19355));
    InMux I__1629 (
            .O(N__19355),
            .I(N__19351));
    InMux I__1628 (
            .O(N__19354),
            .I(N__19348));
    LocalMux I__1627 (
            .O(N__19351),
            .I(cmd_rdadctmp_1));
    LocalMux I__1626 (
            .O(N__19348),
            .I(cmd_rdadctmp_1));
    InMux I__1625 (
            .O(N__19343),
            .I(N__19337));
    InMux I__1624 (
            .O(N__19342),
            .I(N__19337));
    LocalMux I__1623 (
            .O(N__19337),
            .I(cmd_rdadctmp_2));
    CascadeMux I__1622 (
            .O(N__19334),
            .I(N__19330));
    InMux I__1621 (
            .O(N__19333),
            .I(N__19325));
    InMux I__1620 (
            .O(N__19330),
            .I(N__19325));
    LocalMux I__1619 (
            .O(N__19325),
            .I(cmd_rdadctmp_3));
    SRMux I__1618 (
            .O(N__19322),
            .I(N__19319));
    LocalMux I__1617 (
            .O(N__19319),
            .I(N__19316));
    Span4Mux_h I__1616 (
            .O(N__19316),
            .I(N__19313));
    Span4Mux_s3_h I__1615 (
            .O(N__19313),
            .I(N__19310));
    Odrv4 I__1614 (
            .O(N__19310),
            .I(\ADC_VAC.n14822 ));
    InMux I__1613 (
            .O(N__19307),
            .I(\ADC_VAC.n19408 ));
    InMux I__1612 (
            .O(N__19304),
            .I(\ADC_VAC.n19409 ));
    InMux I__1611 (
            .O(N__19301),
            .I(\ADC_VAC.n19410 ));
    InMux I__1610 (
            .O(N__19298),
            .I(\ADC_VAC.n19411 ));
    InMux I__1609 (
            .O(N__19295),
            .I(\ADC_VAC.n19412 ));
    InMux I__1608 (
            .O(N__19292),
            .I(\ADC_VAC.n19413 ));
    InMux I__1607 (
            .O(N__19289),
            .I(\ADC_VAC.n19414 ));
    InMux I__1606 (
            .O(N__19286),
            .I(N__19282));
    InMux I__1605 (
            .O(N__19285),
            .I(N__19279));
    LocalMux I__1604 (
            .O(N__19282),
            .I(\ADC_VAC.bit_cnt_0 ));
    LocalMux I__1603 (
            .O(N__19279),
            .I(\ADC_VAC.bit_cnt_0 ));
    CascadeMux I__1602 (
            .O(N__19274),
            .I(N__19270));
    InMux I__1601 (
            .O(N__19273),
            .I(N__19267));
    InMux I__1600 (
            .O(N__19270),
            .I(N__19264));
    LocalMux I__1599 (
            .O(N__19267),
            .I(\ADC_VAC.bit_cnt_6 ));
    LocalMux I__1598 (
            .O(N__19264),
            .I(\ADC_VAC.bit_cnt_6 ));
    InMux I__1597 (
            .O(N__19259),
            .I(N__19255));
    InMux I__1596 (
            .O(N__19258),
            .I(N__19252));
    LocalMux I__1595 (
            .O(N__19255),
            .I(\ADC_VAC.bit_cnt_4 ));
    LocalMux I__1594 (
            .O(N__19252),
            .I(\ADC_VAC.bit_cnt_4 ));
    InMux I__1593 (
            .O(N__19247),
            .I(N__19243));
    InMux I__1592 (
            .O(N__19246),
            .I(N__19240));
    LocalMux I__1591 (
            .O(N__19243),
            .I(\ADC_VAC.bit_cnt_3 ));
    LocalMux I__1590 (
            .O(N__19240),
            .I(\ADC_VAC.bit_cnt_3 ));
    CascadeMux I__1589 (
            .O(N__19235),
            .I(N__19231));
    InMux I__1588 (
            .O(N__19234),
            .I(N__19228));
    InMux I__1587 (
            .O(N__19231),
            .I(N__19225));
    LocalMux I__1586 (
            .O(N__19228),
            .I(\ADC_VAC.bit_cnt_5 ));
    LocalMux I__1585 (
            .O(N__19225),
            .I(\ADC_VAC.bit_cnt_5 ));
    InMux I__1584 (
            .O(N__19220),
            .I(N__19216));
    InMux I__1583 (
            .O(N__19219),
            .I(N__19213));
    LocalMux I__1582 (
            .O(N__19216),
            .I(\ADC_VAC.bit_cnt_2 ));
    LocalMux I__1581 (
            .O(N__19213),
            .I(\ADC_VAC.bit_cnt_2 ));
    InMux I__1580 (
            .O(N__19208),
            .I(bfn_2_7_0_));
    IoInMux I__1579 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__1578 (
            .O(N__19202),
            .I(N__19199));
    IoSpan4Mux I__1577 (
            .O(N__19199),
            .I(N__19196));
    IoSpan4Mux I__1576 (
            .O(N__19196),
            .I(N__19193));
    Odrv4 I__1575 (
            .O(N__19193),
            .I(ICE_SYSCLK));
    IoInMux I__1574 (
            .O(N__19190),
            .I(N__19187));
    LocalMux I__1573 (
            .O(N__19187),
            .I(N__19184));
    IoSpan4Mux I__1572 (
            .O(N__19184),
            .I(N__19181));
    Span4Mux_s3_v I__1571 (
            .O(N__19181),
            .I(N__19178));
    Sp12to4 I__1570 (
            .O(N__19178),
            .I(N__19175));
    Span12Mux_h I__1569 (
            .O(N__19175),
            .I(N__19172));
    Odrv12 I__1568 (
            .O(N__19172),
            .I(ICE_GPMO_2));
    INV \INVcomm_spi.imiso_83_12208_12209_resetC  (
            .O(\INVcomm_spi.imiso_83_12208_12209_resetC_net ),
            .I(N__56995));
    INV \INVcomm_spi.MISO_48_12202_12203_setC  (
            .O(\INVcomm_spi.MISO_48_12202_12203_setC_net ),
            .I(N__57904));
    INV \INVcomm_spi.MISO_48_12202_12203_resetC  (
            .O(\INVcomm_spi.MISO_48_12202_12203_resetC_net ),
            .I(N__57892));
    INV \INVcomm_spi.imiso_83_12208_12209_setC  (
            .O(\INVcomm_spi.imiso_83_12208_12209_setC_net ),
            .I(N__56998));
    INV \INVcomm_spi.bit_cnt_3778__i3C  (
            .O(\INVcomm_spi.bit_cnt_3778__i3C_net ),
            .I(N__57036));
    INV INVdds0_mclk_304C (
            .O(INVdds0_mclk_304C_net),
            .I(N__45085));
    INV INVdata_cntvec_i0_i8C (
            .O(INVdata_cntvec_i0_i8C_net),
            .I(N__57916));
    INV INVdata_cntvec_i0_i0C (
            .O(INVdata_cntvec_i0_i0C_net),
            .I(N__57899));
    INV \INVcomm_spi.data_valid_85C  (
            .O(\INVcomm_spi.data_valid_85C_net ),
            .I(N__57834));
    INV \INVADC_VDC.genclk.t_clk_24C  (
            .O(\INVADC_VDC.genclk.t_clk_24C_net ),
            .I(N__45079));
    INV INVdds0_mclkcnt_i7_3783__i0C (
            .O(INVdds0_mclkcnt_i7_3783__i0C_net),
            .I(N__45082));
    INV INVeis_state_i2C (
            .O(INVeis_state_i2C_net),
            .I(N__57872));
    INV \INVADC_VDC.genclk.t0on_i8C  (
            .O(\INVADC_VDC.genclk.t0on_i8C_net ),
            .I(N__45078));
    INV \INVADC_VDC.genclk.t0on_i0C  (
            .O(\INVADC_VDC.genclk.t0on_i0C_net ),
            .I(N__45074));
    INV \INVADC_VDC.genclk.div_state_i1C  (
            .O(\INVADC_VDC.genclk.div_state_i1C_net ),
            .I(N__45073));
    INV \INVADC_VDC.genclk.div_state_i0C  (
            .O(\INVADC_VDC.genclk.div_state_i0C_net ),
            .I(N__45072));
    INV INVacadc_skipcnt_i0_i9C (
            .O(INVacadc_skipcnt_i0_i9C_net),
            .I(N__57922));
    INV INVacadc_skipcnt_i0_i1C (
            .O(INVacadc_skipcnt_i0_i1C_net),
            .I(N__57909));
    INV INVacadc_skipcnt_i0_i0C (
            .O(INVacadc_skipcnt_i0_i0C_net),
            .I(N__57894));
    INV INVeis_state_i0C (
            .O(INVeis_state_i0C_net),
            .I(N__57868));
    INV INVeis_end_309C (
            .O(INVeis_end_309C_net),
            .I(N__57859));
    INV \INVADC_VDC.genclk.t0off_i8C  (
            .O(\INVADC_VDC.genclk.t0off_i8C_net ),
            .I(N__45071));
    INV \INVADC_VDC.genclk.t0off_i0C  (
            .O(\INVADC_VDC.genclk.t0off_i0C_net ),
            .I(N__45070));
    INV INVdata_count_i0_i8C (
            .O(INVdata_count_i0_i8C_net),
            .I(N__57861));
    INV INVdata_count_i0_i0C (
            .O(INVdata_count_i0_i0C_net),
            .I(N__57851));
    INV INViac_raw_buf_vac_raw_buf_merged2WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .I(N__57932));
    INV INViac_raw_buf_vac_raw_buf_merged7WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .I(N__57983));
    INV INViac_raw_buf_vac_raw_buf_merged1WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .I(N__57857));
    INV INViac_raw_buf_vac_raw_buf_merged6WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .I(N__57981));
    INV INViac_raw_buf_vac_raw_buf_merged0WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .I(N__57838));
    INV INViac_raw_buf_vac_raw_buf_merged5WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .I(N__57978));
    INV INViac_raw_buf_vac_raw_buf_merged9WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .I(N__57847));
    INV INViac_raw_buf_vac_raw_buf_merged4WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .I(N__57969));
    INV INViac_raw_buf_vac_raw_buf_merged8WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .I(N__57828));
    INV INViac_raw_buf_vac_raw_buf_merged10WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .I(N__57878));
    INV INViac_raw_buf_vac_raw_buf_merged3WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .I(N__57955));
    INV INViac_raw_buf_vac_raw_buf_merged11WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .I(N__57906));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(n19516),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(n19524),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(n19369_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(n19377),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(n19361),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(n19352),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(n19400),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(n19391),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_3_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(\ADC_VDC.genclk.n19475 ),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_13_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_5_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(\ADC_VDC.genclk.n19490 ),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(\ADC_VDC.n19464 ),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_10_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_5_0_));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(\ADC_VDC.n19429 ),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(\ADC_VDC.n19437 ),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(\ADC_VDC.n19445 ),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\ADC_VDC.n19453 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \ADC_VAC.bit_cnt_i0_LC_2_7_0 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i0_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i0_LC_2_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i0_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__19286),
            .in2(_gnd_net_),
            .in3(N__19208),
            .lcout(\ADC_VAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\ADC_VAC.n19408 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i1_LC_2_7_1 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i1_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i1_LC_2_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i1_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__19408),
            .in2(_gnd_net_),
            .in3(N__19307),
            .lcout(\ADC_VAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC.n19408 ),
            .carryout(\ADC_VAC.n19409 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i2_LC_2_7_2 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i2_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i2_LC_2_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i2_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__19220),
            .in2(_gnd_net_),
            .in3(N__19304),
            .lcout(\ADC_VAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC.n19409 ),
            .carryout(\ADC_VAC.n19410 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i3_LC_2_7_3 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i3_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i3_LC_2_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i3_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__19247),
            .in2(_gnd_net_),
            .in3(N__19301),
            .lcout(\ADC_VAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC.n19410 ),
            .carryout(\ADC_VAC.n19411 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i4_LC_2_7_4 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i4_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i4_LC_2_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i4_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__19259),
            .in2(_gnd_net_),
            .in3(N__19298),
            .lcout(\ADC_VAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC.n19411 ),
            .carryout(\ADC_VAC.n19412 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i5_LC_2_7_5 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i5_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i5_LC_2_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i5_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__19234),
            .in2(_gnd_net_),
            .in3(N__19295),
            .lcout(\ADC_VAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC.n19412 ),
            .carryout(\ADC_VAC.n19413 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i6_LC_2_7_6 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i6_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i6_LC_2_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i6_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__19273),
            .in2(_gnd_net_),
            .in3(N__19292),
            .lcout(\ADC_VAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC.n19413 ),
            .carryout(\ADC_VAC.n19414 ),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.bit_cnt_i7_LC_2_7_7 .C_ON=1'b0;
    defparam \ADC_VAC.bit_cnt_i7_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i7_LC_2_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i7_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__19421),
            .in2(_gnd_net_),
            .in3(N__19289),
            .lcout(\ADC_VAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57920),
            .ce(N__19499),
            .sr(N__19322));
    defparam \ADC_VAC.i6_4_lut_LC_2_8_1 .C_ON=1'b0;
    defparam \ADC_VAC.i6_4_lut_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i6_4_lut_LC_2_8_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \ADC_VAC.i6_4_lut_LC_2_8_1  (
            .in0(N__35008),
            .in1(N__19285),
            .in2(N__19274),
            .in3(N__35139),
            .lcout(\ADC_VAC.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19039_4_lut_LC_2_8_6 .C_ON=1'b0;
    defparam \ADC_VAC.i19039_4_lut_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19039_4_lut_LC_2_8_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ADC_VAC.i19039_4_lut_LC_2_8_6  (
            .in0(N__19258),
            .in1(N__19246),
            .in2(N__19235),
            .in3(N__19219),
            .lcout(),
            .ltout(\ADC_VAC.n21054_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i18824_4_lut_LC_2_8_7 .C_ON=1'b0;
    defparam \ADC_VAC.i18824_4_lut_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18824_4_lut_LC_2_8_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ADC_VAC.i18824_4_lut_LC_2_8_7  (
            .in0(N__19420),
            .in1(N__19409),
            .in2(N__19397),
            .in3(N__19394),
            .lcout(\ADC_VAC.n21053 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_3_6_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_3_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_3_6_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i0_LC_3_6_0  (
            .in0(N__19366),
            .in1(N__34296),
            .in2(N__19388),
            .in3(N__35215),
            .lcout(cmd_rdadctmp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57893),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_3_6_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_3_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_3_6_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i1_LC_3_6_5  (
            .in0(N__35214),
            .in1(N__19367),
            .in2(N__34333),
            .in3(N__19354),
            .lcout(cmd_rdadctmp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57893),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_3_7_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_3_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_3_7_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i4_LC_3_7_3  (
            .in0(N__35216),
            .in1(N__21826),
            .in2(N__34332),
            .in3(N__19333),
            .lcout(cmd_rdadctmp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57907),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_3_7_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_3_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_3_7_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i2_LC_3_7_4  (
            .in0(N__19342),
            .in1(N__34291),
            .in2(N__19358),
            .in3(N__35217),
            .lcout(cmd_rdadctmp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57907),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_3_7_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_3_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_3_7_6 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i3_LC_3_7_6  (
            .in0(N__19343),
            .in1(N__34292),
            .in2(N__19334),
            .in3(N__35218),
            .lcout(cmd_rdadctmp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57907),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i12409_2_lut_LC_3_7_7 .C_ON=1'b0;
    defparam \ADC_VAC.i12409_2_lut_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i12409_2_lut_LC_3_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ADC_VAC.i12409_2_lut_LC_3_7_7  (
            .in0(_gnd_net_),
            .in1(N__34938),
            .in2(_gnd_net_),
            .in3(N__19495),
            .lcout(\ADC_VAC.n14822 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i2_LC_3_8_0 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i2_LC_3_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i2_LC_3_8_0 .LUT_INIT=16'b0000111111000000;
    LogicCell40 \ADC_VAC.adc_state_i2_LC_3_8_0  (
            .in0(_gnd_net_),
            .in1(N__35166),
            .in2(N__34959),
            .in3(N__35024),
            .lcout(DTRIG_N_919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57921),
            .ce(N__19511),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i1_LC_3_8_1 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i1_LC_3_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i1_LC_3_8_1 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \ADC_VAC.adc_state_i1_LC_3_8_1  (
            .in0(N__35025),
            .in1(N__34949),
            .in2(_gnd_net_),
            .in3(N__35168),
            .lcout(adc_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57921),
            .ce(N__19511),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_LC_3_9_1 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_LC_3_9_1 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_VAC.i1_4_lut_LC_3_9_1  (
            .in0(N__34926),
            .in1(N__35130),
            .in2(N__19626),
            .in3(N__32228),
            .lcout(),
            .ltout(\ADC_VAC.n20715_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_adj_3_LC_3_9_2 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_adj_3_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_adj_3_LC_3_9_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \ADC_VAC.i1_2_lut_adj_3_LC_3_9_2  (
            .in0(N__35019),
            .in1(_gnd_net_),
            .in2(N__19529),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC.n20716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i0_LC_3_9_3 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i0_LC_3_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i0_LC_3_9_3 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \ADC_VAC.adc_state_i0_LC_3_9_3  (
            .in0(N__35165),
            .in1(N__35020),
            .in2(N__34945),
            .in3(N__19526),
            .lcout(adc_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57933),
            .ce(N__19520),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i30_4_lut_LC_3_9_5 .C_ON=1'b0;
    defparam \ADC_VAC.i30_4_lut_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i30_4_lut_LC_3_9_5 .LUT_INIT=16'b1100100001010001;
    LogicCell40 \ADC_VAC.i30_4_lut_LC_3_9_5  (
            .in0(N__34925),
            .in1(N__35018),
            .in2(N__19628),
            .in3(N__32227),
            .lcout(),
            .ltout(\ADC_VAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19134_2_lut_LC_3_9_6 .C_ON=1'b0;
    defparam \ADC_VAC.i19134_2_lut_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19134_2_lut_LC_3_9_6 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \ADC_VAC.i19134_2_lut_LC_3_9_6  (
            .in0(N__35129),
            .in1(_gnd_net_),
            .in2(N__19514),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_adj_4_LC_3_9_7 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_adj_4_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_adj_4_LC_3_9_7 .LUT_INIT=16'b0000000100100010;
    LogicCell40 \ADC_VAC.i1_4_lut_adj_4_LC_3_9_7  (
            .in0(N__34924),
            .in1(N__35128),
            .in2(N__19627),
            .in3(N__35017),
            .lcout(\ADC_VAC.n12489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.SCLK_35_LC_3_10_2 .C_ON=1'b0;
    defparam \ADC_VAC.SCLK_35_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.SCLK_35_LC_3_10_2 .LUT_INIT=16'b1011000011100010;
    LogicCell40 \ADC_VAC.SCLK_35_LC_3_10_2  (
            .in0(N__34941),
            .in1(N__35167),
            .in2(N__19468),
            .in3(N__35031),
            .lcout(VAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57944),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_140_LC_3_11_0.C_ON=1'b0;
    defparam i1_4_lut_adj_140_LC_3_11_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_140_LC_3_11_0.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_140_LC_3_11_0 (
            .in0(N__35170),
            .in1(N__34940),
            .in2(N__19438),
            .in3(N__35030),
            .lcout(),
            .ltout(n14_adj_1606_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.CS_37_LC_3_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.CS_37_LC_3_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.CS_37_LC_3_11_1 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \ADC_VAC.CS_37_LC_3_11_1  (
            .in0(N__19608),
            .in1(N__19634),
            .in2(N__19451),
            .in3(N__35171),
            .lcout(VAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57956),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_149_LC_3_11_4.C_ON=1'b0;
    defparam i1_2_lut_adj_149_LC_3_11_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_149_LC_3_11_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_149_LC_3_11_4 (
            .in0(_gnd_net_),
            .in1(N__34939),
            .in2(_gnd_net_),
            .in3(N__35029),
            .lcout(n20615),
            .ltout(n20615_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_3_lut_LC_3_11_5 .C_ON=1'b0;
    defparam \ADC_VAC.i1_3_lut_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_3_lut_LC_3_11_5 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \ADC_VAC.i1_3_lut_LC_3_11_5  (
            .in0(N__19609),
            .in1(_gnd_net_),
            .in2(N__19586),
            .in3(N__35169),
            .lcout(n12534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i2_LC_3_11_6 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i2_LC_3_11_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i2_LC_3_11_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \CLK_DDS.dds_state_i2_LC_3_11_6  (
            .in0(N__23393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23358),
            .lcout(dds_state_2_adj_1452),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57956),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_11_7 .C_ON=1'b0;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_11_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \CLK_DDS.i3_3_lut_4_lut_LC_3_11_7  (
            .in0(N__19581),
            .in1(N__23392),
            .in2(N__19567),
            .in3(N__22543),
            .lcout(n8_adj_1608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i3_LC_3_12_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i3_LC_3_12_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i3_LC_3_12_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \CLK_DDS.bit_cnt_i3_LC_3_12_0  (
            .in0(N__19583),
            .in1(N__19910),
            .in2(N__19928),
            .in3(N__19566),
            .lcout(bit_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57962),
            .ce(N__23357),
            .sr(N__19544));
    defparam \CLK_DDS.bit_cnt_i2_LC_3_12_1 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i2_LC_3_12_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i2_LC_3_12_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \CLK_DDS.bit_cnt_i2_LC_3_12_1  (
            .in0(N__19909),
            .in1(_gnd_net_),
            .in2(N__19568),
            .in3(N__19582),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57962),
            .ce(N__23357),
            .sr(N__19544));
    defparam \CLK_DDS.bit_cnt_i1_LC_3_12_2 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i1_LC_3_12_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i1_LC_3_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.bit_cnt_i1_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(N__19562),
            .in2(_gnd_net_),
            .in3(N__19908),
            .lcout(bit_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57962),
            .ce(N__23357),
            .sr(N__19544));
    defparam \CLK_DDS.i1_3_lut_LC_3_13_3 .C_ON=1'b0;
    defparam \CLK_DDS.i1_3_lut_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i1_3_lut_LC_3_13_3 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \CLK_DDS.i1_3_lut_LC_3_13_3  (
            .in0(N__23352),
            .in1(N__23421),
            .in2(_gnd_net_),
            .in3(N__22583),
            .lcout(\CLK_DDS.n16766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.avg_cnt_i0_LC_5_5_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i0_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i0_LC_5_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i0_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__19720),
            .in2(_gnd_net_),
            .in3(N__19532),
            .lcout(\ADC_VDC.avg_cnt_0 ),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\ADC_VDC.n19457 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i1_LC_5_5_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i1_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i1_LC_5_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i1_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__23815),
            .in2(_gnd_net_),
            .in3(N__19661),
            .lcout(\ADC_VDC.avg_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19457 ),
            .carryout(\ADC_VDC.n19458 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i2_LC_5_5_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i2_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i2_LC_5_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i2_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__23836),
            .in2(_gnd_net_),
            .in3(N__19658),
            .lcout(\ADC_VDC.avg_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19458 ),
            .carryout(\ADC_VDC.n19459 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i3_LC_5_5_3 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i3_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i3_LC_5_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i3_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__19765),
            .in2(_gnd_net_),
            .in3(N__19655),
            .lcout(\ADC_VDC.avg_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19459 ),
            .carryout(\ADC_VDC.n19460 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i4_LC_5_5_4 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i4_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i4_LC_5_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i4_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__19798),
            .in2(_gnd_net_),
            .in3(N__19652),
            .lcout(\ADC_VDC.avg_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19460 ),
            .carryout(\ADC_VDC.n19461 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i5_LC_5_5_5 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i5_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i5_LC_5_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i5_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__19750),
            .in2(_gnd_net_),
            .in3(N__19649),
            .lcout(\ADC_VDC.avg_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19461 ),
            .carryout(\ADC_VDC.n19462 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i6_LC_5_5_6 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i6_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i6_LC_5_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i6_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__23797),
            .in2(_gnd_net_),
            .in3(N__19646),
            .lcout(\ADC_VDC.avg_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19462 ),
            .carryout(\ADC_VDC.n19463 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i7_LC_5_5_7 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i7_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i7_LC_5_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i7_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__19783),
            .in2(_gnd_net_),
            .in3(N__19643),
            .lcout(\ADC_VDC.avg_cnt_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19463 ),
            .carryout(\ADC_VDC.n19464 ),
            .clk(N__40135),
            .ce(N__27171),
            .sr(N__27100));
    defparam \ADC_VDC.avg_cnt_i8_LC_5_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i8_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i8_LC_5_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i8_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__19702),
            .in2(_gnd_net_),
            .in3(N__19640),
            .lcout(\ADC_VDC.avg_cnt_8 ),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\ADC_VDC.n19465 ),
            .clk(N__40110),
            .ce(N__27173),
            .sr(N__27095));
    defparam \ADC_VDC.avg_cnt_i9_LC_5_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i9_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i9_LC_5_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i9_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__19735),
            .in2(_gnd_net_),
            .in3(N__19637),
            .lcout(\ADC_VDC.avg_cnt_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19465 ),
            .carryout(\ADC_VDC.n19466 ),
            .clk(N__40110),
            .ce(N__27173),
            .sr(N__27095));
    defparam \ADC_VDC.avg_cnt_i10_LC_5_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i10_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i10_LC_5_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i10_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__19687),
            .in2(_gnd_net_),
            .in3(N__19805),
            .lcout(\ADC_VDC.avg_cnt_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19466 ),
            .carryout(\ADC_VDC.n19467 ),
            .clk(N__40110),
            .ce(N__27173),
            .sr(N__27095));
    defparam \ADC_VDC.avg_cnt_i11_LC_5_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.avg_cnt_i11_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i11_LC_5_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i11_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__23854),
            .in2(_gnd_net_),
            .in3(N__19802),
            .lcout(\ADC_VDC.avg_cnt_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40110),
            .ce(N__27173),
            .sr(N__27095));
    defparam \ADC_VDC.i4_4_lut_adj_31_LC_5_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_31_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_31_LC_5_7_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_31_LC_5_7_0  (
            .in0(N__20971),
            .in1(N__20308),
            .in2(N__21071),
            .in3(N__20170),
            .lcout(\ADC_VDC.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_28_LC_5_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_28_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_28_LC_5_7_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_28_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__20258),
            .in2(_gnd_net_),
            .in3(N__20309),
            .lcout(\ADC_VDC.n6_adj_1410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i8_4_lut_LC_5_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.i8_4_lut_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i8_4_lut_LC_5_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i8_4_lut_LC_5_7_3  (
            .in0(N__19799),
            .in1(N__19784),
            .in2(N__19769),
            .in3(N__19751),
            .lcout(\ADC_VDC.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i1_LC_5_7_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i1_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i1_LC_5_7_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i1_LC_5_7_5  (
            .in0(N__23319),
            .in1(N__23511),
            .in2(N__19940),
            .in3(N__38398),
            .lcout(\CLK_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57879),
            .ce(N__23177),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7_4_lut_LC_5_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.i7_4_lut_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7_4_lut_LC_5_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i7_4_lut_LC_5_8_2  (
            .in0(N__19736),
            .in1(N__19721),
            .in2(N__19706),
            .in3(N__19688),
            .lcout(),
            .ltout(\ADC_VDC.n19_adj_1412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i11_3_lut_LC_5_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.i11_3_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i11_3_lut_LC_5_8_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ADC_VDC.i11_3_lut_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__19673),
            .in2(N__19667),
            .in3(N__23783),
            .lcout(\ADC_VDC.n18479 ),
            .ltout(\ADC_VDC.n18479_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16053_3_lut_LC_5_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.i16053_3_lut_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16053_3_lut_LC_5_8_4 .LUT_INIT=16'b0011001111111100;
    LogicCell40 \ADC_VDC.i16053_3_lut_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__32859),
            .in2(N__19664),
            .in3(N__33517),
            .lcout(\ADC_VDC.n18482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i19_LC_5_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i19_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i19_LC_5_8_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i19_LC_5_8_6  (
            .in0(N__29171),
            .in1(N__33372),
            .in2(N__23875),
            .in3(N__26861),
            .lcout(buf_adcdata_vdc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40132),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.CS_28_LC_5_9_4 .C_ON=1'b0;
    defparam \CLK_DDS.CS_28_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.CS_28_LC_5_9_4 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \CLK_DDS.CS_28_LC_5_9_4  (
            .in0(N__23316),
            .in1(N__23488),
            .in2(_gnd_net_),
            .in3(N__22573),
            .lcout(DDS_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57908),
            .ce(N__21755),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i11_LC_5_10_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i11_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i11_LC_5_10_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i11_LC_5_10_0  (
            .in0(N__23977),
            .in1(N__21545),
            .in2(N__21115),
            .in3(N__22156),
            .lcout(read_buf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i10_LC_5_10_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i10_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i10_LC_5_10_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.read_buf_i10_LC_5_10_1  (
            .in0(N__22155),
            .in1(N__20431),
            .in2(N__21560),
            .in3(N__23976),
            .lcout(read_buf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.mode_53_LC_5_10_2 .C_ON=1'b0;
    defparam \RTD.mode_53_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.mode_53_LC_5_10_2 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \RTD.mode_53_LC_5_10_2  (
            .in0(N__20321),
            .in1(N__21338),
            .in2(N__24102),
            .in3(N__22397),
            .lcout(\RTD.mode ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i12_LC_5_10_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i12_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i12_LC_5_10_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.read_buf_i12_LC_5_10_3  (
            .in0(N__22157),
            .in1(N__21111),
            .in2(N__21561),
            .in3(N__20196),
            .lcout(read_buf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i0_LC_5_10_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i0_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i0_LC_5_10_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.read_buf_i0_LC_5_10_4  (
            .in0(N__24885),
            .in1(N__19820),
            .in2(N__21559),
            .in3(N__22154),
            .lcout(read_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i14_LC_5_10_5 .C_ON=1'b0;
    defparam \RTD.read_buf_i14_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i14_LC_5_10_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i14_LC_5_10_5  (
            .in0(N__22159),
            .in1(N__23925),
            .in2(N__21563),
            .in3(N__20524),
            .lcout(read_buf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i15_LC_5_10_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i15_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i15_LC_5_10_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i15_LC_5_10_6  (
            .in0(N__23926),
            .in1(N__21546),
            .in2(N__21304),
            .in3(N__22160),
            .lcout(read_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i13_LC_5_10_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i13_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i13_LC_5_10_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i13_LC_5_10_7  (
            .in0(N__22158),
            .in1(N__20523),
            .in2(N__21562),
            .in3(N__20197),
            .lcout(read_buf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43760),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i0_LC_5_11_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i0_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i0_LC_5_11_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i0_LC_5_11_1  (
            .in0(N__23318),
            .in1(N__23440),
            .in2(N__23537),
            .in3(N__27539),
            .lcout(\CLK_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57934),
            .ce(N__23170),
            .sr(_gnd_net_));
    defparam i18807_2_lut_LC_5_12_0.C_ON=1'b0;
    defparam i18807_2_lut_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam i18807_2_lut_LC_5_12_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 i18807_2_lut_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(N__19899),
            .in2(_gnd_net_),
            .in3(N__19927),
            .lcout(n21227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i0_LC_5_12_3 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i0_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i0_LC_5_12_3 .LUT_INIT=16'b0001101000001010;
    LogicCell40 \CLK_DDS.bit_cnt_i0_LC_5_12_3  (
            .in0(N__19900),
            .in1(N__23484),
            .in2(N__23353),
            .in3(N__22580),
            .lcout(bit_cnt_0_adj_1456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57945),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_5_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_5_13_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i6_LC_5_13_0  (
            .in0(N__20459),
            .in1(N__52757),
            .in2(N__19853),
            .in3(N__51983),
            .lcout(cmd_rdadctmp_6_adj_1444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57957),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i30_4_lut_LC_5_13_3 .C_ON=1'b0;
    defparam \ADC_IAC.i30_4_lut_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i30_4_lut_LC_5_13_3 .LUT_INIT=16'b1100100001010001;
    LogicCell40 \ADC_IAC.i30_4_lut_LC_5_13_3  (
            .in0(N__35856),
            .in1(N__35789),
            .in2(N__20675),
            .in3(N__32213),
            .lcout(),
            .ltout(\ADC_IAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19132_2_lut_LC_5_13_4 .C_ON=1'b0;
    defparam \ADC_IAC.i19132_2_lut_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19132_2_lut_LC_5_13_4 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \ADC_IAC.i19132_2_lut_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19886),
            .in3(N__52756),
            .lcout(\ADC_IAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.SCLK_27_LC_5_13_5 .C_ON=1'b0;
    defparam \CLK_DDS.SCLK_27_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.SCLK_27_LC_5_13_5 .LUT_INIT=16'b0111001000110001;
    LogicCell40 \CLK_DDS.SCLK_27_LC_5_13_5  (
            .in0(N__23317),
            .in1(N__23483),
            .in2(N__19870),
            .in3(N__22582),
            .lcout(DDS_SCK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57957),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_5_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_5_13_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i7_LC_5_13_6  (
            .in0(N__19852),
            .in1(N__52758),
            .in2(N__25159),
            .in3(N__51984),
            .lcout(cmd_rdadctmp_7_adj_1443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57957),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_adj_5_LC_5_14_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_adj_5_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_adj_5_LC_5_14_0 .LUT_INIT=16'b0000000000110100;
    LogicCell40 \ADC_IAC.i1_4_lut_adj_5_LC_5_14_0  (
            .in0(N__20670),
            .in1(N__35787),
            .in2(N__35867),
            .in3(N__52707),
            .lcout(\ADC_IAC.n12586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i2_LC_5_14_1 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i2_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i2_LC_5_14_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_IAC.adc_state_i2_LC_5_14_1  (
            .in0(N__52708),
            .in1(N__35855),
            .in2(_gnd_net_),
            .in3(N__35786),
            .lcout(DTRIG_N_919_adj_1451),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57963),
            .ce(N__19970),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i1_LC_5_14_2 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i1_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i1_LC_5_14_2 .LUT_INIT=16'b0011000000110011;
    LogicCell40 \ADC_IAC.adc_state_i1_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__35788),
            .in2(N__35868),
            .in3(N__52709),
            .lcout(adc_state_1_adj_1417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57963),
            .ce(N__19970),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_199_LC_5_14_3.C_ON=1'b0;
    defparam i1_2_lut_adj_199_LC_5_14_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_199_LC_5_14_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_199_LC_5_14_3 (
            .in0(_gnd_net_),
            .in1(N__35847),
            .in2(_gnd_net_),
            .in3(N__35784),
            .lcout(n20612),
            .ltout(n20612_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_3_lut_LC_5_14_4 .C_ON=1'b0;
    defparam \ADC_IAC.i1_3_lut_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_3_lut_LC_5_14_4 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \ADC_IAC.i1_3_lut_LC_5_14_4  (
            .in0(N__20669),
            .in1(_gnd_net_),
            .in2(N__19955),
            .in3(N__52706),
            .lcout(n12663),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_5_14_7.C_ON=1'b0;
    defparam i1_2_lut_LC_5_14_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_5_14_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_LC_5_14_7 (
            .in0(_gnd_net_),
            .in1(N__35851),
            .in2(_gnd_net_),
            .in3(N__35785),
            .lcout(n20584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_2_lut_LC_5_15_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_2_lut_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_2_lut_LC_5_15_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \ADC_IAC.i1_2_lut_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__35790),
            .in2(_gnd_net_),
            .in3(N__19952),
            .lcout(\ADC_IAC.n20714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_LC_5_15_1 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_LC_5_15_1 .LUT_INIT=16'b1010101111101111;
    LogicCell40 \ADC_IAC.i1_4_lut_LC_5_15_1  (
            .in0(N__52720),
            .in1(N__35857),
            .in2(N__20657),
            .in3(N__32226),
            .lcout(\ADC_IAC.n20713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i18169_4_lut_LC_5_15_2 .C_ON=1'b0;
    defparam \ADC_IAC.i18169_4_lut_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i18169_4_lut_LC_5_15_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_IAC.i18169_4_lut_LC_5_15_2  (
            .in0(N__20866),
            .in1(N__20545),
            .in2(N__20579),
            .in3(N__20560),
            .lcout(),
            .ltout(\ADC_IAC.n20783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i18181_4_lut_LC_5_15_3 .C_ON=1'b0;
    defparam \ADC_IAC.i18181_4_lut_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i18181_4_lut_LC_5_15_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_IAC.i18181_4_lut_LC_5_15_3  (
            .in0(N__20836),
            .in1(N__20593),
            .in2(N__19946),
            .in3(N__20818),
            .lcout(),
            .ltout(\ADC_IAC.n20795_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i18845_4_lut_LC_5_15_4 .C_ON=1'b0;
    defparam \ADC_IAC.i18845_4_lut_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i18845_4_lut_LC_5_15_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_IAC.i18845_4_lut_LC_5_15_4  (
            .in0(N__20851),
            .in1(N__52721),
            .in2(N__19943),
            .in3(N__35791),
            .lcout(),
            .ltout(\ADC_IAC.n21068_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i0_LC_5_15_5 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i0_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i0_LC_5_15_5 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \ADC_IAC.adc_state_i0_LC_5_15_5  (
            .in0(N__35792),
            .in1(N__52755),
            .in2(N__20063),
            .in3(N__35858),
            .lcout(adc_state_0_adj_1418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57971),
            .ce(N__20060),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_5_16_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_5_16_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i1_LC_5_16_0  (
            .in0(N__52754),
            .in1(N__20030),
            .in2(N__20774),
            .in3(N__52015),
            .lcout(cmd_rdadctmp_1_adj_1449),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57975),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_5_16_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_5_16_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i0_LC_5_16_2  (
            .in0(N__52753),
            .in1(N__20029),
            .in2(N__20051),
            .in3(N__52014),
            .lcout(cmd_rdadctmp_0_adj_1450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57975),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.SCLK_35_LC_5_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.SCLK_35_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.SCLK_35_LC_5_16_4 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_IAC.SCLK_35_LC_5_16_4  (
            .in0(N__52752),
            .in1(N__35869),
            .in2(N__20011),
            .in3(N__35803),
            .lcout(IAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57975),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i1_LC_5_17_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i1_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i1_LC_5_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.dds_state_i1_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__23510),
            .in2(_gnd_net_),
            .in3(N__22581),
            .lcout(dds_state_1_adj_1453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57979),
            .ce(N__22492),
            .sr(N__23359));
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_6_4_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_6_4_1 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i29_LC_6_4_1  (
            .in0(N__35320),
            .in1(N__21909),
            .in2(N__19993),
            .in3(N__34335),
            .lcout(cmd_rdadctmp_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57830),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_6_4_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_6_4_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i28_LC_6_4_5  (
            .in0(N__35319),
            .in1(N__29459),
            .in2(N__19992),
            .in3(N__34334),
            .lcout(cmd_rdadctmp_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57830),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i20_LC_6_5_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i20_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i20_LC_6_5_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i20_LC_6_5_0  (
            .in0(N__34653),
            .in1(N__35306),
            .in2(N__19994),
            .in3(N__21942),
            .lcout(buf_adcdata_vac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57840),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16066_3_lut_LC_6_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i16066_3_lut_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16066_3_lut_LC_6_5_4 .LUT_INIT=16'b1101110110101010;
    LogicCell40 \ADC_VDC.i16066_3_lut_LC_6_5_4  (
            .in0(N__33612),
            .in1(N__32872),
            .in2(_gnd_net_),
            .in3(N__33519),
            .lcout(\ADC_VDC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18135_2_lut_LC_6_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i18135_2_lut_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18135_2_lut_LC_6_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VDC.i18135_2_lut_LC_6_5_5  (
            .in0(N__32871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33613),
            .lcout(\ADC_VDC.n20748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i15177_2_lut_LC_6_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i15177_2_lut_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i15177_2_lut_LC_6_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i15177_2_lut_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__32870),
            .in2(_gnd_net_),
            .in3(N__33518),
            .lcout(\ADC_VDC.n7_adj_1411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.bit_cnt_3780__i0_LC_6_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i0_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i0_LC_6_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i0_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__20975),
            .in2(_gnd_net_),
            .in3(N__20087),
            .lcout(\ADC_VDC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\ADC_VDC.n19531 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i1_LC_6_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i1_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i1_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i1_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__21070),
            .in2(_gnd_net_),
            .in3(N__20084),
            .lcout(\ADC_VDC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19531 ),
            .carryout(\ADC_VDC.n19532 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i2_LC_6_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i2_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i2_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i2_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__20314),
            .in2(_gnd_net_),
            .in3(N__20081),
            .lcout(\ADC_VDC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19532 ),
            .carryout(\ADC_VDC.n19533 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i3_LC_6_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i3_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i3_LC_6_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i3_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__20267),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\ADC_VDC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19533 ),
            .carryout(\ADC_VDC.n19534 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i4_LC_6_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i4_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i4_LC_6_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i4_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__21020),
            .in2(_gnd_net_),
            .in3(N__20075),
            .lcout(\ADC_VDC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19534 ),
            .carryout(\ADC_VDC.n19535 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i5_LC_6_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i5_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i5_LC_6_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i5_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__20171),
            .in2(_gnd_net_),
            .in3(N__20072),
            .lcout(\ADC_VDC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19535 ),
            .carryout(\ADC_VDC.n19536 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i6_LC_6_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3780__i6_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i6_LC_6_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i6_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__20129),
            .in2(_gnd_net_),
            .in3(N__20069),
            .lcout(\ADC_VDC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19536 ),
            .carryout(\ADC_VDC.n19537 ),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.bit_cnt_3780__i7_LC_6_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.bit_cnt_3780__i7_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3780__i7_LC_6_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3780__i7_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__20144),
            .in2(_gnd_net_),
            .in3(N__20066),
            .lcout(\ADC_VDC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40109),
            .ce(N__33647),
            .sr(N__21134));
    defparam \ADC_VDC.i18857_4_lut_LC_6_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.i18857_4_lut_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18857_4_lut_LC_6_7_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \ADC_VDC.i18857_4_lut_LC_6_7_0  (
            .in0(N__20114),
            .in1(N__33521),
            .in2(N__21027),
            .in3(N__21041),
            .lcout(\ADC_VDC.n21079 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_3_lut_LC_6_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.i2_3_lut_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_3_lut_LC_6_7_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i2_3_lut_LC_6_7_1  (
            .in0(N__20169),
            .in1(N__20142),
            .in2(_gnd_net_),
            .in3(N__20127),
            .lcout(\ADC_VDC.n20534 ),
            .ltout(\ADC_VDC.n20534_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_6_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_6_7_2 .LUT_INIT=16'b1111111011111110;
    LogicCell40 \ADC_VDC.i1_2_lut_3_lut_LC_6_7_2  (
            .in0(N__20972),
            .in1(N__21067),
            .in2(N__20153),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i5_3_lut_LC_6_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.i5_3_lut_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i5_3_lut_LC_6_7_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \ADC_VDC.i5_3_lut_LC_6_7_3  (
            .in0(N__20150),
            .in1(N__20143),
            .in2(_gnd_net_),
            .in3(N__20128),
            .lcout(\ADC_VDC.n20562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i8_LC_6_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i8_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i8_LC_6_7_5 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.ADC_DATA_i8_LC_6_7_5  (
            .in0(N__26621),
            .in1(N__30535),
            .in2(N__29177),
            .in3(N__33346),
            .lcout(buf_adcdata_vdc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40120),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i23_LC_6_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i23_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i23_LC_6_7_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i23_LC_6_7_6  (
            .in0(N__33345),
            .in1(N__29173),
            .in2(N__22294),
            .in3(N__27029),
            .lcout(buf_adcdata_vdc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40120),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19094_4_lut_LC_6_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.i19094_4_lut_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19094_4_lut_LC_6_7_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ADC_VDC.i19094_4_lut_LC_6_7_7  (
            .in0(N__21068),
            .in1(N__20973),
            .in2(N__20268),
            .in3(N__20310),
            .lcout(\ADC_VDC.n21082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.n21974_bdd_4_lut_4_lut_LC_6_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.n21974_bdd_4_lut_4_lut_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.n21974_bdd_4_lut_4_lut_LC_6_8_0 .LUT_INIT=16'b1101110100110000;
    LogicCell40 \ADC_VDC.n21974_bdd_4_lut_4_lut_LC_6_8_0  (
            .in0(N__33516),
            .in1(N__33349),
            .in2(N__20108),
            .in3(N__20276),
            .lcout(),
            .ltout(\ADC_VDC.n21977_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i1_LC_6_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i1_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i1_LC_6_8_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.adc_state_i1_LC_6_8_1  (
            .in0(N__33350),
            .in1(N__33022),
            .in2(N__20096),
            .in3(N__20093),
            .lcout(\ADC_VDC.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40111),
            .ce(N__20213),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_LC_6_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_LC_6_8_2 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \ADC_VDC.i4_4_lut_LC_6_8_2  (
            .in0(N__20269),
            .in1(N__20315),
            .in2(N__21028),
            .in3(N__20285),
            .lcout(\ADC_VDC.n10552 ),
            .ltout(\ADC_VDC.n10552_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_6_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_6_8_3 .LUT_INIT=16'b0110011001001100;
    LogicCell40 \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_6_8_3  (
            .in0(N__33348),
            .in1(N__32858),
            .in2(N__20279),
            .in3(N__33515),
            .lcout(\ADC_VDC.n21974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18952_4_lut_LC_6_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.i18952_4_lut_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18952_4_lut_LC_6_8_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \ADC_VDC.i18952_4_lut_LC_6_8_4  (
            .in0(N__20270),
            .in1(N__33011),
            .in2(N__21029),
            .in3(N__20237),
            .lcout(),
            .ltout(\ADC_VDC.n21224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i37_4_lut_LC_6_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.i37_4_lut_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i37_4_lut_LC_6_8_5 .LUT_INIT=16'b1101000110101010;
    LogicCell40 \ADC_VDC.i37_4_lut_LC_6_8_5  (
            .in0(N__33588),
            .in1(N__32857),
            .in2(N__20228),
            .in3(N__33514),
            .lcout(),
            .ltout(\ADC_VDC.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_LC_6_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_LC_6_8_6 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \ADC_VDC.i1_4_lut_LC_6_8_6  (
            .in0(N__20225),
            .in1(N__33012),
            .in2(N__20216),
            .in3(N__33347),
            .lcout(\ADC_VDC.n20555 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i6_LC_6_9_1 .C_ON=1'b0;
    defparam \RTD.adress_i6_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i6_LC_6_9_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \RTD.adress_i6_LC_6_9_1  (
            .in0(N__21283),
            .in1(N__20490),
            .in2(N__20360),
            .in3(N__21211),
            .lcout(adress_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43813),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i12_LC_6_9_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i12_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i12_LC_6_9_2 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i12_LC_6_9_2  (
            .in0(N__25408),
            .in1(N__24201),
            .in2(N__20201),
            .in3(N__24473),
            .lcout(buf_readRTD_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43813),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i4_LC_6_9_3 .C_ON=1'b0;
    defparam \RTD.adress_i4_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i4_LC_6_9_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \RTD.adress_i4_LC_6_9_3  (
            .in0(N__20368),
            .in1(N__20486),
            .in2(N__20183),
            .in3(N__21209),
            .lcout(adress_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43813),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i3_LC_6_9_4 .C_ON=1'b0;
    defparam \RTD.adress_i3_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i3_LC_6_9_4 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \RTD.adress_i3_LC_6_9_4  (
            .in0(N__21208),
            .in1(N__20378),
            .in2(N__20491),
            .in3(N__20179),
            .lcout(adress_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43813),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i2_LC_6_9_5 .C_ON=1'b0;
    defparam \RTD.adress_i2_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i2_LC_6_9_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \RTD.adress_i2_LC_6_9_5  (
            .in0(N__20377),
            .in1(N__20482),
            .in2(N__20414),
            .in3(N__21207),
            .lcout(adress_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43813),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i5_LC_6_9_6 .C_ON=1'b0;
    defparam \RTD.adress_i5_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i5_LC_6_9_6 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \RTD.adress_i5_LC_6_9_6  (
            .in0(N__21210),
            .in1(N__20369),
            .in2(N__20492),
            .in3(N__20356),
            .lcout(adress_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43813),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.MOSI_59_LC_6_10_0 .C_ON=1'b0;
    defparam \RTD.MOSI_59_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.MOSI_59_LC_6_10_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \RTD.MOSI_59_LC_6_10_0  (
            .in0(N__24447),
            .in1(N__21238),
            .in2(N__21398),
            .in3(N__24847),
            .lcout(RTD_SDI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43815),
            .ce(N__21347),
            .sr(N__24514));
    defparam \RTD.i18150_rep_64_2_lut_LC_6_10_1 .C_ON=1'b0;
    defparam \RTD.i18150_rep_64_2_lut_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i18150_rep_64_2_lut_LC_6_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i18150_rep_64_2_lut_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__24443),
            .in2(_gnd_net_),
            .in3(N__24843),
            .lcout(\RTD.n22370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19089_3_lut_LC_6_10_2 .C_ON=1'b0;
    defparam \RTD.i19089_3_lut_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i19089_3_lut_LC_6_10_2 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \RTD.i19089_3_lut_LC_6_10_2  (
            .in0(N__22425),
            .in1(N__24845),
            .in2(_gnd_net_),
            .in3(N__21333),
            .lcout(),
            .ltout(\RTD.n21309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_7_LC_6_10_3 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_7_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_7_LC_6_10_3 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \RTD.i1_4_lut_adj_7_LC_6_10_3  (
            .in0(N__24673),
            .in1(N__24445),
            .in2(N__20324),
            .in3(N__22454),
            .lcout(\RTD.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i16303_3_lut_LC_6_10_4 .C_ON=1'b0;
    defparam \RTD.i16303_3_lut_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i16303_3_lut_LC_6_10_4 .LUT_INIT=16'b1111101001010101;
    LogicCell40 \RTD.i16303_3_lut_LC_6_10_4  (
            .in0(N__24444),
            .in1(_gnd_net_),
            .in2(N__22461),
            .in3(N__24844),
            .lcout(\RTD.n20762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_11_LC_6_10_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_11_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_11_LC_6_10_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \RTD.i1_2_lut_adj_11_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__24842),
            .in2(_gnd_net_),
            .in3(N__24664),
            .lcout(\RTD.n20631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i34_4_lut_4_lut_LC_6_10_6 .C_ON=1'b0;
    defparam \RTD.i34_4_lut_4_lut_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i34_4_lut_4_lut_LC_6_10_6 .LUT_INIT=16'b1100111111000111;
    LogicCell40 \RTD.i34_4_lut_4_lut_LC_6_10_6  (
            .in0(N__22426),
            .in1(N__24846),
            .in2(N__25049),
            .in3(N__22387),
            .lcout(),
            .ltout(\RTD.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i36_4_lut_4_lut_LC_6_10_7 .C_ON=1'b0;
    defparam \RTD.i36_4_lut_4_lut_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i36_4_lut_4_lut_LC_6_10_7 .LUT_INIT=16'b1000100000110000;
    LogicCell40 \RTD.i36_4_lut_4_lut_LC_6_10_7  (
            .in0(N__22637),
            .in1(N__24446),
            .in2(N__20435),
            .in3(N__24665),
            .lcout(n13181),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i9_LC_6_11_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i9_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i9_LC_6_11_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i9_LC_6_11_0  (
            .in0(N__20510),
            .in1(N__21524),
            .in2(N__20432),
            .in3(N__22163),
            .lcout(read_buf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i9_LC_6_11_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i9_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i9_LC_6_11_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \RTD.READ_DATA_i9_LC_6_11_1  (
            .in0(N__24470),
            .in1(N__20430),
            .in2(N__24235),
            .in3(N__27562),
            .lcout(buf_readRTD_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i1_LC_6_11_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i1_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i1_LC_6_11_2 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i1_LC_6_11_2  (
            .in0(N__43339),
            .in1(N__24222),
            .in2(N__20396),
            .in3(N__24472),
            .lcout(buf_readRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i2_LC_6_11_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i2_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i2_LC_6_11_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.read_buf_i2_LC_6_11_3  (
            .in0(N__22162),
            .in1(N__20394),
            .in2(N__21607),
            .in3(N__21525),
            .lcout(read_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i3_LC_6_11_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i3_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i3_LC_6_11_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \RTD.READ_DATA_i3_LC_6_11_4  (
            .in0(N__38311),
            .in1(N__24471),
            .in2(N__21587),
            .in3(N__24223),
            .lcout(buf_readRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i1_LC_6_11_5 .C_ON=1'b0;
    defparam \RTD.adress_i1_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i1_LC_6_11_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.adress_i1_LC_6_11_5  (
            .in0(N__20470),
            .in1(N__20407),
            .in2(N__21227),
            .in3(N__21206),
            .lcout(adress_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i1_LC_6_11_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i1_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i1_LC_6_11_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i1_LC_6_11_6  (
            .in0(N__24893),
            .in1(N__21523),
            .in2(N__20395),
            .in3(N__22161),
            .lcout(read_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43805),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12602_2_lut_LC_6_11_7 .C_ON=1'b0;
    defparam \RTD.i12602_2_lut_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i12602_2_lut_LC_6_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RTD.i12602_2_lut_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(N__24676),
            .in2(_gnd_net_),
            .in3(N__21376),
            .lcout(\RTD.n15015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i8_LC_6_12_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i8_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i8_LC_6_12_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \RTD.READ_DATA_i8_LC_6_12_1  (
            .in0(N__24468),
            .in1(N__25375),
            .in2(N__24236),
            .in3(N__20506),
            .lcout(buf_readRTD_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43761),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i7_LC_6_12_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i7_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i7_LC_6_12_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.read_buf_i7_LC_6_12_2  (
            .in0(N__21521),
            .in1(N__21621),
            .in2(N__24259),
            .in3(N__22168),
            .lcout(read_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43761),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i13_LC_6_12_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i13_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i13_LC_6_12_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i13_LC_6_12_4  (
            .in0(N__25132),
            .in1(N__24229),
            .in2(N__20531),
            .in3(N__24469),
            .lcout(buf_readRTD_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43761),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i8_LC_6_12_5 .C_ON=1'b0;
    defparam \RTD.read_buf_i8_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i8_LC_6_12_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i8_LC_6_12_5  (
            .in0(N__22169),
            .in1(N__20505),
            .in2(N__21628),
            .in3(N__21522),
            .lcout(read_buf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43761),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i6_LC_6_12_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i6_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i6_LC_6_12_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i6_LC_6_12_6  (
            .in0(N__21520),
            .in1(N__21464),
            .in2(N__24258),
            .in3(N__22167),
            .lcout(read_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43761),
            .ce(),
            .sr(_gnd_net_));
    defparam i18141_2_lut_LC_6_12_7.C_ON=1'b0;
    defparam i18141_2_lut_LC_6_12_7.SEQ_MODE=4'b0000;
    defparam i18141_2_lut_LC_6_12_7.LUT_INIT=16'b1101110111011101;
    LogicCell40 i18141_2_lut_LC_6_12_7 (
            .in0(N__25040),
            .in1(N__24643),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n20754),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_6_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_6_13_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i30_LC_6_13_0  (
            .in0(N__51981),
            .in1(N__21735),
            .in2(N__52916),
            .in3(N__21444),
            .lcout(cmd_rdadctmp_30_adj_1420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57935),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_6_13_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_6_13_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i29_LC_6_13_5  (
            .in0(N__20706),
            .in1(N__52850),
            .in2(N__21448),
            .in3(N__51982),
            .lcout(cmd_rdadctmp_29_adj_1421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57935),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_6_14_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_6_14_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i28_LC_6_14_0  (
            .in0(N__52747),
            .in1(N__25297),
            .in2(N__20710),
            .in3(N__51979),
            .lcout(cmd_rdadctmp_28_adj_1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57946),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_6_14_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_6_14_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i5_LC_6_14_1  (
            .in0(N__51978),
            .in1(N__20458),
            .in2(N__20447),
            .in3(N__52751),
            .lcout(cmd_rdadctmp_5_adj_1445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57946),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_6_14_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_6_14_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i4_LC_6_14_2  (
            .in0(N__52748),
            .in1(N__20443),
            .in2(N__20687),
            .in3(N__51980),
            .lcout(cmd_rdadctmp_4_adj_1446),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57946),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i3_LC_6_14_3  (
            .in0(N__51977),
            .in1(N__20683),
            .in2(N__20759),
            .in3(N__52750),
            .lcout(cmd_rdadctmp_3_adj_1447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57946),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_137_LC_6_14_4.C_ON=1'b0;
    defparam i1_4_lut_adj_137_LC_6_14_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_137_LC_6_14_4.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_137_LC_6_14_4 (
            .in0(N__52746),
            .in1(N__35859),
            .in2(N__20611),
            .in3(N__35799),
            .lcout(),
            .ltout(n14_adj_1604_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.CS_37_LC_6_14_5 .C_ON=1'b0;
    defparam \ADC_IAC.CS_37_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.CS_37_LC_6_14_5 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \ADC_IAC.CS_37_LC_6_14_5  (
            .in0(N__20671),
            .in1(N__20630),
            .in2(N__20624),
            .in3(N__52749),
            .lcout(IAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57946),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i12447_2_lut_LC_6_14_6 .C_ON=1'b0;
    defparam \ADC_IAC.i12447_2_lut_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i12447_2_lut_LC_6_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ADC_IAC.i12447_2_lut_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__35860),
            .in2(_gnd_net_),
            .in3(N__20797),
            .lcout(\ADC_IAC.n14860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.bit_cnt_i0_LC_6_15_0 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i0_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i0_LC_6_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i0_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__20594),
            .in2(_gnd_net_),
            .in3(N__20582),
            .lcout(\ADC_IAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\ADC_IAC.n19415 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i1_LC_6_15_1 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i1_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i1_LC_6_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i1_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__20578),
            .in2(_gnd_net_),
            .in3(N__20564),
            .lcout(\ADC_IAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_IAC.n19415 ),
            .carryout(\ADC_IAC.n19416 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i2_LC_6_15_2 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i2_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i2_LC_6_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i2_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__20561),
            .in2(_gnd_net_),
            .in3(N__20549),
            .lcout(\ADC_IAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_IAC.n19416 ),
            .carryout(\ADC_IAC.n19417 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i3_LC_6_15_3 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i3_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i3_LC_6_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i3_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__20546),
            .in2(_gnd_net_),
            .in3(N__20534),
            .lcout(\ADC_IAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_IAC.n19417 ),
            .carryout(\ADC_IAC.n19418 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i4_LC_6_15_4 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i4_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i4_LC_6_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i4_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__20867),
            .in2(_gnd_net_),
            .in3(N__20855),
            .lcout(\ADC_IAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_IAC.n19418 ),
            .carryout(\ADC_IAC.n19419 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i5_LC_6_15_5 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i5_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i5_LC_6_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i5_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(N__20852),
            .in2(_gnd_net_),
            .in3(N__20840),
            .lcout(\ADC_IAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_IAC.n19419 ),
            .carryout(\ADC_IAC.n19420 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i6_LC_6_15_6 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i6_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i6_LC_6_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i6_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(N__20837),
            .in2(_gnd_net_),
            .in3(N__20825),
            .lcout(\ADC_IAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_IAC.n19420 ),
            .carryout(\ADC_IAC.n19421 ),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \ADC_IAC.bit_cnt_i7_LC_6_15_7 .C_ON=1'b0;
    defparam \ADC_IAC.bit_cnt_i7_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i7_LC_6_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i7_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(N__20819),
            .in2(_gnd_net_),
            .in3(N__20822),
            .lcout(\ADC_IAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57958),
            .ce(N__20807),
            .sr(N__20786));
    defparam \CLK_DDS.i19097_4_lut_LC_6_16_2 .C_ON=1'b0;
    defparam \CLK_DDS.i19097_4_lut_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19097_4_lut_LC_6_16_2 .LUT_INIT=16'b1000100111001100;
    LogicCell40 \CLK_DDS.i19097_4_lut_LC_6_16_2  (
            .in0(N__23228),
            .in1(N__23489),
            .in2(N__23126),
            .in3(N__22574),
            .lcout(\CLK_DDS.n12800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_6_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_6_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_6_17_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i2_LC_6_17_7  (
            .in0(N__20773),
            .in1(N__52819),
            .in2(N__20755),
            .in3(N__52016),
            .lcout(cmd_rdadctmp_2_adj_1448),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57972),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_main.i19670_1_lut_LC_7_1_7 .C_ON=1'b0;
    defparam \pll_main.i19670_1_lut_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \pll_main.i19670_1_lut_LC_7_1_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_main.i19670_1_lut_LC_7_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45097),
            .lcout(DDS_MCLK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i20_LC_7_3_2 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i20_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i20_LC_7_3_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i20_LC_7_3_2  (
            .in0(N__53184),
            .in1(N__52995),
            .in2(N__20720),
            .in3(N__40362),
            .lcout(buf_adcdata_iac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57817),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i2_LC_7_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i2_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i2_LC_7_4_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \ADC_VDC.adc_state_i2_LC_7_4_2  (
            .in0(N__33240),
            .in1(N__32896),
            .in2(_gnd_net_),
            .in3(N__33523),
            .lcout(adc_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40108),
            .ce(N__20915),
            .sr(N__20909));
    defparam \ADC_VDC.ADC_DATA_i2_LC_7_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i2_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i2_LC_7_5_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i2_LC_7_5_0  (
            .in0(N__29131),
            .in1(N__33239),
            .in2(N__28636),
            .in3(N__26315),
            .lcout(buf_adcdata_vdc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40134),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_7_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_7_5_1 .LUT_INIT=16'b1010110100100101;
    LogicCell40 \ADC_VDC.i40_3_lut_4_lut_LC_7_5_1  (
            .in0(N__33492),
            .in1(N__32898),
            .in2(N__33632),
            .in3(N__20947),
            .lcout(),
            .ltout(\ADC_VDC.n19_adj_1413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19163_4_lut_LC_7_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i19163_4_lut_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19163_4_lut_LC_7_5_2 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_VDC.i19163_4_lut_LC_7_5_2  (
            .in0(N__33044),
            .in1(N__33238),
            .in2(N__20918),
            .in3(N__20884),
            .lcout(\ADC_VDC.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19168_4_lut_LC_7_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i19168_4_lut_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19168_4_lut_LC_7_5_3 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \ADC_VDC.i19168_4_lut_LC_7_5_3  (
            .in0(N__20894),
            .in1(N__33235),
            .in2(N__33631),
            .in3(N__33043),
            .lcout(\ADC_VDC.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7717_3_lut_4_lut_LC_7_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i7717_3_lut_4_lut_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7717_3_lut_4_lut_LC_7_5_4 .LUT_INIT=16'b0101001111001100;
    LogicCell40 \ADC_VDC.i7717_3_lut_4_lut_LC_7_5_4  (
            .in0(N__20948),
            .in1(N__33628),
            .in2(N__32906),
            .in3(N__33493),
            .lcout(),
            .ltout(\ADC_VDC.n10132_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_7_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_7_5_5 .LUT_INIT=16'b1101110111111100;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_LC_7_5_5  (
            .in0(N__20885),
            .in1(N__33236),
            .in2(N__20897),
            .in3(N__33045),
            .lcout(\ADC_VDC.n12823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18137_2_lut_LC_7_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i18137_2_lut_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18137_2_lut_LC_7_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i18137_2_lut_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__33621),
            .in2(_gnd_net_),
            .in3(N__20893),
            .lcout(\ADC_VDC.n20750 ),
            .ltout(\ADC_VDC.n20750_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_32_LC_7_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_32_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_32_LC_7_5_7 .LUT_INIT=16'b1100111111101110;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_32_LC_7_5_7  (
            .in0(N__20876),
            .in1(N__33234),
            .in2(N__20870),
            .in3(N__33042),
            .lcout(\ADC_VDC.n72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19101_4_lut_4_lut_LC_7_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.i19101_4_lut_4_lut_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19101_4_lut_4_lut_LC_7_6_0 .LUT_INIT=16'b1111111011110001;
    LogicCell40 \ADC_VDC.i19101_4_lut_4_lut_LC_7_6_0  (
            .in0(N__33476),
            .in1(N__32904),
            .in2(N__33126),
            .in3(N__33283),
            .lcout(),
            .ltout(\ADC_VDC.n11692_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.SCLK_46_LC_7_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.SCLK_46_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.SCLK_46_LC_7_6_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.SCLK_46_LC_7_6_1  (
            .in0(N__32905),
            .in1(N__21088),
            .in2(N__21095),
            .in3(N__25820),
            .lcout(VDC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40060),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i1_LC_7_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i1_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i1_LC_7_6_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i1_LC_7_6_2  (
            .in0(N__29110),
            .in1(N__33285),
            .in2(N__28933),
            .in3(N__26348),
            .lcout(buf_adcdata_vdc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40060),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_LC_7_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_LC_7_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__21069),
            .in2(_gnd_net_),
            .in3(N__21040),
            .lcout(),
            .ltout(\ADC_VDC.n11281_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_adj_29_LC_7_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_29_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_29_LC_7_6_4 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_29_LC_7_6_4  (
            .in0(N__21016),
            .in1(N__20990),
            .in2(N__20978),
            .in3(N__20974),
            .lcout(\ADC_VDC.n15 ),
            .ltout(\ADC_VDC.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18133_2_lut_LC_7_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i18133_2_lut_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18133_2_lut_LC_7_6_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ADC_VDC.i18133_2_lut_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20939),
            .in3(N__33475),
            .lcout(),
            .ltout(\ADC_VDC.n20746_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_33_LC_7_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_33_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_33_LC_7_6_6 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_33_LC_7_6_6  (
            .in0(N__21146),
            .in1(N__32903),
            .in2(N__20936),
            .in3(N__20933),
            .lcout(\ADC_VDC.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i7_LC_7_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i7_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i7_LC_7_6_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i7_LC_7_6_7  (
            .in0(N__33284),
            .in1(N__29111),
            .in2(N__23671),
            .in3(N__26660),
            .lcout(buf_adcdata_vdc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40060),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i3_LC_7_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i3_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i3_LC_7_7_1 .LUT_INIT=16'b0010010000001100;
    LogicCell40 \ADC_VDC.adc_state_i3_LC_7_7_1  (
            .in0(N__33472),
            .in1(N__32988),
            .in2(N__33340),
            .in3(N__32860),
            .lcout(adc_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40133),
            .ce(N__20927),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_7_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_7_7_2 .LUT_INIT=16'b1110101000001000;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_7_7_2  (
            .in0(N__32983),
            .in1(N__32845),
            .in2(N__33520),
            .in3(N__33270),
            .lcout(\ADC_VDC.n13038 ),
            .ltout(\ADC_VDC.n13038_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i12557_2_lut_LC_7_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.i12557_2_lut_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i12557_2_lut_LC_7_7_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ADC_VDC.i12557_2_lut_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21149),
            .in3(N__32985),
            .lcout(\ADC_VDC.n14931 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_30_LC_7_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_30_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_30_LC_7_7_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_30_LC_7_7_4  (
            .in0(N__32984),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33271),
            .lcout(\ADC_VDC.n20659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_36_LC_7_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_36_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_36_LC_7_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_36_LC_7_7_5  (
            .in0(N__33273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32986),
            .lcout(\ADC_VDC.n20392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i15034_2_lut_LC_7_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.i15034_2_lut_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i15034_2_lut_LC_7_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i15034_2_lut_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__33272),
            .in2(_gnd_net_),
            .in3(N__32846),
            .lcout(),
            .ltout(\ADC_VDC.n17432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_35_LC_7_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_35_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_35_LC_7_7_7 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_adj_35_LC_7_7_7  (
            .in0(N__33471),
            .in1(N__32987),
            .in2(N__21137),
            .in3(N__32768),
            .lcout(\ADC_VDC.n18466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i1_LC_7_8_0 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i1_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i1_LC_7_8_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.cfg_buf_i1_LC_7_8_0  (
            .in0(N__24140),
            .in1(N__24107),
            .in2(N__27626),
            .in3(N__22316),
            .lcout(\RTD.cfg_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i5_LC_7_8_1 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i5_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i5_LC_7_8_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i5_LC_7_8_1  (
            .in0(N__24110),
            .in1(N__24143),
            .in2(N__27505),
            .in3(N__21182),
            .lcout(\RTD.cfg_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i3_LC_7_8_2 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i3_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i3_LC_7_8_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.cfg_buf_i3_LC_7_8_2  (
            .in0(N__24142),
            .in1(N__24109),
            .in2(N__21170),
            .in3(N__25205),
            .lcout(\RTD.cfg_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i0_LC_7_8_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i0_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i0_LC_7_8_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i0_LC_7_8_3  (
            .in0(N__24106),
            .in1(N__24139),
            .in2(N__25364),
            .in3(N__21260),
            .lcout(\RTD.cfg_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i11_LC_7_8_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i11_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i11_LC_7_8_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i11_LC_7_8_4  (
            .in0(N__23902),
            .in1(N__24202),
            .in2(N__21122),
            .in3(N__24436),
            .lcout(buf_readRTD_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i6_LC_7_8_5 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i6_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i6_LC_7_8_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i6_LC_7_8_5  (
            .in0(N__24108),
            .in1(N__24141),
            .in2(N__29515),
            .in3(N__21272),
            .lcout(\RTD.cfg_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_17_LC_7_8_6 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_17_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_17_LC_7_8_6 .LUT_INIT=16'b1110000010000000;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_17_LC_7_8_6  (
            .in0(N__24808),
            .in1(N__24435),
            .in2(N__24680),
            .in3(N__25038),
            .lcout(n11730),
            .ltout(n11730_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i15_LC_7_8_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i15_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i15_LC_7_8_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \RTD.READ_DATA_i15_LC_7_8_7  (
            .in0(N__24437),
            .in1(N__21311),
            .in2(N__21287),
            .in3(N__22231),
            .lcout(buf_readRTD_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43820),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i7_LC_7_9_0 .C_ON=1'b0;
    defparam \RTD.adress_i7_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i7_LC_7_9_0 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.adress_i7_LC_7_9_0  (
            .in0(N__25011),
            .in1(N__21284),
            .in2(N__24806),
            .in3(N__22390),
            .lcout(\RTD.adress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43806),
            .ce(N__21215),
            .sr(N__24518));
    defparam \RTD.i1_4_lut_adj_14_LC_7_9_1 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_14_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_14_LC_7_9_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i1_4_lut_adj_14_LC_7_9_1  (
            .in0(N__25360),
            .in1(N__21271),
            .in2(N__29508),
            .in3(N__21259),
            .lcout(),
            .ltout(\RTD.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i7_4_lut_LC_7_9_2 .C_ON=1'b0;
    defparam \RTD.i7_4_lut_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i7_4_lut_LC_7_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \RTD.i7_4_lut_LC_7_9_2  (
            .in0(N__22304),
            .in1(N__24914),
            .in2(N__21248),
            .in3(N__21155),
            .lcout(\RTD.adress_7_N_1340_7 ),
            .ltout(\RTD.adress_7_N_1340_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_LC_7_9_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_LC_7_9_3 .LUT_INIT=16'b0000000011110011;
    LogicCell40 \RTD.i1_2_lut_3_lut_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__24765),
            .in2(N__21245),
            .in3(N__25009),
            .lcout(\RTD.n20587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i0_LC_7_9_4 .C_ON=1'b0;
    defparam \RTD.adress_i0_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i0_LC_7_9_4 .LUT_INIT=16'b1011000111110101;
    LogicCell40 \RTD.adress_i0_LC_7_9_4  (
            .in0(N__25010),
            .in1(N__24799),
            .in2(N__21242),
            .in3(N__22389),
            .lcout(adress_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43806),
            .ce(N__21215),
            .sr(N__24518));
    defparam \RTD.i3_4_lut_adj_13_LC_7_9_5 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_adj_13_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_adj_13_LC_7_9_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i3_4_lut_adj_13_LC_7_9_5  (
            .in0(N__25204),
            .in1(N__21181),
            .in2(N__27506),
            .in3(N__21166),
            .lcout(\RTD.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4918_2_lut_LC_7_10_0 .C_ON=1'b0;
    defparam \RTD.i4918_2_lut_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i4918_2_lut_LC_7_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i4918_2_lut_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__24369),
            .in2(_gnd_net_),
            .in3(N__25012),
            .lcout(\RTD.n7333 ),
            .ltout(\RTD.n7333_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i3_4_lut_LC_7_10_1 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_LC_7_10_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \RTD.i3_4_lut_LC_7_10_1  (
            .in0(N__24666),
            .in1(N__24839),
            .in2(N__21353),
            .in3(N__22364),
            .lcout(\RTD.n11742 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i30_3_lut_4_lut_3_lut_LC_7_10_2 .C_ON=1'b0;
    defparam \RTD.i30_3_lut_4_lut_3_lut_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i30_3_lut_4_lut_3_lut_LC_7_10_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \RTD.i30_3_lut_4_lut_3_lut_LC_7_10_2  (
            .in0(N__24659),
            .in1(N__24793),
            .in2(_gnd_net_),
            .in3(N__25013),
            .lcout(),
            .ltout(\RTD.n13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i29_4_lut_LC_7_10_3 .C_ON=1'b0;
    defparam \RTD.i29_4_lut_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i29_4_lut_LC_7_10_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \RTD.i29_4_lut_LC_7_10_3  (
            .in0(N__24370),
            .in1(N__24660),
            .in2(N__21350),
            .in3(N__22615),
            .lcout(\RTD.n13228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i27_4_lut_4_lut_LC_7_10_5 .C_ON=1'b0;
    defparam \RTD.i27_4_lut_4_lut_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i27_4_lut_4_lut_LC_7_10_5 .LUT_INIT=16'b1110110100000010;
    LogicCell40 \RTD.i27_4_lut_4_lut_LC_7_10_5  (
            .in0(N__25014),
            .in1(N__24841),
            .in2(N__24682),
            .in3(N__24417),
            .lcout(\RTD.n11734 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19144_4_lut_4_lut_LC_7_10_6 .C_ON=1'b0;
    defparam \RTD.i19144_4_lut_4_lut_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i19144_4_lut_4_lut_LC_7_10_6 .LUT_INIT=16'b1101111110111111;
    LogicCell40 \RTD.i19144_4_lut_4_lut_LC_7_10_6  (
            .in0(N__24840),
            .in1(N__24371),
            .in2(N__24681),
            .in3(N__25015),
            .lcout(\RTD.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i1_LC_7_10_7 .C_ON=1'b0;
    defparam \RTD.adc_state_i1_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i1_LC_7_10_7 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \RTD.adc_state_i1_LC_7_10_7  (
            .in0(N__24794),
            .in1(N__21334),
            .in2(N__24683),
            .in3(N__22706),
            .lcout(adc_state_1_adj_1483),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43814),
            .ce(N__22683),
            .sr(_gnd_net_));
    defparam \RTD.cfg_tmp_i1_LC_7_11_0 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i1_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i1_LC_7_11_0 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i1_LC_7_11_0  (
            .in0(N__24420),
            .in1(N__27615),
            .in2(N__24863),
            .in3(N__21383),
            .lcout(\RTD.cfg_tmp_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i2_LC_7_11_1 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i2_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i2_LC_7_11_1 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \RTD.cfg_tmp_i2_LC_7_11_1  (
            .in0(N__21317),
            .in1(N__24801),
            .in2(N__25102),
            .in3(N__24427),
            .lcout(\RTD.cfg_tmp_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i3_LC_7_11_2 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i3_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i3_LC_7_11_2 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i3_LC_7_11_2  (
            .in0(N__24421),
            .in1(N__21428),
            .in2(N__24864),
            .in3(N__25197),
            .lcout(\RTD.cfg_tmp_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i4_LC_7_11_3 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i4_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i4_LC_7_11_3 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \RTD.cfg_tmp_i4_LC_7_11_3  (
            .in0(N__21422),
            .in1(N__24424),
            .in2(N__25256),
            .in3(N__24849),
            .lcout(\RTD.cfg_tmp_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i5_LC_7_11_4 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i5_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i5_LC_7_11_4 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i5_LC_7_11_4  (
            .in0(N__24422),
            .in1(N__27501),
            .in2(N__24865),
            .in3(N__21416),
            .lcout(\RTD.cfg_tmp_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i6_LC_7_11_5 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i6_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i6_LC_7_11_5 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \RTD.cfg_tmp_i6_LC_7_11_5  (
            .in0(N__21410),
            .in1(N__24425),
            .in2(N__29516),
            .in3(N__24850),
            .lcout(\RTD.cfg_tmp_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i7_LC_7_11_6 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i7_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i7_LC_7_11_6 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i7_LC_7_11_6  (
            .in0(N__24423),
            .in1(N__24065),
            .in2(N__24866),
            .in3(N__21404),
            .lcout(\RTD.cfg_tmp_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.cfg_tmp_i0_LC_7_11_7 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i0_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i0_LC_7_11_7 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \RTD.cfg_tmp_i0_LC_7_11_7  (
            .in0(N__21394),
            .in1(N__24800),
            .in2(N__25359),
            .in3(N__24426),
            .lcout(\RTD.cfg_tmp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43804),
            .ce(N__21377),
            .sr(N__21365));
    defparam \RTD.READ_DATA_i4_LC_7_12_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i4_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i4_LC_7_12_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i4_LC_7_12_0  (
            .in0(N__24218),
            .in1(N__21478),
            .in2(N__38182),
            .in3(N__24442),
            .lcout(buf_readRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i2_LC_7_12_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i2_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i2_LC_7_12_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i2_LC_7_12_1  (
            .in0(N__24439),
            .in1(N__46891),
            .in2(N__21608),
            .in3(N__24219),
            .lcout(buf_readRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i4_LC_7_12_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i4_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i4_LC_7_12_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i4_LC_7_12_2  (
            .in0(N__22165),
            .in1(N__21477),
            .in2(N__21586),
            .in3(N__21519),
            .lcout(read_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i7_LC_7_12_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i7_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i7_LC_7_12_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i7_LC_7_12_3  (
            .in0(N__24441),
            .in1(N__35653),
            .in2(N__21629),
            .in3(N__24221),
            .lcout(buf_readRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i3_LC_7_12_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i3_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i3_LC_7_12_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.read_buf_i3_LC_7_12_4  (
            .in0(N__22164),
            .in1(N__21606),
            .in2(N__21585),
            .in3(N__21518),
            .lcout(read_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i5_LC_7_12_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i5_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i5_LC_7_12_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i5_LC_7_12_5  (
            .in0(N__24440),
            .in1(N__21463),
            .in2(N__43600),
            .in3(N__24220),
            .lcout(buf_readRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_adj_9_LC_7_12_6 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_adj_9_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_adj_9_LC_7_12_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RTD.i2_3_lut_adj_9_LC_7_12_6  (
            .in0(N__24848),
            .in1(N__24584),
            .in2(_gnd_net_),
            .in3(N__24438),
            .lcout(n1_adj_1601),
            .ltout(n1_adj_1601_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i5_LC_7_12_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i5_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i5_LC_7_12_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.read_buf_i5_LC_7_12_7  (
            .in0(N__21479),
            .in1(N__21462),
            .in2(N__21467),
            .in3(N__22166),
            .lcout(read_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43759),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_7_13_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_7_13_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i26_LC_7_13_1  (
            .in0(N__22950),
            .in1(N__52849),
            .in2(N__21667),
            .in3(N__52047),
            .lcout(cmd_rdadctmp_26_adj_1424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57923),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i15_LC_7_13_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i15_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i15_LC_7_13_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i15_LC_7_13_3  (
            .in0(N__53127),
            .in1(N__52846),
            .in2(N__21704),
            .in3(N__44949),
            .lcout(buf_adcdata_iac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57923),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i21_LC_7_13_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i21_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i21_LC_7_13_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i21_LC_7_13_5  (
            .in0(N__53128),
            .in1(N__52847),
            .in2(N__21449),
            .in3(N__22881),
            .lcout(buf_adcdata_iac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57923),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_7_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_7_13_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i31_LC_7_13_6  (
            .in0(N__52046),
            .in1(N__21736),
            .in2(N__22930),
            .in3(N__52854),
            .lcout(cmd_rdadctmp_31_adj_1419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57923),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i22_LC_7_13_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i22_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i22_LC_7_13_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i22_LC_7_13_7  (
            .in0(N__53129),
            .in1(N__52848),
            .in2(N__21740),
            .in3(N__36795),
            .lcout(buf_adcdata_iac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57923),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_7_14_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_7_14_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i27_LC_7_14_0  (
            .in0(N__52880),
            .in1(N__25296),
            .in2(N__21668),
            .in3(N__52003),
            .lcout(cmd_rdadctmp_27_adj_1423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i16_LC_7_14_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i16_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i16_LC_7_14_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i16_LC_7_14_1  (
            .in0(N__53068),
            .in1(N__52875),
            .in2(N__21686),
            .in3(N__22782),
            .lcout(buf_adcdata_iac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.MOSI_31_LC_7_14_2 .C_ON=1'b0;
    defparam \CLK_DDS.MOSI_31_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.MOSI_31_LC_7_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CLK_DDS.MOSI_31_LC_7_14_2  (
            .in0(N__23533),
            .in1(N__21715),
            .in2(_gnd_net_),
            .in3(N__23342),
            .lcout(DDS_MOSI1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_7_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_7_14_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i23_LC_7_14_3  (
            .in0(N__21699),
            .in1(N__52877),
            .in2(N__30881),
            .in3(N__52004),
            .lcout(cmd_rdadctmp_23_adj_1427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_7_14_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_7_14_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i24_LC_7_14_5  (
            .in0(N__21700),
            .in1(N__52878),
            .in2(N__21685),
            .in3(N__52005),
            .lcout(cmd_rdadctmp_24_adj_1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_7_14_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_7_14_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i25_LC_7_14_6  (
            .in0(N__52879),
            .in1(N__21681),
            .in2(N__22954),
            .in3(N__52002),
            .lcout(cmd_rdadctmp_25_adj_1425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i18_LC_7_14_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i18_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i18_LC_7_14_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i18_LC_7_14_7  (
            .in0(N__53069),
            .in1(N__52876),
            .in2(N__27447),
            .in3(N__21666),
            .lcout(buf_adcdata_iac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57936),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i5_LC_7_15_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i5_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i5_LC_7_15_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i5_LC_7_15_1  (
            .in0(N__23333),
            .in1(N__23497),
            .in2(N__21785),
            .in3(N__36302),
            .lcout(\CLK_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57947),
            .ce(N__23145),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i2_LC_7_15_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i2_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i2_LC_7_15_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i2_LC_7_15_5  (
            .in0(N__23331),
            .in1(N__23496),
            .in2(N__21647),
            .in3(N__27884),
            .lcout(\CLK_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57947),
            .ce(N__23145),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i3_LC_7_15_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i3_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i3_LC_7_15_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i3_LC_7_15_6  (
            .in0(N__23495),
            .in1(N__23334),
            .in2(N__21803),
            .in3(N__27656),
            .lcout(\CLK_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57947),
            .ce(N__23145),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i4_LC_7_15_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i4_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i4_LC_7_15_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \CLK_DDS.tmp_buf_i4_LC_7_15_7  (
            .in0(N__23332),
            .in1(N__25745),
            .in2(N__21794),
            .in3(N__23498),
            .lcout(\CLK_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57947),
            .ce(N__23145),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i6_LC_7_16_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i6_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i6_LC_7_16_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \CLK_DDS.tmp_buf_i6_LC_7_16_2  (
            .in0(N__21776),
            .in1(N__23494),
            .in2(N__31286),
            .in3(N__23326),
            .lcout(\CLK_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57959),
            .ce(N__23144),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i7_LC_7_16_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i7_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i7_LC_7_16_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i7_LC_7_16_3  (
            .in0(N__23325),
            .in1(N__23499),
            .in2(N__21770),
            .in3(N__44588),
            .lcout(\CLK_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57959),
            .ce(N__23144),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i8_LC_7_16_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i8_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i8_LC_7_16_4 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i8_LC_7_16_4  (
            .in0(N__21761),
            .in1(N__23327),
            .in2(N__23513),
            .in3(N__25592),
            .lcout(\CLK_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57959),
            .ce(N__23144),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i23_4_lut_LC_7_16_6 .C_ON=1'b0;
    defparam \CLK_DDS.i23_4_lut_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i23_4_lut_LC_7_16_6 .LUT_INIT=16'b1110111000010011;
    LogicCell40 \CLK_DDS.i23_4_lut_LC_7_16_6  (
            .in0(N__22575),
            .in1(N__23323),
            .in2(N__23121),
            .in3(N__23490),
            .lcout(\CLK_DDS.n9_adj_1395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19153_4_lut_LC_7_16_7 .C_ON=1'b0;
    defparam \CLK_DDS.i19153_4_lut_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19153_4_lut_LC_7_16_7 .LUT_INIT=16'b1111101111111110;
    LogicCell40 \CLK_DDS.i19153_4_lut_LC_7_16_7  (
            .in0(N__23324),
            .in1(N__22576),
            .in2(N__23512),
            .in3(N__23114),
            .lcout(\CLK_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_8_2_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_8_2_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i12_LC_8_2_0  (
            .in0(N__25968),
            .in1(N__34454),
            .in2(N__28835),
            .in3(N__35305),
            .lcout(cmd_rdadctmp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57809),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i4_LC_8_3_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i4_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i4_LC_8_3_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i4_LC_8_3_0  (
            .in0(N__25972),
            .in1(N__34658),
            .in2(N__35423),
            .in3(N__21886),
            .lcout(buf_adcdata_vac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57814),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i4_LC_8_3_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i4_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i4_LC_8_3_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i4_LC_8_3_1  (
            .in0(N__53185),
            .in1(N__52996),
            .in2(N__28763),
            .in3(N__21862),
            .lcout(buf_adcdata_iac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57814),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_5_i22_3_lut_LC_8_3_2.C_ON=1'b0;
    defparam mux_136_Mux_5_i22_3_lut_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_5_i22_3_lut_LC_8_3_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_136_Mux_5_i22_3_lut_LC_8_3_2 (
            .in0(N__21983),
            .in1(N__25861),
            .in2(_gnd_net_),
            .in3(N__49056),
            .lcout(n22_adj_1632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_4_i19_3_lut_LC_8_3_4.C_ON=1'b0;
    defparam mux_136_Mux_4_i19_3_lut_LC_8_3_4.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_4_i19_3_lut_LC_8_3_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_136_Mux_4_i19_3_lut_LC_8_3_4 (
            .in0(N__22043),
            .in1(N__21885),
            .in2(_gnd_net_),
            .in3(N__56358),
            .lcout(),
            .ltout(n19_adj_1636_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_4_i22_3_lut_LC_8_3_5.C_ON=1'b0;
    defparam mux_136_Mux_4_i22_3_lut_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_4_i22_3_lut_LC_8_3_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_136_Mux_4_i22_3_lut_LC_8_3_5 (
            .in0(N__49057),
            .in1(_gnd_net_),
            .in2(N__21872),
            .in3(N__21861),
            .lcout(),
            .ltout(n22_adj_1637_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_4_i30_3_lut_LC_8_3_6.C_ON=1'b0;
    defparam mux_136_Mux_4_i30_3_lut_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_4_i30_3_lut_LC_8_3_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_136_Mux_4_i30_3_lut_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(N__21848),
            .in2(N__21836),
            .in3(N__48669),
            .lcout(n30_adj_1638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_8_4_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_8_4_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i16_LC_8_4_0  (
            .in0(N__35368),
            .in1(N__21994),
            .in2(N__30576),
            .in3(N__34337),
            .lcout(cmd_rdadctmp_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_8_4_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_8_4_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i5_LC_8_4_1  (
            .in0(N__34338),
            .in1(N__35372),
            .in2(N__21815),
            .in3(N__21833),
            .lcout(cmd_rdadctmp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i21_LC_8_4_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i21_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i21_LC_8_4_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i21_LC_8_4_2  (
            .in0(N__35366),
            .in1(N__34657),
            .in2(N__21923),
            .in3(N__25470),
            .lcout(buf_adcdata_vac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i7_LC_8_4_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i7_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i7_LC_8_4_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i7_LC_8_4_3  (
            .in0(N__34656),
            .in1(N__35371),
            .in2(N__21998),
            .in3(N__23650),
            .lcout(buf_adcdata_vac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_8_4_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_8_4_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i6_LC_8_4_4  (
            .in0(N__35369),
            .in1(N__21814),
            .in2(N__25921),
            .in3(N__34339),
            .lcout(cmd_rdadctmp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i6_LC_8_4_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i6_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i6_LC_8_4_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i6_LC_8_4_5  (
            .in0(N__34655),
            .in1(N__35370),
            .in2(N__23590),
            .in3(N__23695),
            .lcout(buf_adcdata_vac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_8_4_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_8_4_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i15_LC_8_4_6  (
            .in0(N__35367),
            .in1(N__21993),
            .in2(N__23696),
            .in3(N__34336),
            .lcout(cmd_rdadctmp_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57818),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_5_i19_3_lut_LC_8_4_7.C_ON=1'b0;
    defparam mux_136_Mux_5_i19_3_lut_LC_8_4_7.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_5_i19_3_lut_LC_8_4_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_136_Mux_5_i19_3_lut_LC_8_4_7 (
            .in0(N__21969),
            .in1(N__56295),
            .in2(_gnd_net_),
            .in3(N__22058),
            .lcout(n19_adj_1631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i5_LC_8_5_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i5_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i5_LC_8_5_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i5_LC_8_5_0  (
            .in0(N__35361),
            .in1(N__34661),
            .in2(N__25952),
            .in3(N__21973),
            .lcout(buf_adcdata_vac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57822),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i23_LC_8_5_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i23_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i23_LC_8_5_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i23_LC_8_5_1  (
            .in0(N__34660),
            .in1(N__35364),
            .in2(N__22073),
            .in3(N__22263),
            .lcout(buf_adcdata_vac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57822),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3 .LUT_INIT=16'b1101000011000000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_LC_8_5_3  (
            .in0(N__32897),
            .in1(N__33237),
            .in2(N__33124),
            .in3(N__33491),
            .lcout(n13109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22202_bdd_4_lut_LC_8_5_4.C_ON=1'b0;
    defparam n22202_bdd_4_lut_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam n22202_bdd_4_lut_LC_8_5_4.LUT_INIT=16'b1010101011100100;
    LogicCell40 n22202_bdd_4_lut_LC_8_5_4 (
            .in0(N__25397),
            .in1(N__21943),
            .in2(N__22028),
            .in3(N__48419),
            .lcout(n22205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i22_LC_8_5_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i22_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i22_LC_8_5_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i22_LC_8_5_5  (
            .in0(N__34659),
            .in1(N__35363),
            .in2(N__31965),
            .in3(N__22087),
            .lcout(buf_adcdata_vac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57822),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_8_5_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_8_5_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i30_LC_8_5_6  (
            .in0(N__35362),
            .in1(N__21922),
            .in2(N__22088),
            .in3(N__34439),
            .lcout(cmd_rdadctmp_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57822),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_8_5_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_8_5_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i31_LC_8_5_7  (
            .in0(N__34440),
            .in1(N__22086),
            .in2(N__22072),
            .in3(N__35365),
            .lcout(cmd_rdadctmp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57822),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i5_LC_8_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i5_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i5_LC_8_6_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i5_LC_8_6_0  (
            .in0(N__33294),
            .in1(N__22054),
            .in2(N__29162),
            .in3(N__26744),
            .lcout(buf_adcdata_vdc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i10_LC_8_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i10_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i10_LC_8_6_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \ADC_VDC.ADC_DATA_i10_LC_8_6_1  (
            .in0(N__30484),
            .in1(N__33295),
            .in2(N__26552),
            .in3(N__29124),
            .lcout(buf_adcdata_vdc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i4_LC_8_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i4_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i4_LC_8_6_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i4_LC_8_6_2  (
            .in0(N__33293),
            .in1(N__22039),
            .in2(N__29161),
            .in3(N__26786),
            .lcout(buf_adcdata_vdc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i17_LC_8_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i17_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i17_LC_8_6_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \ADC_VDC.ADC_DATA_i17_LC_8_6_3  (
            .in0(N__43978),
            .in1(N__29125),
            .in2(N__26903),
            .in3(N__33296),
            .lcout(buf_adcdata_vdc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i20_LC_8_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i20_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i20_LC_8_6_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i20_LC_8_6_4  (
            .in0(N__33291),
            .in1(N__22021),
            .in2(N__29159),
            .in3(N__27239),
            .lcout(buf_adcdata_vdc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i6_LC_8_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i6_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i6_LC_8_6_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \ADC_VDC.ADC_DATA_i6_LC_8_6_5  (
            .in0(N__23557),
            .in1(N__33298),
            .in2(N__26705),
            .in3(N__29127),
            .lcout(buf_adcdata_vdc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i3_LC_8_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i3_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i3_LC_8_6_6 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i3_LC_8_6_6  (
            .in0(N__33292),
            .in1(N__28510),
            .in2(N__29160),
            .in3(N__26825),
            .lcout(buf_adcdata_vdc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i21_LC_8_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i21_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i21_LC_8_6_7 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \ADC_VDC.ADC_DATA_i21_LC_8_6_7  (
            .in0(N__25435),
            .in1(N__29126),
            .in2(N__27218),
            .in3(N__33297),
            .lcout(buf_adcdata_vdc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40112),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i0_LC_8_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i0_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i0_LC_8_7_0 .LUT_INIT=16'b0000000001110110;
    LogicCell40 \ADC_VDC.adc_state_i0_LC_8_7_0  (
            .in0(N__33344),
            .in1(N__33086),
            .in2(N__33614),
            .in3(N__33477),
            .lcout(\ADC_VDC.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40136),
            .ce(N__22010),
            .sr(_gnd_net_));
    defparam i15243_2_lut_3_lut_LC_8_7_1.C_ON=1'b0;
    defparam i15243_2_lut_3_lut_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam i15243_2_lut_3_lut_LC_8_7_1.LUT_INIT=16'b0000000000001010;
    LogicCell40 i15243_2_lut_3_lut_LC_8_7_1 (
            .in0(N__37981),
            .in1(_gnd_net_),
            .in2(N__54172),
            .in3(N__52436),
            .lcout(n14_adj_1579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15253_2_lut_3_lut_LC_8_7_2.C_ON=1'b0;
    defparam i15253_2_lut_3_lut_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam i15253_2_lut_3_lut_LC_8_7_2.LUT_INIT=16'b0001000100000000;
    LogicCell40 i15253_2_lut_3_lut_LC_8_7_2 (
            .in0(N__52437),
            .in1(N__54145),
            .in2(_gnd_net_),
            .in3(N__43149),
            .lcout(n14_adj_1570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15255_2_lut_3_lut_LC_8_7_4.C_ON=1'b0;
    defparam i15255_2_lut_3_lut_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam i15255_2_lut_3_lut_LC_8_7_4.LUT_INIT=16'b0001000100000000;
    LogicCell40 i15255_2_lut_3_lut_LC_8_7_4 (
            .in0(N__52435),
            .in1(N__54141),
            .in2(_gnd_net_),
            .in3(N__44291),
            .lcout(n14_adj_1572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15256_2_lut_3_lut_LC_8_7_5.C_ON=1'b0;
    defparam i15256_2_lut_3_lut_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam i15256_2_lut_3_lut_LC_8_7_5.LUT_INIT=16'b0000000000001010;
    LogicCell40 i15256_2_lut_3_lut_LC_8_7_5 (
            .in0(N__42971),
            .in1(_gnd_net_),
            .in2(N__54173),
            .in3(N__52439),
            .lcout(n14_adj_1573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15257_2_lut_3_lut_LC_8_7_6.C_ON=1'b0;
    defparam i15257_2_lut_3_lut_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam i15257_2_lut_3_lut_LC_8_7_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15257_2_lut_3_lut_LC_8_7_6 (
            .in0(N__52438),
            .in1(N__45545),
            .in2(_gnd_net_),
            .in3(N__54149),
            .lcout(n14_adj_1574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.SCLK_51_LC_8_8_0 .C_ON=1'b0;
    defparam \RTD.SCLK_51_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.SCLK_51_LC_8_8_0 .LUT_INIT=16'b0011100100011100;
    LogicCell40 \RTD.SCLK_51_LC_8_8_0  (
            .in0(N__24805),
            .in1(N__24434),
            .in2(N__24679),
            .in3(N__25034),
            .lcout(RTD_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43816),
            .ce(N__22181),
            .sr(_gnd_net_));
    defparam \RTD.i19171_4_lut_4_lut_LC_8_8_2 .C_ON=1'b0;
    defparam \RTD.i19171_4_lut_4_lut_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i19171_4_lut_4_lut_LC_8_8_2 .LUT_INIT=16'b1100011110111000;
    LogicCell40 \RTD.i19171_4_lut_4_lut_LC_8_8_2  (
            .in0(N__24802),
            .in1(N__24431),
            .in2(N__24677),
            .in3(N__25031),
            .lcout(\RTD.n11756 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_3_lut_4_lut_LC_8_8_3 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_LC_8_8_3 .LUT_INIT=16'b1101000010000110;
    LogicCell40 \RTD.i1_3_lut_4_lut_LC_8_8_3  (
            .in0(N__25030),
            .in1(N__24644),
            .in2(N__24467),
            .in3(N__24803),
            .lcout(\RTD.n15081 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_16_LC_8_8_4 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_16_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_16_LC_8_8_4 .LUT_INIT=16'b1100000010110001;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_16_LC_8_8_4  (
            .in0(N__24804),
            .in1(N__24433),
            .in2(N__24678),
            .in3(N__25033),
            .lcout(n13309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19100_3_lut_3_lut_LC_8_8_6 .C_ON=1'b0;
    defparam \RTD.i19100_3_lut_3_lut_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i19100_3_lut_3_lut_LC_8_8_6 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \RTD.i19100_3_lut_3_lut_LC_8_8_6  (
            .in0(N__24648),
            .in1(N__24432),
            .in2(_gnd_net_),
            .in3(N__25032),
            .lcout(\RTD.n11703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_15_LC_8_9_1 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_15_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_15_LC_8_9_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \RTD.i1_2_lut_adj_15_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__22430),
            .in2(_gnd_net_),
            .in3(N__22388),
            .lcout(\RTD.n16669 ),
            .ltout(\RTD.n16669_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.CS_52_LC_8_9_2 .C_ON=1'b0;
    defparam \RTD.CS_52_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.CS_52_LC_8_9_2 .LUT_INIT=16'b0000001101110111;
    LogicCell40 \RTD.CS_52_LC_8_9_2  (
            .in0(N__25039),
            .in1(N__24658),
            .in2(N__22358),
            .in3(N__24797),
            .lcout(RTD_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43780),
            .ce(N__22334),
            .sr(_gnd_net_));
    defparam \RTD.i4_4_lut_LC_8_9_3 .C_ON=1'b0;
    defparam \RTD.i4_4_lut_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i4_4_lut_LC_8_9_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i4_4_lut_LC_8_9_3  (
            .in0(N__24022),
            .in1(N__24063),
            .in2(N__27622),
            .in3(N__22315),
            .lcout(\RTD.n12_adj_1397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16108_3_lut_LC_8_9_4 .C_ON=1'b0;
    defparam \ADC_VDC.i16108_3_lut_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16108_3_lut_LC_8_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \ADC_VDC.i16108_3_lut_LC_8_9_4  (
            .in0(N__22298),
            .in1(N__22264),
            .in2(_gnd_net_),
            .in3(N__56248),
            .lcout(),
            .ltout(n19_adj_1526_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19474_LC_8_9_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19474_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19474_LC_8_9_5.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19474_LC_8_9_5 (
            .in0(N__22220),
            .in1(N__48398),
            .in2(N__22244),
            .in3(N__49054),
            .lcout(),
            .ltout(n22076_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22076_bdd_4_lut_LC_8_9_6.C_ON=1'b0;
    defparam n22076_bdd_4_lut_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam n22076_bdd_4_lut_LC_8_9_6.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22076_bdd_4_lut_LC_8_9_6 (
            .in0(N__49055),
            .in1(N__24491),
            .in2(N__22241),
            .in3(N__22805),
            .lcout(n22079),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_7_i20_3_lut_LC_8_9_7.C_ON=1'b0;
    defparam mux_134_Mux_7_i20_3_lut_LC_8_9_7.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i20_3_lut_LC_8_9_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_134_Mux_7_i20_3_lut_LC_8_9_7 (
            .in0(N__56247),
            .in1(N__22238),
            .in2(_gnd_net_),
            .in3(N__24062),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i0_LC_8_10_0 .C_ON=1'b0;
    defparam \RTD.adc_state_i0_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i0_LC_8_10_0 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \RTD.adc_state_i0_LC_8_10_0  (
            .in0(N__22652),
            .in1(N__22214),
            .in2(N__24675),
            .in3(N__22727),
            .lcout(\RTD.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43740),
            .ce(N__22684),
            .sr(_gnd_net_));
    defparam \RTD.i19088_2_lut_LC_8_10_1 .C_ON=1'b0;
    defparam \RTD.i19088_2_lut_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i19088_2_lut_LC_8_10_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \RTD.i19088_2_lut_LC_8_10_1  (
            .in0(N__25017),
            .in1(N__33845),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\RTD.n21323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i45_4_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \RTD.i45_4_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i45_4_lut_LC_8_10_2 .LUT_INIT=16'b0111001000100010;
    LogicCell40 \RTD.i45_4_lut_LC_8_10_2  (
            .in0(N__24411),
            .in1(N__22632),
            .in2(N__22655),
            .in3(N__31703),
            .lcout(\RTD.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19023_4_lut_LC_8_10_3 .C_ON=1'b0;
    defparam \RTD.i19023_4_lut_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i19023_4_lut_LC_8_10_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \RTD.i19023_4_lut_LC_8_10_3  (
            .in0(N__22643),
            .in1(N__24636),
            .in2(N__22468),
            .in3(N__22721),
            .lcout(),
            .ltout(\RTD.n21325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i2_LC_8_10_4 .C_ON=1'b0;
    defparam \RTD.adc_state_i2_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i2_LC_8_10_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.adc_state_i2_LC_8_10_4  (
            .in0(N__24413),
            .in1(N__22633),
            .in2(N__22646),
            .in3(N__24635),
            .lcout(adc_state_2_adj_1482),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43740),
            .ce(N__22684),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_12_LC_8_10_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_12_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_12_LC_8_10_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \RTD.i1_2_lut_adj_12_LC_8_10_5  (
            .in0(N__25018),
            .in1(_gnd_net_),
            .in2(N__24807),
            .in3(_gnd_net_),
            .lcout(\RTD.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4948_2_lut_LC_8_10_6 .C_ON=1'b0;
    defparam \RTD.i4948_2_lut_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i4948_2_lut_LC_8_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i4948_2_lut_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__24769),
            .in2(_gnd_net_),
            .in3(N__25016),
            .lcout(\RTD.n1 ),
            .ltout(\RTD.n1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i22_4_lut_4_lut_LC_8_10_7 .C_ON=1'b0;
    defparam \RTD.i22_4_lut_4_lut_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i22_4_lut_4_lut_LC_8_10_7 .LUT_INIT=16'b1001000110000000;
    LogicCell40 \RTD.i22_4_lut_4_lut_LC_8_10_7  (
            .in0(N__24634),
            .in1(N__24412),
            .in2(N__22619),
            .in3(N__22616),
            .lcout(\RTD.n13192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i0_LC_8_11_1 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i0_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i0_LC_8_11_1 .LUT_INIT=16'b1010001100000011;
    LogicCell40 \CLK_DDS.dds_state_i0_LC_8_11_1  (
            .in0(N__22604),
            .in1(N__22532),
            .in2(N__23360),
            .in3(N__22595),
            .lcout(dds_state_0_adj_1454),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57881),
            .ce(N__22493),
            .sr(_gnd_net_));
    defparam \RTD.i18725_4_lut_LC_8_11_3 .C_ON=1'b0;
    defparam \RTD.i18725_4_lut_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i18725_4_lut_LC_8_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \RTD.i18725_4_lut_LC_8_11_3  (
            .in0(N__24409),
            .in1(N__25019),
            .in2(N__22469),
            .in3(N__22720),
            .lcout(),
            .ltout(\RTD.n21276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19037_3_lut_LC_8_11_4 .C_ON=1'b0;
    defparam \RTD.i19037_3_lut_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19037_3_lut_LC_8_11_4 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \RTD.i19037_3_lut_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__24795),
            .in2(N__22730),
            .in3(N__24928),
            .lcout(\RTD.n21275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_LC_8_11_6 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_LC_8_11_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \RTD.i1_2_lut_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__33840),
            .in2(_gnd_net_),
            .in3(N__31701),
            .lcout(\RTD.adc_state_3_N_1368_1 ),
            .ltout(\RTD.adc_state_3_N_1368_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_8_11_7 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_8_11_7 .LUT_INIT=16'b1011100111101110;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_8_11_7  (
            .in0(N__24410),
            .in1(N__24798),
            .in2(N__22709),
            .in3(N__25020),
            .lcout(\RTD.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i3_LC_8_12_0 .C_ON=1'b0;
    defparam \RTD.adc_state_i3_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i3_LC_8_12_0 .LUT_INIT=16'b0100010001000111;
    LogicCell40 \RTD.adc_state_i3_LC_8_12_0  (
            .in0(N__24466),
            .in1(N__24591),
            .in2(N__22700),
            .in3(N__24929),
            .lcout(adc_state_3_adj_1481),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43758),
            .ce(N__22685),
            .sr(_gnd_net_));
    defparam i15266_2_lut_3_lut_LC_8_12_1.C_ON=1'b0;
    defparam i15266_2_lut_3_lut_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam i15266_2_lut_3_lut_LC_8_12_1.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15266_2_lut_3_lut_LC_8_12_1 (
            .in0(N__41499),
            .in1(N__54171),
            .in2(_gnd_net_),
            .in3(N__52433),
            .lcout(n14_adj_1545),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_3_i16_3_lut_LC_8_12_3.C_ON=1'b0;
    defparam mux_135_Mux_3_i16_3_lut_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_3_i16_3_lut_LC_8_12_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 mux_135_Mux_3_i16_3_lut_LC_8_12_3 (
            .in0(N__28287),
            .in1(_gnd_net_),
            .in2(N__27655),
            .in3(N__56286),
            .lcout(),
            .ltout(n16_adj_1512_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18264_3_lut_LC_8_12_4.C_ON=1'b0;
    defparam i18264_3_lut_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam i18264_3_lut_LC_8_12_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 i18264_3_lut_LC_8_12_4 (
            .in0(N__53230),
            .in1(_gnd_net_),
            .in2(N__22658),
            .in3(N__48374),
            .lcout(n20878),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18225_3_lut_LC_8_12_5.C_ON=1'b0;
    defparam i18225_3_lut_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam i18225_3_lut_LC_8_12_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 i18225_3_lut_LC_8_12_5 (
            .in0(N__23011),
            .in1(N__56287),
            .in2(_gnd_net_),
            .in3(N__32345),
            .lcout(n20839),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_218_LC_8_12_7.C_ON=1'b0;
    defparam i1_3_lut_adj_218_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_218_LC_8_12_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_3_lut_adj_218_LC_8_12_7 (
            .in0(N__53591),
            .in1(N__48503),
            .in2(_gnd_net_),
            .in3(N__31882),
            .lcout(n20670),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i3_LC_8_13_0.C_ON=1'b0;
    defparam buf_dds0_i3_LC_8_13_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i3_LC_8_13_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i3_LC_8_13_0 (
            .in0(N__49871),
            .in1(N__28288),
            .in2(N__37985),
            .in3(N__38967),
            .lcout(buf_dds0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57910),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i17_LC_8_13_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i17_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i17_LC_8_13_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i17_LC_8_13_1  (
            .in0(N__53130),
            .in1(N__52845),
            .in2(N__22955),
            .in3(N__25545),
            .lcout(buf_adcdata_iac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57910),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i8_LC_8_13_2.C_ON=1'b0;
    defparam buf_device_acadc_i8_LC_8_13_2.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i8_LC_8_13_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_device_acadc_i8_LC_8_13_2 (
            .in0(N__41370),
            .in1(N__46059),
            .in2(N__49915),
            .in3(N__22819),
            .lcout(VAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57910),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i6_LC_8_13_3.C_ON=1'b0;
    defparam buf_device_acadc_i6_LC_8_13_3.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i6_LC_8_13_3.LUT_INIT=16'b0010001011100010;
    LogicCell40 buf_device_acadc_i6_LC_8_13_3 (
            .in0(N__22906),
            .in1(N__41371),
            .in2(N__46421),
            .in3(N__49875),
            .lcout(VAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57910),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i23_LC_8_13_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i23_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i23_LC_8_13_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i23_LC_8_13_4  (
            .in0(N__52844),
            .in1(N__53131),
            .in2(N__22931),
            .in3(N__22849),
            .lcout(buf_adcdata_iac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57910),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19469_LC_8_13_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19469_LC_8_13_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19469_LC_8_13_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19469_LC_8_13_5 (
            .in0(N__22905),
            .in1(N__48373),
            .in2(N__22882),
            .in3(N__56246),
            .lcout(n22100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14314_3_lut_LC_8_13_6.C_ON=1'b0;
    defparam i14314_3_lut_LC_8_13_6.SEQ_MODE=4'b0000;
    defparam i14314_3_lut_LC_8_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i14314_3_lut_LC_8_13_6 (
            .in0(N__56245),
            .in1(N__22848),
            .in2(_gnd_net_),
            .in3(N__22818),
            .lcout(n17_adj_1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19444_LC_8_14_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19444_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19444_LC_8_14_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19444_LC_8_14_0 (
            .in0(N__22743),
            .in1(N__48375),
            .in2(N__22783),
            .in3(N__56304),
            .lcout(n22040),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i1_LC_8_14_2.C_ON=1'b0;
    defparam buf_device_acadc_i1_LC_8_14_2.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i1_LC_8_14_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 buf_device_acadc_i1_LC_8_14_2 (
            .in0(N__22744),
            .in1(N__44477),
            .in2(_gnd_net_),
            .in3(N__41388),
            .lcout(IAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57924),
            .ce(),
            .sr(_gnd_net_));
    defparam n22100_bdd_4_lut_LC_8_14_3.C_ON=1'b0;
    defparam n22100_bdd_4_lut_LC_8_14_3.SEQ_MODE=4'b0000;
    defparam n22100_bdd_4_lut_LC_8_14_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22100_bdd_4_lut_LC_8_14_3 (
            .in0(N__48376),
            .in1(N__28117),
            .in2(N__23033),
            .in3(N__30994),
            .lcout(n22103),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i5_LC_8_14_4.C_ON=1'b0;
    defparam buf_control_i5_LC_8_14_4.SEQ_MODE=4'b1000;
    defparam buf_control_i5_LC_8_14_4.LUT_INIT=16'b0010111000100010;
    LogicCell40 buf_control_i5_LC_8_14_4 (
            .in0(N__30942),
            .in1(N__44430),
            .in2(N__49925),
            .in3(N__46406),
            .lcout(AMPV_POW),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57924),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i7_LC_8_14_5.C_ON=1'b0;
    defparam buf_cfgRTD_i7_LC_8_14_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i7_LC_8_14_5.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_cfgRTD_i7_LC_8_14_5 (
            .in0(N__28979),
            .in1(N__49910),
            .in2(N__46067),
            .in3(N__24047),
            .lcout(buf_cfgRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57924),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i2_LC_8_14_6.C_ON=1'b0;
    defparam buf_control_i2_LC_8_14_6.SEQ_MODE=4'b1000;
    defparam buf_control_i2_LC_8_14_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i2_LC_8_14_6 (
            .in0(N__49909),
            .in1(N__44429),
            .in2(N__43005),
            .in3(N__23007),
            .lcout(SELIRNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57924),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_4_i16_3_lut_LC_8_14_7.C_ON=1'b0;
    defparam mux_135_Mux_4_i16_3_lut_LC_8_14_7.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_4_i16_3_lut_LC_8_14_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_135_Mux_4_i16_3_lut_LC_8_14_7 (
            .in0(N__56305),
            .in1(N__25740),
            .in2(_gnd_net_),
            .in3(N__28414),
            .lcout(n16_adj_1508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i10_LC_8_15_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i10_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i10_LC_8_15_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i10_LC_8_15_0  (
            .in0(N__23335),
            .in1(N__23506),
            .in2(N__23186),
            .in3(N__25798),
            .lcout(\CLK_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i11_LC_8_15_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i11_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i11_LC_8_15_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i11_LC_8_15_1  (
            .in0(N__23503),
            .in1(N__23339),
            .in2(N__22988),
            .in3(N__40483),
            .lcout(\CLK_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i12_LC_8_15_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i12_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i12_LC_8_15_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i12_LC_8_15_2  (
            .in0(N__23336),
            .in1(N__23507),
            .in2(N__22979),
            .in3(N__40293),
            .lcout(\CLK_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i13_LC_8_15_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i13_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i13_LC_8_15_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i13_LC_8_15_4  (
            .in0(N__23337),
            .in1(N__23508),
            .in2(N__22970),
            .in3(N__30995),
            .lcout(\CLK_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i14_LC_8_15_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i14_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i14_LC_8_15_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \CLK_DDS.tmp_buf_i14_LC_8_15_5  (
            .in0(N__23504),
            .in1(N__23340),
            .in2(N__36964),
            .in3(N__22961),
            .lcout(\CLK_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i15_LC_8_15_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i15_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i15_LC_8_15_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i15_LC_8_15_6  (
            .in0(N__23338),
            .in1(N__23509),
            .in2(N__23546),
            .in3(N__25280),
            .lcout(tmp_buf_15_adj_1455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i9_LC_8_15_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i9_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i9_LC_8_15_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i9_LC_8_15_7  (
            .in0(N__23505),
            .in1(N__23341),
            .in2(N__23195),
            .in3(N__25609),
            .lcout(\CLK_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57937),
            .ce(N__23169),
            .sr(_gnd_net_));
    defparam trig_dds1_315_LC_8_16_0.C_ON=1'b0;
    defparam trig_dds1_315_LC_8_16_0.SEQ_MODE=4'b1000;
    defparam trig_dds1_315_LC_8_16_0.LUT_INIT=16'b0110000001100100;
    LogicCell40 trig_dds1_315_LC_8_16_0 (
            .in0(N__49904),
            .in1(N__54981),
            .in2(N__23125),
            .in3(N__34796),
            .lcout(trig_dds1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57948),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_219_LC_8_16_1.C_ON=1'b0;
    defparam i1_4_lut_adj_219_LC_8_16_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_219_LC_8_16_1.LUT_INIT=16'b1100000011010000;
    LogicCell40 i1_4_lut_adj_219_LC_8_16_1 (
            .in0(N__34829),
            .in1(N__49900),
            .in2(N__54983),
            .in3(N__36587),
            .lcout(n12411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i13_LC_8_16_3.C_ON=1'b0;
    defparam buf_dds0_i13_LC_8_16_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i13_LC_8_16_3.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i13_LC_8_16_3 (
            .in0(N__49918),
            .in1(N__28116),
            .in2(N__46420),
            .in3(N__38957),
            .lcout(buf_dds0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57948),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i4_LC_8_16_4.C_ON=1'b0;
    defparam buf_dds0_i4_LC_8_16_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i4_LC_8_16_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_dds0_i4_LC_8_16_4 (
            .in0(N__38955),
            .in1(N__51183),
            .in2(N__49923),
            .in3(N__28413),
            .lcout(buf_dds0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57948),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_8_16_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_8_16_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_8_16_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_4_lut_LC_8_16_5 (
            .in0(N__48360),
            .in1(N__56360),
            .in2(N__34834),
            .in3(N__49100),
            .lcout(n20673),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i9_LC_8_16_6.C_ON=1'b0;
    defparam buf_dds0_i9_LC_8_16_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i9_LC_8_16_6.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i9_LC_8_16_6 (
            .in0(N__38956),
            .in1(N__49919),
            .in2(N__45576),
            .in3(N__28030),
            .lcout(buf_dds0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57948),
            .ce(),
            .sr(_gnd_net_));
    defparam ICE_GPMO_1_I_0_3_lut_LC_9_2_6.C_ON=1'b0;
    defparam ICE_GPMO_1_I_0_3_lut_LC_9_2_6.SEQ_MODE=4'b0000;
    defparam ICE_GPMO_1_I_0_3_lut_LC_9_2_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 ICE_GPMO_1_I_0_3_lut_LC_9_2_6 (
            .in0(N__31373),
            .in1(N__23093),
            .in2(_gnd_net_),
            .in3(N__35720),
            .lcout(IAC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_9_3_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_9_3_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i14_LC_9_3_0  (
            .in0(N__35417),
            .in1(N__23686),
            .in2(N__25948),
            .in3(N__34455),
            .lcout(cmd_rdadctmp_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57810),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i7_LC_9_3_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i7_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i7_LC_9_3_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i7_LC_9_3_1  (
            .in0(N__53199),
            .in1(N__52994),
            .in2(N__23717),
            .in3(N__23623),
            .lcout(buf_adcdata_iac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57810),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_7_i19_3_lut_LC_9_3_2.C_ON=1'b0;
    defparam mux_136_Mux_7_i19_3_lut_LC_9_3_2.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_7_i19_3_lut_LC_9_3_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_136_Mux_7_i19_3_lut_LC_9_3_2 (
            .in0(N__23675),
            .in1(N__23646),
            .in2(_gnd_net_),
            .in3(N__56359),
            .lcout(),
            .ltout(n19_adj_1625_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_7_i22_3_lut_LC_9_3_3.C_ON=1'b0;
    defparam mux_136_Mux_7_i22_3_lut_LC_9_3_3.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_7_i22_3_lut_LC_9_3_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_136_Mux_7_i22_3_lut_LC_9_3_3 (
            .in0(_gnd_net_),
            .in1(N__23622),
            .in2(N__23609),
            .in3(N__49116),
            .lcout(),
            .ltout(n22_adj_1626_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_7_i30_3_lut_LC_9_3_4.C_ON=1'b0;
    defparam mux_136_Mux_7_i30_3_lut_LC_9_3_4.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_7_i30_3_lut_LC_9_3_4.LUT_INIT=16'b1101100011011000;
    LogicCell40 mux_136_Mux_7_i30_3_lut_LC_9_3_4 (
            .in0(N__48723),
            .in1(N__23606),
            .in2(N__23594),
            .in3(_gnd_net_),
            .lcout(n30_adj_1627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i0_LC_9_3_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i0_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i0_LC_9_3_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i0_LC_9_3_7  (
            .in0(N__34654),
            .in1(N__35418),
            .in2(N__33957),
            .in3(N__26970),
            .lcout(buf_adcdata_vac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57810),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_9_4_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_9_4_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i13_LC_9_4_0  (
            .in0(N__52951),
            .in1(N__25878),
            .in2(N__28762),
            .in3(N__52073),
            .lcout(cmd_rdadctmp_13_adj_1437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57815),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i6_LC_9_4_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i6_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i6_LC_9_4_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_IAC.ADC_DATA_i6_LC_9_4_1  (
            .in0(N__53198),
            .in1(N__23767),
            .in2(N__52997),
            .in3(N__23731),
            .lcout(buf_adcdata_iac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57815),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_6_i19_3_lut_LC_9_4_2.C_ON=1'b0;
    defparam mux_136_Mux_6_i19_3_lut_LC_9_4_2.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_6_i19_3_lut_LC_9_4_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_136_Mux_6_i19_3_lut_LC_9_4_2 (
            .in0(N__23583),
            .in1(N__23564),
            .in2(_gnd_net_),
            .in3(N__56361),
            .lcout(),
            .ltout(n19_adj_1628_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_6_i22_3_lut_LC_9_4_3.C_ON=1'b0;
    defparam mux_136_Mux_6_i22_3_lut_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_6_i22_3_lut_LC_9_4_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_136_Mux_6_i22_3_lut_LC_9_4_3 (
            .in0(_gnd_net_),
            .in1(N__23766),
            .in2(N__23750),
            .in3(N__49117),
            .lcout(),
            .ltout(n22_adj_1629_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_6_i30_3_lut_LC_9_4_4.C_ON=1'b0;
    defparam mux_136_Mux_6_i30_3_lut_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_6_i30_3_lut_LC_9_4_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_136_Mux_6_i30_3_lut_LC_9_4_4 (
            .in0(_gnd_net_),
            .in1(N__23747),
            .in2(N__23735),
            .in3(N__48668),
            .lcout(n30_adj_1630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_9_4_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_9_4_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i14_LC_9_4_5  (
            .in0(N__52071),
            .in1(N__23727),
            .in2(N__25885),
            .in3(N__52953),
            .lcout(cmd_rdadctmp_14_adj_1436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57815),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_9_4_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_9_4_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i15_LC_9_4_6  (
            .in0(N__52952),
            .in1(N__23709),
            .in2(N__23732),
            .in3(N__52074),
            .lcout(cmd_rdadctmp_15_adj_1435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57815),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_9_4_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_9_4_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i16_LC_9_4_7  (
            .in0(N__52072),
            .in1(N__52105),
            .in2(N__23716),
            .in3(N__52954),
            .lcout(cmd_rdadctmp_16_adj_1434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57815),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_9_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_9_5_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i1_LC_9_5_0  (
            .in0(N__33116),
            .in1(N__26242),
            .in2(N__26180),
            .in3(N__26151),
            .lcout(cmd_rdadctmp_1_adj_1478),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_9_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_9_5_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i7_LC_9_5_1  (
            .in0(N__26001),
            .in1(N__26520),
            .in2(N__26277),
            .in3(N__33121),
            .lcout(cmd_rdadctmp_7_adj_1472),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_9_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_9_5_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i6_LC_9_5_2  (
            .in0(N__33117),
            .in1(N__26002),
            .in2(N__26036),
            .in3(N__26246),
            .lcout(cmd_rdadctmp_6_adj_1473),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_9_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_9_5_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i0_LC_9_5_3  (
            .in0(N__26241),
            .in1(N__26175),
            .in2(N__33629),
            .in3(N__33119),
            .lcout(cmd_rdadctmp_0_adj_1479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_5_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i9_LC_9_5_4  (
            .in0(N__33118),
            .in1(N__26492),
            .in2(N__26459),
            .in3(N__26250),
            .lcout(cmd_rdadctmp_9_adj_1470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_5  (
            .in0(N__26031),
            .in1(N__26065),
            .in2(N__26276),
            .in3(N__33120),
            .lcout(cmd_rdadctmp_5_adj_1474),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i12_LC_9_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i12_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i12_LC_9_5_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i12_LC_9_5_7  (
            .in0(N__33339),
            .in1(N__35614),
            .in2(N__29163),
            .in3(N__26933),
            .lcout(buf_adcdata_vdc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40121),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_0  (
            .in0(N__33109),
            .in1(N__26392),
            .in2(N__26426),
            .in3(N__26232),
            .lcout(cmd_rdadctmp_11_adj_1468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_1  (
            .in0(N__26391),
            .in1(N__26364),
            .in2(N__26274),
            .in3(N__33113),
            .lcout(cmd_rdadctmp_12_adj_1467),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_27_LC_9_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_27_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_27_LC_9_6_2 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_27_LC_9_6_2  (
            .in0(N__33108),
            .in1(N__32902),
            .in2(N__33358),
            .in3(N__33473),
            .lcout(n12875),
            .ltout(n12875_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_3 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_3  (
            .in0(N__26330),
            .in1(N__26842),
            .in2(N__23774),
            .in3(N__33114),
            .lcout(cmd_rdadctmp_14_adj_1465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_4  (
            .in0(N__33110),
            .in1(N__26236),
            .in2(N__26371),
            .in3(N__26329),
            .lcout(cmd_rdadctmp_13_adj_1466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_9_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_9_6_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i19_LC_9_6_5  (
            .in0(N__26637),
            .in1(N__26680),
            .in2(N__26275),
            .in3(N__33115),
            .lcout(cmd_rdadctmp_19_adj_1460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_6  (
            .in0(N__33111),
            .in1(N__26638),
            .in2(N__26603),
            .in3(N__26240),
            .lcout(cmd_rdadctmp_20_adj_1459),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_6_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i10_LC_9_6_7  (
            .in0(N__26421),
            .in1(N__26454),
            .in2(N__26273),
            .in3(N__33112),
            .lcout(cmd_rdadctmp_10_adj_1469),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40053),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i18_LC_9_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i18_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i18_LC_9_7_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ADC_VDC.ADC_DATA_i18_LC_9_7_0  (
            .in0(N__26879),
            .in1(N__29150),
            .in2(N__23956),
            .in3(N__33338),
            .lcout(buf_adcdata_vdc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i11_LC_9_7_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i11_LC_9_7_1  (
            .in0(N__33337),
            .in1(N__38248),
            .in2(N__29172),
            .in3(N__26948),
            .lcout(buf_adcdata_vdc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam n22214_bdd_4_lut_LC_9_7_2.C_ON=1'b0;
    defparam n22214_bdd_4_lut_LC_9_7_2.SEQ_MODE=4'b0000;
    defparam n22214_bdd_4_lut_LC_9_7_2.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22214_bdd_4_lut_LC_9_7_2 (
            .in0(N__48340),
            .in1(N__29428),
            .in2(N__23882),
            .in3(N__23891),
            .lcout(n20828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_7_3 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i15_LC_9_7_3  (
            .in0(N__26802),
            .in1(N__26843),
            .in2(N__26278),
            .in3(N__33083),
            .lcout(cmd_rdadctmp_15_adj_1464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_9_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_9_7_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i17_LC_9_7_4  (
            .in0(N__33082),
            .in1(N__26721),
            .in2(N__26768),
            .in3(N__26255),
            .lcout(cmd_rdadctmp_17_adj_1462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i8_LC_9_7_5  (
            .in0(N__26487),
            .in1(N__26525),
            .in2(N__26280),
            .in3(N__33085),
            .lcout(cmd_rdadctmp_8_adj_1471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_9_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_9_7_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i16_LC_9_7_6  (
            .in0(N__33081),
            .in1(N__26803),
            .in2(N__26767),
            .in3(N__26254),
            .lcout(cmd_rdadctmp_16_adj_1463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_9_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_9_7_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i18_LC_9_7_7  (
            .in0(N__26722),
            .in1(N__26679),
            .in2(N__26279),
            .in3(N__33084),
            .lcout(cmd_rdadctmp_18_adj_1461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40118),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i9_4_lut_LC_9_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.i9_4_lut_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i9_4_lut_LC_9_8_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \ADC_VDC.i9_4_lut_LC_9_8_1  (
            .in0(N__23858),
            .in1(N__23840),
            .in2(N__23822),
            .in3(N__23801),
            .lcout(\ADC_VDC.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18888_3_lut_LC_9_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.i18888_3_lut_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18888_3_lut_LC_9_8_2 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \ADC_VDC.i18888_3_lut_LC_9_8_2  (
            .in0(N__27022),
            .in1(N__33354),
            .in2(_gnd_net_),
            .in3(N__24011),
            .lcout(),
            .ltout(\ADC_VDC.n21145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_8_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i34_LC_9_8_3  (
            .in0(N__33123),
            .in1(N__27002),
            .in2(N__24002),
            .in3(N__32867),
            .lcout(cmd_rdadcbuf_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40088),
            .ce(N__23999),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_9_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_9_8_5 .LUT_INIT=16'b1110000010101010;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_9_8_5  (
            .in0(N__33122),
            .in1(N__32866),
            .in2(N__33371),
            .in3(N__33474),
            .lcout(\ADC_VDC.n13050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i10_LC_9_9_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i10_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i10_LC_9_9_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \RTD.READ_DATA_i10_LC_9_9_0  (
            .in0(N__24418),
            .in1(N__24233),
            .in2(N__23990),
            .in3(N__25120),
            .lcout(buf_readRTD_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43779),
            .ce(),
            .sr(_gnd_net_));
    defparam i12112_2_lut_LC_9_9_1.C_ON=1'b0;
    defparam i12112_2_lut_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam i12112_2_lut_LC_9_9_1.LUT_INIT=16'b0000000010101010;
    LogicCell40 i12112_2_lut_LC_9_9_1 (
            .in0(N__54106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54846),
            .lcout(n14522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18219_3_lut_LC_9_9_2.C_ON=1'b0;
    defparam i18219_3_lut_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam i18219_3_lut_LC_9_9_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18219_3_lut_LC_9_9_2 (
            .in0(N__23963),
            .in1(N__29029),
            .in2(_gnd_net_),
            .in3(N__56250),
            .lcout(),
            .ltout(n20833_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19484_LC_9_9_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19484_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19484_LC_9_9_3.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19484_LC_9_9_3 (
            .in0(N__25058),
            .in1(N__48309),
            .in2(N__23939),
            .in3(N__49059),
            .lcout(n22118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i14_LC_9_9_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i14_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i14_LC_9_9_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \RTD.READ_DATA_i14_LC_9_9_4  (
            .in0(N__24419),
            .in1(N__24234),
            .in2(N__23936),
            .in3(N__28885),
            .lcout(buf_readRTD_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43779),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19562_LC_9_9_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19562_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19562_LC_9_9_5.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19562_LC_9_9_5 (
            .in0(N__56249),
            .in1(N__25196),
            .in2(N__23912),
            .in3(N__48308),
            .lcout(n22214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_4_lut_LC_9_9_6 .C_ON=1'b0;
    defparam \RTD.i2_4_lut_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_4_lut_LC_9_9_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i2_4_lut_LC_9_9_6  (
            .in0(N__25103),
            .in1(N__24484),
            .in2(N__25255),
            .in3(N__24904),
            .lcout(\RTD.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i2_LC_9_10_0 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i2_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i2_LC_9_10_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i2_LC_9_10_0  (
            .in0(N__24103),
            .in1(N__24125),
            .in2(N__25095),
            .in3(N__24905),
            .lcout(\RTD.cfg_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43736),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i0_LC_9_10_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i0_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i0_LC_9_10_1 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i0_LC_9_10_1  (
            .in0(N__24449),
            .in1(N__24892),
            .in2(N__41251),
            .in3(N__24227),
            .lcout(buf_readRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43736),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_9_10_2 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_9_10_2 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \RTD.i1_2_lut_3_lut_4_lut_LC_9_10_2  (
            .in0(N__24796),
            .in1(N__24448),
            .in2(N__25048),
            .in3(N__24674),
            .lcout(\RTD.n14717 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_7_i16_3_lut_LC_9_10_3.C_ON=1'b0;
    defparam mux_134_Mux_7_i16_3_lut_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i16_3_lut_LC_9_10_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_134_Mux_7_i16_3_lut_LC_9_10_3 (
            .in0(N__25276),
            .in1(N__28064),
            .in2(_gnd_net_),
            .in3(N__56180),
            .lcout(n16_adj_1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i4_LC_9_10_4 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i4_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i4_LC_9_10_4 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i4_LC_9_10_4  (
            .in0(N__24104),
            .in1(N__24126),
            .in2(N__25248),
            .in3(N__24485),
            .lcout(\RTD.cfg_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43736),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i6_LC_9_10_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i6_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i6_LC_9_10_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i6_LC_9_10_5  (
            .in0(N__24450),
            .in1(N__38044),
            .in2(N__24266),
            .in3(N__24228),
            .lcout(buf_readRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43736),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i7_LC_9_10_7 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i7_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i7_LC_9_10_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.cfg_buf_i7_LC_9_10_7  (
            .in0(N__24127),
            .in1(N__24105),
            .in2(N__24026),
            .in3(N__24064),
            .lcout(\RTD.cfg_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43736),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i3_LC_9_11_0.C_ON=1'b0;
    defparam comm_cmd_i3_LC_9_11_0.SEQ_MODE=4'b1000;
    defparam comm_cmd_i3_LC_9_11_0.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i3_LC_9_11_0 (
            .in0(N__40802),
            .in1(N__32053),
            .in2(N__48620),
            .in3(N__32099),
            .lcout(comm_cmd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57869),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i3_LC_9_11_2.C_ON=1'b0;
    defparam buf_cfgRTD_i3_LC_9_11_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i3_LC_9_11_2.LUT_INIT=16'b0011101100001000;
    LogicCell40 buf_cfgRTD_i3_LC_9_11_2 (
            .in0(N__44307),
            .in1(N__29001),
            .in2(N__49917),
            .in3(N__25187),
            .lcout(buf_cfgRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57869),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i8_LC_9_11_3  (
            .in0(N__52089),
            .in1(N__25163),
            .in2(N__29394),
            .in3(N__52911),
            .lcout(cmd_rdadctmp_8_adj_1442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57869),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i2_LC_9_11_4.C_ON=1'b0;
    defparam buf_cfgRTD_i2_LC_9_11_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i2_LC_9_11_4.LUT_INIT=16'b0010111000100010;
    LogicCell40 buf_cfgRTD_i2_LC_9_11_4 (
            .in0(N__25085),
            .in1(N__29000),
            .in2(N__49916),
            .in3(N__43009),
            .lcout(buf_cfgRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57869),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19542_LC_9_11_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19542_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19542_LC_9_11_5.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19542_LC_9_11_5 (
            .in0(N__56263),
            .in1(N__27473),
            .in2(N__25142),
            .in3(N__48299),
            .lcout(n22184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18220_3_lut_LC_9_11_6.C_ON=1'b0;
    defparam i18220_3_lut_LC_9_11_6.SEQ_MODE=4'b0000;
    defparam i18220_3_lut_LC_9_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18220_3_lut_LC_9_11_6 (
            .in0(N__25121),
            .in1(N__25084),
            .in2(_gnd_net_),
            .in3(N__56264),
            .lcout(n20834),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_adj_19_LC_9_11_7 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_adj_19_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_adj_19_LC_9_11_7 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \RTD.i1_2_lut_3_lut_adj_19_LC_9_11_7  (
            .in0(N__33844),
            .in1(N__25047),
            .in2(_gnd_net_),
            .in3(N__31702),
            .lcout(\RTD.n20656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_216_LC_9_12_0.C_ON=1'b0;
    defparam i1_4_lut_adj_216_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_216_LC_9_12_0.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_216_LC_9_12_0 (
            .in0(N__46609),
            .in1(N__54922),
            .in2(N__49895),
            .in3(N__34830),
            .lcout(n12397),
            .ltout(n12397_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i7_LC_9_12_1.C_ON=1'b0;
    defparam buf_device_acadc_i7_LC_9_12_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i7_LC_9_12_1.LUT_INIT=16'b0010111100100000;
    LogicCell40 buf_device_acadc_i7_LC_9_12_1 (
            .in0(N__43161),
            .in1(N__49839),
            .in2(N__24917),
            .in3(N__36843),
            .lcout(VAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57882),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_251_LC_9_12_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_251_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_251_LC_9_12_2.LUT_INIT=16'b1111111111011101;
    LogicCell40 i1_2_lut_3_lut_adj_251_LC_9_12_2 (
            .in0(N__27672),
            .in1(N__27255),
            .in2(_gnd_net_),
            .in3(N__27270),
            .lcout(n20646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22184_bdd_4_lut_LC_9_12_4.C_ON=1'b0;
    defparam n22184_bdd_4_lut_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam n22184_bdd_4_lut_LC_9_12_4.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22184_bdd_4_lut_LC_9_12_4 (
            .in0(N__48344),
            .in1(N__25483),
            .in2(N__25448),
            .in3(N__25424),
            .lcout(n20849),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19552_LC_9_12_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19552_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19552_LC_9_12_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19552_LC_9_12_5 (
            .in0(N__25228),
            .in1(N__48342),
            .in2(N__25418),
            .in3(N__56281),
            .lcout(n22202),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i1_LC_9_12_6.C_ON=1'b0;
    defparam buf_cfgRTD_i1_LC_9_12_6.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i1_LC_9_12_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i1_LC_9_12_6 (
            .in0(N__49838),
            .in1(N__28996),
            .in2(N__45581),
            .in3(N__27596),
            .lcout(buf_cfgRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57882),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19395_LC_9_12_7.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19395_LC_9_12_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19395_LC_9_12_7.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19395_LC_9_12_7 (
            .in0(N__25340),
            .in1(N__48343),
            .in2(N__25385),
            .in3(N__56282),
            .lcout(n22016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i0_LC_9_13_0.C_ON=1'b0;
    defparam buf_cfgRTD_i0_LC_9_13_0.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i0_LC_9_13_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i0_LC_9_13_0 (
            .in0(N__44467),
            .in1(N__28994),
            .in2(_gnd_net_),
            .in3(N__25332),
            .lcout(buf_cfgRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57895),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_13_2 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_13_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i19_LC_9_13_2  (
            .in0(N__53166),
            .in1(N__52915),
            .in2(N__25313),
            .in3(N__40893),
            .lcout(buf_adcdata_iac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57895),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i15_LC_9_13_3.C_ON=1'b0;
    defparam buf_dds1_i15_LC_9_13_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i15_LC_9_13_3.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i15_LC_9_13_3 (
            .in0(N__25275),
            .in1(N__38574),
            .in2(N__46066),
            .in3(N__38479),
            .lcout(buf_dds1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57895),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i4_LC_9_13_4.C_ON=1'b0;
    defparam buf_cfgRTD_i4_LC_9_13_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i4_LC_9_13_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i4_LC_9_13_4 (
            .in0(N__49921),
            .in1(N__28995),
            .in2(N__44174),
            .in3(N__25229),
            .lcout(buf_cfgRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57895),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i3_LC_9_13_5.C_ON=1'b0;
    defparam buf_device_acadc_i3_LC_9_13_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i3_LC_9_13_5.LUT_INIT=16'b0010001011100010;
    LogicCell40 buf_device_acadc_i3_LC_9_13_5 (
            .in0(N__27399),
            .in1(N__41375),
            .in2(N__43010),
            .in3(N__49922),
            .lcout(IAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57895),
            .ce(),
            .sr(_gnd_net_));
    defparam n22106_bdd_4_lut_LC_9_13_6.C_ON=1'b0;
    defparam n22106_bdd_4_lut_LC_9_13_6.SEQ_MODE=4'b0000;
    defparam n22106_bdd_4_lut_LC_9_13_6.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22106_bdd_4_lut_LC_9_13_6 (
            .in0(N__25571),
            .in1(N__25505),
            .in2(N__25565),
            .in3(N__48538),
            .lcout(n22109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19405_LC_9_14_1.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19405_LC_9_14_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19405_LC_9_14_1.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19405_LC_9_14_1 (
            .in0(N__48297),
            .in1(N__27703),
            .in2(N__25546),
            .in3(N__56301),
            .lcout(n22022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18262_4_lut_LC_9_14_3.C_ON=1'b0;
    defparam i18262_4_lut_LC_9_14_3.SEQ_MODE=4'b0000;
    defparam i18262_4_lut_LC_9_14_3.LUT_INIT=16'b0101000010001000;
    LogicCell40 i18262_4_lut_LC_9_14_3 (
            .in0(N__48298),
            .in1(N__25523),
            .in2(N__32153),
            .in3(N__56302),
            .lcout(),
            .ltout(n20876_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19479_LC_9_14_4.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19479_LC_9_14_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19479_LC_9_14_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19479_LC_9_14_4 (
            .in0(N__25499),
            .in1(N__48574),
            .in2(N__25508),
            .in3(N__49058),
            .lcout(n22106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i12_LC_9_14_5.C_ON=1'b0;
    defparam buf_dds1_i12_LC_9_14_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i12_LC_9_14_5.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i12_LC_9_14_5 (
            .in0(N__40294),
            .in1(N__38573),
            .in2(N__44168),
            .in3(N__38472),
            .lcout(buf_dds1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57911),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_1_i16_3_lut_LC_9_14_6.C_ON=1'b0;
    defparam mux_135_Mux_1_i16_3_lut_LC_9_14_6.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_1_i16_3_lut_LC_9_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_135_Mux_1_i16_3_lut_LC_9_14_6 (
            .in0(N__56303),
            .in1(N__38399),
            .in2(_gnd_net_),
            .in3(N__28339),
            .lcout(n16_adj_1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18261_4_lut_LC_9_14_7.C_ON=1'b0;
    defparam i18261_4_lut_LC_9_14_7.SEQ_MODE=4'b0000;
    defparam i18261_4_lut_LC_9_14_7.LUT_INIT=16'b0111001001010000;
    LogicCell40 i18261_4_lut_LC_9_14_7 (
            .in0(N__48296),
            .in1(N__56300),
            .in2(N__30923),
            .in3(N__47555),
            .lcout(n20875),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i7_LC_9_15_0.C_ON=1'b0;
    defparam data_index_i7_LC_9_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i7_LC_9_15_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i7_LC_9_15_0 (
            .in0(N__27845),
            .in1(N__54949),
            .in2(N__49823),
            .in3(N__27836),
            .lcout(data_index_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57925),
            .ce(),
            .sr(_gnd_net_));
    defparam n22022_bdd_4_lut_LC_9_15_3.C_ON=1'b0;
    defparam n22022_bdd_4_lut_LC_9_15_3.SEQ_MODE=4'b0000;
    defparam n22022_bdd_4_lut_LC_9_15_3.LUT_INIT=16'b1100101111001000;
    LogicCell40 n22022_bdd_4_lut_LC_9_15_3 (
            .in0(N__25608),
            .in1(N__25493),
            .in2(N__48424),
            .in3(N__28023),
            .lcout(n22025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i4_LC_9_15_4.C_ON=1'b0;
    defparam buf_dds1_i4_LC_9_15_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i4_LC_9_15_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i4_LC_9_15_4 (
            .in0(N__25744),
            .in1(N__38562),
            .in2(N__51188),
            .in3(N__38455),
            .lcout(buf_dds1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57925),
            .ce(),
            .sr(_gnd_net_));
    defparam i6394_3_lut_LC_9_15_5.C_ON=1'b0;
    defparam i6394_3_lut_LC_9_15_5.SEQ_MODE=4'b0000;
    defparam i6394_3_lut_LC_9_15_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6394_3_lut_LC_9_15_5 (
            .in0(N__41498),
            .in1(N__27920),
            .in2(_gnd_net_),
            .in3(N__41749),
            .lcout(n8_adj_1555),
            .ltout(n8_adj_1555_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_8_i15_4_lut_LC_9_15_6.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_8_i15_4_lut_LC_9_15_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_8_i15_4_lut_LC_9_15_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_365_Mux_8_i15_4_lut_LC_9_15_6 (
            .in0(N__49734),
            .in1(N__54948),
            .in2(N__25724),
            .in3(N__27898),
            .lcout(data_index_9_N_216_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i8_LC_9_15_7.C_ON=1'b0;
    defparam data_index_i8_LC_9_15_7.SEQ_MODE=4'b1000;
    defparam data_index_i8_LC_9_15_7.LUT_INIT=16'b0011101000001010;
    LogicCell40 data_index_i8_LC_9_15_7 (
            .in0(N__27899),
            .in1(N__49735),
            .in2(N__54977),
            .in3(N__25625),
            .lcout(data_index_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57925),
            .ce(),
            .sr(_gnd_net_));
    defparam n22040_bdd_4_lut_LC_9_16_0.C_ON=1'b0;
    defparam n22040_bdd_4_lut_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam n22040_bdd_4_lut_LC_9_16_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22040_bdd_4_lut_LC_9_16_0 (
            .in0(N__25587),
            .in1(N__25619),
            .in2(N__28372),
            .in3(N__48377),
            .lcout(n22043),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i10_LC_9_16_1.C_ON=1'b0;
    defparam buf_dds1_i10_LC_9_16_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i10_LC_9_16_1.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i10_LC_9_16_1 (
            .in0(N__25802),
            .in1(N__38557),
            .in2(N__43004),
            .in3(N__38448),
            .lcout(buf_dds1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57938),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i9_LC_9_16_2.C_ON=1'b0;
    defparam buf_dds1_i9_LC_9_16_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i9_LC_9_16_2.LUT_INIT=16'b1010000010001000;
    LogicCell40 buf_dds1_i9_LC_9_16_2 (
            .in0(N__38450),
            .in1(N__25610),
            .in2(N__45577),
            .in3(N__38563),
            .lcout(buf_dds1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57938),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i8_LC_9_16_3.C_ON=1'b0;
    defparam buf_dds1_i8_LC_9_16_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i8_LC_9_16_3.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i8_LC_9_16_3 (
            .in0(N__25591),
            .in1(N__38558),
            .in2(N__41510),
            .in3(N__38449),
            .lcout(buf_dds1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57938),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i1_LC_9_16_4.C_ON=1'b0;
    defparam buf_dds0_i1_LC_9_16_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i1_LC_9_16_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i1_LC_9_16_4 (
            .in0(N__49899),
            .in1(N__38932),
            .in2(N__45467),
            .in3(N__28335),
            .lcout(buf_dds0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57938),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i15_LC_9_16_5.C_ON=1'b0;
    defparam buf_dds0_i15_LC_9_16_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i15_LC_9_16_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i15_LC_9_16_5 (
            .in0(N__28060),
            .in1(N__49897),
            .in2(N__46058),
            .in3(N__38935),
            .lcout(buf_dds0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57938),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_213_LC_9_16_6.C_ON=1'b0;
    defparam i1_3_lut_adj_213_LC_9_16_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_213_LC_9_16_6.LUT_INIT=16'b1011101100000000;
    LogicCell40 i1_3_lut_adj_213_LC_9_16_6 (
            .in0(N__49896),
            .in1(N__25781),
            .in2(_gnd_net_),
            .in3(N__54963),
            .lcout(n12383),
            .ltout(n12383_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i8_LC_9_16_7.C_ON=1'b0;
    defparam buf_dds0_i8_LC_9_16_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i8_LC_9_16_7.LUT_INIT=16'b0010111100100000;
    LogicCell40 buf_dds0_i8_LC_9_16_7 (
            .in0(N__41506),
            .in1(N__49898),
            .in2(N__25805),
            .in3(N__28368),
            .lcout(buf_dds0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57938),
            .ce(),
            .sr(_gnd_net_));
    defparam i18210_3_lut_LC_9_17_2.C_ON=1'b0;
    defparam i18210_3_lut_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam i18210_3_lut_LC_9_17_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18210_3_lut_LC_9_17_2 (
            .in0(N__25797),
            .in1(N__28143),
            .in2(_gnd_net_),
            .in3(N__56339),
            .lcout(n20824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i2_LC_9_17_4.C_ON=1'b0;
    defparam buf_dds0_i2_LC_9_17_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i2_LC_9_17_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i2_LC_9_17_4 (
            .in0(N__38933),
            .in1(N__49914),
            .in2(N__47150),
            .in3(N__28440),
            .lcout(buf_dds0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57949),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i10_LC_9_17_5.C_ON=1'b0;
    defparam buf_dds0_i10_LC_9_17_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i10_LC_9_17_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i10_LC_9_17_5 (
            .in0(N__28144),
            .in1(N__49908),
            .in2(N__43003),
            .in3(N__38934),
            .lcout(buf_dds0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57949),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_253_LC_9_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_253_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_253_LC_9_17_6.LUT_INIT=16'b1011101100001011;
    LogicCell40 i1_4_lut_adj_253_LC_9_17_6 (
            .in0(N__51589),
            .in1(N__25780),
            .in2(N__49924),
            .in3(N__54964),
            .lcout(),
            .ltout(n11412_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds0_314_LC_9_17_7.C_ON=1'b0;
    defparam trig_dds0_314_LC_9_17_7.SEQ_MODE=4'b1000;
    defparam trig_dds0_314_LC_9_17_7.LUT_INIT=16'b0000110010101100;
    LogicCell40 trig_dds0_314_LC_9_17_7 (
            .in0(N__54965),
            .in1(N__44789),
            .in2(N__25769),
            .in3(N__49920),
            .lcout(trig_dds0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57949),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_I_0_1_lut_LC_9_20_2.C_ON=1'b0;
    defparam acadc_rst_I_0_1_lut_LC_9_20_2.SEQ_MODE=4'b0000;
    defparam acadc_rst_I_0_1_lut_LC_9_20_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 acadc_rst_I_0_1_lut_LC_9_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36359),
            .lcout(AC_ADC_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_10_2_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_10_2_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_10_2_2 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i8_LC_10_2_2  (
            .in0(N__25901),
            .in1(N__34424),
            .in2(N__26971),
            .in3(N__35421),
            .lcout(cmd_rdadctmp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57804),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_10_3_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_10_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_10_3_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i13_LC_10_3_0  (
            .in0(N__25944),
            .in1(N__34456),
            .in2(N__25979),
            .in3(N__35420),
            .lcout(cmd_rdadctmp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57807),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_10_3_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_10_3_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_10_3_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i7_LC_10_3_3  (
            .in0(N__35419),
            .in1(N__25900),
            .in2(N__34460),
            .in3(N__25922),
            .lcout(cmd_rdadctmp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57807),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i2_LC_10_3_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i2_LC_10_3_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i2_LC_10_3_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i2_LC_10_3_4  (
            .in0(N__53206),
            .in1(N__52993),
            .in2(N__28676),
            .in3(N__28585),
            .lcout(buf_adcdata_iac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57807),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i5_LC_10_3_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i5_LC_10_3_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i5_LC_10_3_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i5_LC_10_3_5  (
            .in0(N__52992),
            .in1(N__53207),
            .in2(N__25889),
            .in3(N__25860),
            .lcout(buf_adcdata_iac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57807),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_5_i30_3_lut_LC_10_3_7.C_ON=1'b0;
    defparam mux_136_Mux_5_i30_3_lut_LC_10_3_7.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_5_i30_3_lut_LC_10_3_7.LUT_INIT=16'b1010110010101100;
    LogicCell40 mux_136_Mux_5_i30_3_lut_LC_10_3_7 (
            .in0(N__25841),
            .in1(N__25829),
            .in2(N__48741),
            .in3(_gnd_net_),
            .lcout(n30_adj_1634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_10_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_10_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_10_4_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i2_LC_10_4_0  (
            .in0(N__33100),
            .in1(N__26121),
            .in2(N__26291),
            .in3(N__26152),
            .lcout(cmd_rdadctmp_2_adj_1477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40048),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_10_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_10_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_10_4_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i22_LC_10_4_1  (
            .in0(N__26569),
            .in1(N__31782),
            .in2(N__33127),
            .in3(N__26284),
            .lcout(cmd_rdadctmp_22_adj_1457),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40048),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19104_2_lut_LC_10_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i19104_2_lut_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19104_2_lut_LC_10_4_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ADC_VDC.i19104_2_lut_LC_10_4_3  (
            .in0(_gnd_net_),
            .in1(N__33301),
            .in2(_gnd_net_),
            .in3(N__33098),
            .lcout(\ADC_VDC.n21718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_10_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_10_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_10_4_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i21_LC_10_4_4  (
            .in0(N__33099),
            .in1(N__26568),
            .in2(N__26290),
            .in3(N__26602),
            .lcout(cmd_rdadctmp_21_adj_1458),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40048),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_10_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_10_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_10_4_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i4_LC_10_4_6  (
            .in0(N__26289),
            .in1(N__33101),
            .in2(N__26096),
            .in3(N__26064),
            .lcout(cmd_rdadctmp_4_adj_1475),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40048),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_10_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_10_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_10_4_7 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i3_LC_10_4_7  (
            .in0(N__26122),
            .in1(N__26091),
            .in2(N__33128),
            .in3(N__26288),
            .lcout(cmd_rdadctmp_3_adj_1476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40048),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_10_5_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_10_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_10_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i0_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__26159),
            .in2(N__26179),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.cmd_rdadcbuf_0 ),
            .ltout(),
            .carryin(bfn_10_5_0_),
            .carryout(\ADC_VDC.n19422 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_10_5_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_10_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i1_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__26132),
            .in2(N__26153),
            .in3(N__26126),
            .lcout(\ADC_VDC.cmd_rdadcbuf_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19422 ),
            .carryout(\ADC_VDC.n19423 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_10_5_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_10_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i2_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__26105),
            .in2(N__26123),
            .in3(N__26099),
            .lcout(\ADC_VDC.cmd_rdadcbuf_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19423 ),
            .carryout(\ADC_VDC.n19424 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_10_5_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_10_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i3_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(N__26075),
            .in2(N__26095),
            .in3(N__26069),
            .lcout(\ADC_VDC.cmd_rdadcbuf_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19424 ),
            .carryout(\ADC_VDC.n19425 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_10_5_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_10_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_10_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i4_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(N__26045),
            .in2(N__26066),
            .in3(N__26039),
            .lcout(\ADC_VDC.cmd_rdadcbuf_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19425 ),
            .carryout(\ADC_VDC.n19426 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_10_5_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_10_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i5_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__26012),
            .in2(N__26035),
            .in3(N__26006),
            .lcout(\ADC_VDC.cmd_rdadcbuf_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19426 ),
            .carryout(\ADC_VDC.n19427 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_10_5_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_10_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i6_LC_10_5_6  (
            .in0(_gnd_net_),
            .in1(N__25985),
            .in2(N__26003),
            .in3(N__26528),
            .lcout(\ADC_VDC.cmd_rdadcbuf_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19427 ),
            .carryout(\ADC_VDC.n19428 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_10_5_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_10_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i7_LC_10_5_7  (
            .in0(_gnd_net_),
            .in1(N__26501),
            .in2(N__26524),
            .in3(N__26495),
            .lcout(\ADC_VDC.cmd_rdadcbuf_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19428 ),
            .carryout(\ADC_VDC.n19429 ),
            .clk(N__40034),
            .ce(N__27190),
            .sr(N__27107));
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_10_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_10_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i8_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__26468),
            .in2(N__26491),
            .in3(N__26462),
            .lcout(\ADC_VDC.cmd_rdadcbuf_8 ),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\ADC_VDC.n19430 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_10_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_10_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i9_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__26435),
            .in2(N__26458),
            .in3(N__26429),
            .lcout(\ADC_VDC.cmd_rdadcbuf_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19430 ),
            .carryout(\ADC_VDC.n19431 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_10_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_10_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i10_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__26402),
            .in2(N__26425),
            .in3(N__26396),
            .lcout(\ADC_VDC.cmd_rdadcbuf_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19431 ),
            .carryout(\ADC_VDC.n19432 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_10_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_10_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i11_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__29200),
            .in2(N__26393),
            .in3(N__26375),
            .lcout(cmd_rdadcbuf_11),
            .ltout(),
            .carryin(\ADC_VDC.n19432 ),
            .carryout(\ADC_VDC.n19433 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_10_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_10_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i12_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__26344),
            .in2(N__26372),
            .in3(N__26333),
            .lcout(cmd_rdadcbuf_12),
            .ltout(),
            .carryin(\ADC_VDC.n19433 ),
            .carryout(\ADC_VDC.n19434 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_10_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_10_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i13_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__26328),
            .in2(N__26311),
            .in3(N__26294),
            .lcout(cmd_rdadcbuf_13),
            .ltout(),
            .carryin(\ADC_VDC.n19434 ),
            .carryout(\ADC_VDC.n19435 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_10_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_10_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i14_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__26841),
            .in2(N__26824),
            .in3(N__26807),
            .lcout(cmd_rdadcbuf_14),
            .ltout(),
            .carryin(\ADC_VDC.n19435 ),
            .carryout(\ADC_VDC.n19436 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_10_6_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_10_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i15_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__26782),
            .in2(N__26804),
            .in3(N__26771),
            .lcout(cmd_rdadcbuf_15),
            .ltout(),
            .carryin(\ADC_VDC.n19436 ),
            .carryout(\ADC_VDC.n19437 ),
            .clk(N__40049),
            .ce(N__27183),
            .sr(N__27106));
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_10_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_10_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i16_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__26737),
            .in2(N__26766),
            .in3(N__26726),
            .lcout(cmd_rdadcbuf_16),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\ADC_VDC.n19438 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_10_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_10_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i17_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__26695),
            .in2(N__26723),
            .in3(N__26684),
            .lcout(cmd_rdadcbuf_17),
            .ltout(),
            .carryin(\ADC_VDC.n19438 ),
            .carryout(\ADC_VDC.n19439 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_10_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_10_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i18_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__26653),
            .in2(N__26681),
            .in3(N__26642),
            .lcout(cmd_rdadcbuf_18),
            .ltout(),
            .carryin(\ADC_VDC.n19439 ),
            .carryout(\ADC_VDC.n19440 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_10_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_10_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i19_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__26617),
            .in2(N__26639),
            .in3(N__26606),
            .lcout(cmd_rdadcbuf_19),
            .ltout(),
            .carryin(\ADC_VDC.n19440 ),
            .carryout(\ADC_VDC.n19441 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_10_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_10_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i20_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__29044),
            .in2(N__26601),
            .in3(N__26576),
            .lcout(cmd_rdadcbuf_20),
            .ltout(),
            .carryin(\ADC_VDC.n19441 ),
            .carryout(\ADC_VDC.n19442 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_10_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_10_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i21_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__26542),
            .in2(N__26573),
            .in3(N__26531),
            .lcout(cmd_rdadcbuf_21),
            .ltout(),
            .carryin(\ADC_VDC.n19442 ),
            .carryout(\ADC_VDC.n19443 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_10_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_10_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i22_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__26947),
            .in2(N__31789),
            .in3(N__26936),
            .lcout(cmd_rdadcbuf_22),
            .ltout(),
            .carryin(\ADC_VDC.n19443 ),
            .carryout(\ADC_VDC.n19444 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_10_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_10_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i23_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(N__26929),
            .in2(N__31751),
            .in3(N__26918),
            .lcout(cmd_rdadcbuf_23),
            .ltout(),
            .carryin(\ADC_VDC.n19444 ),
            .carryout(\ADC_VDC.n19445 ),
            .clk(N__40117),
            .ce(N__27159),
            .sr(N__27105));
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_10_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_10_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i24_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__28846),
            .in2(_gnd_net_),
            .in3(N__26915),
            .lcout(cmd_rdadcbuf_24),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\ADC_VDC.n19446 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_10_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_10_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i25_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__28858),
            .in2(_gnd_net_),
            .in3(N__26912),
            .lcout(cmd_rdadcbuf_25),
            .ltout(),
            .carryin(\ADC_VDC.n19446 ),
            .carryout(\ADC_VDC.n19447 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_10_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_10_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i26_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__28870),
            .in2(_gnd_net_),
            .in3(N__26909),
            .lcout(cmd_rdadcbuf_26),
            .ltout(),
            .carryin(\ADC_VDC.n19447 ),
            .carryout(\ADC_VDC.n19448 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_10_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_10_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i27_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__29215),
            .in2(_gnd_net_),
            .in3(N__26906),
            .lcout(cmd_rdadcbuf_27),
            .ltout(),
            .carryin(\ADC_VDC.n19448 ),
            .carryout(\ADC_VDC.n19449 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_10_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_10_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i28_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__26893),
            .in2(_gnd_net_),
            .in3(N__26882),
            .lcout(cmd_rdadcbuf_28),
            .ltout(),
            .carryin(\ADC_VDC.n19449 ),
            .carryout(\ADC_VDC.n19450 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_10_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_10_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i29_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__26875),
            .in2(_gnd_net_),
            .in3(N__26864),
            .lcout(cmd_rdadcbuf_29),
            .ltout(),
            .carryin(\ADC_VDC.n19450 ),
            .carryout(\ADC_VDC.n19451 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_10_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_10_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i30_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__26857),
            .in2(_gnd_net_),
            .in3(N__26846),
            .lcout(cmd_rdadcbuf_30),
            .ltout(),
            .carryin(\ADC_VDC.n19451 ),
            .carryout(\ADC_VDC.n19452 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_10_8_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_10_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i31_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__27232),
            .in2(_gnd_net_),
            .in3(N__27221),
            .lcout(cmd_rdadcbuf_31),
            .ltout(),
            .carryin(\ADC_VDC.n19452 ),
            .carryout(\ADC_VDC.n19453 ),
            .clk(N__40116),
            .ce(N__27172),
            .sr(N__27099));
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_10_9_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_10_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i32_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__27208),
            .in2(_gnd_net_),
            .in3(N__27197),
            .lcout(cmd_rdadcbuf_32),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\ADC_VDC.n19454 ),
            .clk(N__40119),
            .ce(N__27191),
            .sr(N__27104));
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_10_9_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i33_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__29188),
            .in2(_gnd_net_),
            .in3(N__27194),
            .lcout(cmd_rdadcbuf_33),
            .ltout(),
            .carryin(\ADC_VDC.n19454 ),
            .carryout(\ADC_VDC.n19455 ),
            .clk(N__40119),
            .ce(N__27191),
            .sr(N__27104));
    defparam \ADC_VDC.add_23_36_lut_LC_10_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.add_23_36_lut_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.add_23_36_lut_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.add_23_36_lut_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__27021),
            .in2(_gnd_net_),
            .in3(N__27005),
            .lcout(\ADC_VDC.cmd_rdadcbuf_35_N_1139_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_376_i9_2_lut_3_lut_LC_10_10_0.C_ON=1'b0;
    defparam comm_cmd_6__I_0_376_i9_2_lut_3_lut_LC_10_10_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_376_i9_2_lut_3_lut_LC_10_10_0.LUT_INIT=16'b1111111111101110;
    LogicCell40 comm_cmd_6__I_0_376_i9_2_lut_3_lut_LC_10_10_0 (
            .in0(N__48171),
            .in1(N__56182),
            .in2(_gnd_net_),
            .in3(N__48952),
            .lcout(n9_adj_1416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_10_10_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_10_10_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i10_LC_10_10_1  (
            .in0(N__34761),
            .in1(N__34380),
            .in2(N__28531),
            .in3(N__35345),
            .lcout(cmd_rdadctmp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57850),
            .ce(),
            .sr(_gnd_net_));
    defparam n22118_bdd_4_lut_LC_10_10_3.C_ON=1'b0;
    defparam n22118_bdd_4_lut_LC_10_10_3.SEQ_MODE=4'b0000;
    defparam n22118_bdd_4_lut_LC_10_10_3.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22118_bdd_4_lut_LC_10_10_3 (
            .in0(N__48953),
            .in1(N__27380),
            .in2(N__26996),
            .in3(N__26978),
            .lcout(n22121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_194_i9_2_lut_3_lut_LC_10_10_4.C_ON=1'b0;
    defparam equal_194_i9_2_lut_3_lut_LC_10_10_4.SEQ_MODE=4'b0000;
    defparam equal_194_i9_2_lut_3_lut_LC_10_10_4.LUT_INIT=16'b1111111111011101;
    LogicCell40 equal_194_i9_2_lut_3_lut_LC_10_10_4 (
            .in0(N__48170),
            .in1(N__56181),
            .in2(_gnd_net_),
            .in3(N__48951),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_10_10_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_10_10_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i9_LC_10_10_5  (
            .in0(N__26972),
            .in1(N__34382),
            .in2(N__34765),
            .in3(N__35347),
            .lcout(cmd_rdadctmp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57850),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i5_LC_10_10_6.C_ON=1'b0;
    defparam buf_cfgRTD_i5_LC_10_10_6.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i5_LC_10_10_6.LUT_INIT=16'b0111010000110000;
    LogicCell40 buf_cfgRTD_i5_LC_10_10_6 (
            .in0(N__49828),
            .in1(N__29006),
            .in2(N__27483),
            .in3(N__46405),
            .lcout(buf_cfgRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57850),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_10_10_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_10_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_10_10_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i25_LC_10_10_7  (
            .in0(N__29239),
            .in1(N__34381),
            .in2(N__34482),
            .in3(N__35346),
            .lcout(cmd_rdadctmp_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57850),
            .ce(),
            .sr(_gnd_net_));
    defparam i18211_3_lut_LC_10_11_0.C_ON=1'b0;
    defparam i18211_3_lut_LC_10_11_0.SEQ_MODE=4'b0000;
    defparam i18211_3_lut_LC_10_11_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18211_3_lut_LC_10_11_0 (
            .in0(N__56166),
            .in1(N__27451),
            .in2(_gnd_net_),
            .in3(N__27403),
            .lcout(n20825),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i14_LC_10_11_1.C_ON=1'b0;
    defparam buf_dds0_i14_LC_10_11_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i14_LC_10_11_1.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_dds0_i14_LC_10_11_1 (
            .in0(N__38964),
            .in1(N__43153),
            .in2(N__49825),
            .in3(N__36909),
            .lcout(buf_dds0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57860),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_0_i16_3_lut_LC_10_11_2.C_ON=1'b0;
    defparam mux_135_Mux_0_i16_3_lut_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_0_i16_3_lut_LC_10_11_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_135_Mux_0_i16_3_lut_LC_10_11_2 (
            .in0(N__56167),
            .in1(_gnd_net_),
            .in2(N__27538),
            .in3(N__31189),
            .lcout(n16_adj_1488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_0_i15_4_lut_LC_10_11_3.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_0_i15_4_lut_LC_10_11_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_0_i15_4_lut_LC_10_11_3.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_365_Mux_0_i15_4_lut_LC_10_11_3 (
            .in0(N__54923),
            .in1(N__31013),
            .in2(N__49824),
            .in3(N__30896),
            .lcout(data_index_9_N_216_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15049_2_lut_3_lut_LC_10_11_4.C_ON=1'b0;
    defparam i15049_2_lut_3_lut_LC_10_11_4.SEQ_MODE=4'b0000;
    defparam i15049_2_lut_3_lut_LC_10_11_4.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15049_2_lut_3_lut_LC_10_11_4 (
            .in0(N__27673),
            .in1(N__27256),
            .in2(_gnd_net_),
            .in3(N__27271),
            .lcout(comm_state_3_N_436_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i5_LC_10_11_6.C_ON=1'b0;
    defparam comm_cmd_i5_LC_10_11_6.SEQ_MODE=4'b1000;
    defparam comm_cmd_i5_LC_10_11_6.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i5_LC_10_11_6 (
            .in0(N__32045),
            .in1(N__32101),
            .in2(N__51059),
            .in3(N__27272),
            .lcout(comm_cmd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57860),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i6_LC_10_11_7.C_ON=1'b0;
    defparam comm_cmd_i6_LC_10_11_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i6_LC_10_11_7.LUT_INIT=16'b1010000011001100;
    LogicCell40 comm_cmd_i6_LC_10_11_7 (
            .in0(N__40247),
            .in1(N__27257),
            .in2(N__32116),
            .in3(N__32046),
            .lcout(comm_cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57860),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i2_LC_10_12_1.C_ON=1'b0;
    defparam buf_device_acadc_i2_LC_10_12_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i2_LC_10_12_1.LUT_INIT=16'b0010111100100000;
    LogicCell40 buf_device_acadc_i2_LC_10_12_1 (
            .in0(N__45544),
            .in1(N__49749),
            .in2(N__41382),
            .in3(N__27693),
            .lcout(IAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57870),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i4_LC_10_12_2.C_ON=1'b0;
    defparam comm_cmd_i4_LC_10_12_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i4_LC_10_12_2.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i4_LC_10_12_2 (
            .in0(N__32122),
            .in1(N__32054),
            .in2(N__40661),
            .in3(N__27674),
            .lcout(comm_cmd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57870),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i3_LC_10_12_4.C_ON=1'b0;
    defparam buf_dds1_i3_LC_10_12_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i3_LC_10_12_4.LUT_INIT=16'b1110001011101110;
    LogicCell40 buf_dds1_i3_LC_10_12_4 (
            .in0(N__27648),
            .in1(N__38578),
            .in2(N__47841),
            .in3(N__54946),
            .lcout(buf_dds1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57870),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_LC_10_12_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_LC_10_12_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_LC_10_12_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_LC_10_12_5 (
            .in0(N__27595),
            .in1(N__48341),
            .in2(N__27572),
            .in3(N__56159),
            .lcout(n22226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_210_LC_10_12_6.C_ON=1'b0;
    defparam i1_4_lut_adj_210_LC_10_12_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_210_LC_10_12_6.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_210_LC_10_12_6 (
            .in0(N__27551),
            .in1(N__54945),
            .in2(N__49826),
            .in3(N__46571),
            .lcout(n11931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i0_LC_10_12_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i0_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i0_LC_10_12_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i0_LC_10_12_7  (
            .in0(N__53175),
            .in1(N__52989),
            .in2(N__29398),
            .in3(N__34051),
            .lcout(buf_adcdata_iac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57870),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i14_LC_10_13_0.C_ON=1'b0;
    defparam buf_dds1_i14_LC_10_13_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i14_LC_10_13_0.LUT_INIT=16'b1101100000000000;
    LogicCell40 buf_dds1_i14_LC_10_13_0 (
            .in0(N__38571),
            .in1(N__43168),
            .in2(N__36954),
            .in3(N__38471),
            .lcout(buf_dds1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57883),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i0_LC_10_13_1.C_ON=1'b0;
    defparam buf_dds1_i0_LC_10_13_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i0_LC_10_13_1.LUT_INIT=16'b1000100010100000;
    LogicCell40 buf_dds1_i0_LC_10_13_1 (
            .in0(N__38470),
            .in1(N__41163),
            .in2(N__27537),
            .in3(N__38572),
            .lcout(buf_dds1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57883),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_240_LC_10_13_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_240_LC_10_13_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_240_LC_10_13_2.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_240_LC_10_13_2 (
            .in0(N__53568),
            .in1(N__48537),
            .in2(_gnd_net_),
            .in3(N__31880),
            .lcout(n20663),
            .ltout(n20663_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_10_13_3.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_10_13_3.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_10_13_3.LUT_INIT=16'b1111111111111011;
    LogicCell40 i2_3_lut_4_lut_LC_10_13_3 (
            .in0(N__53995),
            .in1(N__52378),
            .in2(N__27731),
            .in3(N__36582),
            .lcout(n10614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_243_LC_10_13_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_243_LC_10_13_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_243_LC_10_13_4.LUT_INIT=16'b1111111101110111;
    LogicCell40 i1_2_lut_3_lut_adj_243_LC_10_13_4 (
            .in0(N__56144),
            .in1(N__48536),
            .in2(_gnd_net_),
            .in3(N__31881),
            .lcout(n11354),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15263_2_lut_3_lut_LC_10_13_5.C_ON=1'b0;
    defparam i15263_2_lut_3_lut_LC_10_13_5.SEQ_MODE=4'b0000;
    defparam i15263_2_lut_3_lut_LC_10_13_5.LUT_INIT=16'b0000000001010000;
    LogicCell40 i15263_2_lut_3_lut_LC_10_13_5 (
            .in0(N__53997),
            .in1(_gnd_net_),
            .in2(N__46028),
            .in3(N__52380),
            .lcout(n14_adj_1544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i0_LC_10_13_6.C_ON=1'b0;
    defparam buf_dds0_i0_LC_10_13_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i0_LC_10_13_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i0_LC_10_13_6 (
            .in0(N__49754),
            .in1(N__31188),
            .in2(N__41168),
            .in3(N__38965),
            .lcout(buf_dds0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57883),
            .ce(),
            .sr(_gnd_net_));
    defparam i15302_2_lut_3_lut_LC_10_13_7.C_ON=1'b0;
    defparam i15302_2_lut_3_lut_LC_10_13_7.SEQ_MODE=4'b0000;
    defparam i15302_2_lut_3_lut_LC_10_13_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15302_2_lut_3_lut_LC_10_13_7 (
            .in0(N__53996),
            .in1(N__41162),
            .in2(_gnd_net_),
            .in3(N__52379),
            .lcout(n14_adj_1533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_2_lut_LC_10_14_0.C_ON=1'b1;
    defparam add_131_2_lut_LC_10_14_0.SEQ_MODE=4'b0000;
    defparam add_131_2_lut_LC_10_14_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_2_lut_LC_10_14_0 (
            .in0(N__31031),
            .in1(N__31029),
            .in2(N__39136),
            .in3(N__27728),
            .lcout(n7_adj_1531),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(n19384),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_3_lut_LC_10_14_1.C_ON=1'b1;
    defparam add_131_3_lut_LC_10_14_1.SEQ_MODE=4'b0000;
    defparam add_131_3_lut_LC_10_14_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_3_lut_LC_10_14_1 (
            .in0(N__38606),
            .in1(N__38605),
            .in2(N__39140),
            .in3(N__27725),
            .lcout(n7_adj_1566),
            .ltout(),
            .carryin(n19384),
            .carryout(n19385),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_4_lut_LC_10_14_2.C_ON=1'b1;
    defparam add_131_4_lut_LC_10_14_2.SEQ_MODE=4'b0000;
    defparam add_131_4_lut_LC_10_14_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_4_lut_LC_10_14_2 (
            .in0(N__36182),
            .in1(N__36181),
            .in2(N__39137),
            .in3(N__27722),
            .lcout(n7_adj_1564),
            .ltout(),
            .carryin(n19385),
            .carryout(n19386),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_5_lut_LC_10_14_3.C_ON=1'b1;
    defparam add_131_5_lut_LC_10_14_3.SEQ_MODE=4'b0000;
    defparam add_131_5_lut_LC_10_14_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_5_lut_LC_10_14_3 (
            .in0(N__36047),
            .in1(N__36046),
            .in2(N__39141),
            .in3(N__27719),
            .lcout(n7_adj_1562),
            .ltout(),
            .carryin(n19386),
            .carryout(n19387),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_6_lut_LC_10_14_4.C_ON=1'b1;
    defparam add_131_6_lut_LC_10_14_4.SEQ_MODE=4'b0000;
    defparam add_131_6_lut_LC_10_14_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_6_lut_LC_10_14_4 (
            .in0(N__38768),
            .in1(N__38767),
            .in2(N__39138),
            .in3(N__27716),
            .lcout(n7_adj_1560),
            .ltout(),
            .carryin(n19387),
            .carryout(n19388),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_7_lut_LC_10_14_5.C_ON=1'b1;
    defparam add_131_7_lut_LC_10_14_5.SEQ_MODE=4'b0000;
    defparam add_131_7_lut_LC_10_14_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_7_lut_LC_10_14_5 (
            .in0(N__31051),
            .in1(N__31050),
            .in2(N__39142),
            .in3(N__27929),
            .lcout(n17409),
            .ltout(),
            .carryin(n19388),
            .carryout(n19389),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_8_lut_LC_10_14_6.C_ON=1'b1;
    defparam add_131_8_lut_LC_10_14_6.SEQ_MODE=4'b0000;
    defparam add_131_8_lut_LC_10_14_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_8_lut_LC_10_14_6 (
            .in0(N__41963),
            .in1(N__41962),
            .in2(N__39139),
            .in3(N__27926),
            .lcout(n7_adj_1558),
            .ltout(),
            .carryin(n19389),
            .carryout(n19390),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_9_lut_LC_10_14_7.C_ON=1'b1;
    defparam add_131_9_lut_LC_10_14_7.SEQ_MODE=4'b0000;
    defparam add_131_9_lut_LC_10_14_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_9_lut_LC_10_14_7 (
            .in0(N__27862),
            .in1(N__27861),
            .in2(N__39143),
            .in3(N__27923),
            .lcout(n7_adj_1556),
            .ltout(),
            .carryin(n19390),
            .carryout(n19391),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_10_lut_LC_10_15_0.C_ON=1'b1;
    defparam add_131_10_lut_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam add_131_10_lut_LC_10_15_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_10_lut_LC_10_15_0 (
            .in0(N__27919),
            .in1(N__27912),
            .in2(N__39153),
            .in3(N__27890),
            .lcout(n7_adj_1554),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(n19392),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_131_11_lut_LC_10_15_1.C_ON=1'b0;
    defparam add_131_11_lut_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam add_131_11_lut_LC_10_15_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_131_11_lut_LC_10_15_1 (
            .in0(N__27985),
            .in1(N__27986),
            .in2(N__39158),
            .in3(N__27887),
            .lcout(n7_adj_1552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_2_i16_3_lut_LC_10_15_2.C_ON=1'b0;
    defparam mux_135_Mux_2_i16_3_lut_LC_10_15_2.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_2_i16_3_lut_LC_10_15_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_2_i16_3_lut_LC_10_15_2 (
            .in0(N__27879),
            .in1(N__28442),
            .in2(_gnd_net_),
            .in3(N__56309),
            .lcout(n16_adj_1515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i2_LC_10_15_3.C_ON=1'b0;
    defparam buf_dds1_i2_LC_10_15_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i2_LC_10_15_3.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i2_LC_10_15_3 (
            .in0(N__27883),
            .in1(N__38559),
            .in2(N__47143),
            .in3(N__38451),
            .lcout(buf_dds1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57912),
            .ce(),
            .sr(_gnd_net_));
    defparam i6404_3_lut_LC_10_15_4.C_ON=1'b0;
    defparam i6404_3_lut_LC_10_15_4.SEQ_MODE=4'b0000;
    defparam i6404_3_lut_LC_10_15_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6404_3_lut_LC_10_15_4 (
            .in0(N__47672),
            .in1(N__27863),
            .in2(_gnd_net_),
            .in3(N__41709),
            .lcout(n8_adj_1557),
            .ltout(n8_adj_1557_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_7_i15_4_lut_LC_10_15_5.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_7_i15_4_lut_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_7_i15_4_lut_LC_10_15_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_365_Mux_7_i15_4_lut_LC_10_15_5 (
            .in0(N__49830),
            .in1(N__54953),
            .in2(N__27839),
            .in3(N__27835),
            .lcout(data_index_9_N_216_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6384_3_lut_LC_10_15_6.C_ON=1'b0;
    defparam i6384_3_lut_LC_10_15_6.SEQ_MODE=4'b0000;
    defparam i6384_3_lut_LC_10_15_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6384_3_lut_LC_10_15_6 (
            .in0(N__45521),
            .in1(N__27984),
            .in2(_gnd_net_),
            .in3(N__41708),
            .lcout(n8_adj_1553),
            .ltout(n8_adj_1553_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i9_LC_10_15_7.C_ON=1'b0;
    defparam data_index_i9_LC_10_15_7.SEQ_MODE=4'b1000;
    defparam data_index_i9_LC_10_15_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i9_LC_10_15_7 (
            .in0(N__49831),
            .in1(N__54954),
            .in2(N__27989),
            .in3(N__28255),
            .lcout(data_index_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57912),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_response_312_LC_10_16_0.C_ON=1'b0;
    defparam comm_response_312_LC_10_16_0.SEQ_MODE=4'b1000;
    defparam comm_response_312_LC_10_16_0.LUT_INIT=16'b0000001001010010;
    LogicCell40 comm_response_312_LC_10_16_0 (
            .in0(N__54976),
            .in1(N__52389),
            .in2(N__54140),
            .in3(N__53590),
            .lcout(ICE_GPMI_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57926),
            .ce(N__27944),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_297_LC_10_16_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_297_LC_10_16_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_297_LC_10_16_1.LUT_INIT=16'b1111101000110010;
    LogicCell40 i1_3_lut_4_lut_adj_297_LC_10_16_1 (
            .in0(N__53589),
            .in1(N__52416),
            .in2(N__51590),
            .in3(N__54975),
            .lcout(n11401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_227_LC_10_16_3.C_ON=1'b0;
    defparam i1_3_lut_adj_227_LC_10_16_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_227_LC_10_16_3.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_3_lut_adj_227_LC_10_16_3 (
            .in0(N__51585),
            .in1(N__39482),
            .in2(_gnd_net_),
            .in3(N__54971),
            .lcout(n11866),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18158_2_lut_3_lut_LC_10_16_4.C_ON=1'b0;
    defparam i18158_2_lut_3_lut_LC_10_16_4.SEQ_MODE=4'b0000;
    defparam i18158_2_lut_3_lut_LC_10_16_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i18158_2_lut_3_lut_LC_10_16_4 (
            .in0(N__54090),
            .in1(N__52387),
            .in2(_gnd_net_),
            .in3(N__53587),
            .lcout(),
            .ltout(n20772_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_183_LC_10_16_5.C_ON=1'b0;
    defparam i1_4_lut_adj_183_LC_10_16_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_183_LC_10_16_5.LUT_INIT=16'b1000101011001111;
    LogicCell40 i1_4_lut_adj_183_LC_10_16_5 (
            .in0(N__51584),
            .in1(N__54973),
            .in2(N__27935),
            .in3(N__34795),
            .lcout(n11835),
            .ltout(n11835_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_69_LC_10_16_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_69_LC_10_16_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_69_LC_10_16_6.LUT_INIT=16'b0000111100101111;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_69_LC_10_16_6 (
            .in0(N__54974),
            .in1(N__54005),
            .in2(N__27932),
            .in3(N__52388),
            .lcout(n16763),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_282_LC_10_16_7.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_282_LC_10_16_7.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_282_LC_10_16_7.LUT_INIT=16'b1110111011111111;
    LogicCell40 i2_2_lut_3_lut_adj_282_LC_10_16_7 (
            .in0(N__53588),
            .in1(N__54091),
            .in2(_gnd_net_),
            .in3(N__54972),
            .lcout(n11377),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i14_LC_10_17_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i14_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i14_LC_10_17_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \SIG_DDS.tmp_buf_i14_LC_10_17_0  (
            .in0(N__50306),
            .in1(N__50138),
            .in2(N__36925),
            .in3(N__28097),
            .lcout(\SIG_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i11_LC_10_17_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i11_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i11_LC_10_17_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i11_LC_10_17_1  (
            .in0(N__50133),
            .in1(N__50303),
            .in2(N__28130),
            .in3(N__40457),
            .lcout(\SIG_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i10_LC_10_17_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i10_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i10_LC_10_17_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i10_LC_10_17_2  (
            .in0(N__50302),
            .in1(N__50132),
            .in2(N__28007),
            .in3(N__28145),
            .lcout(\SIG_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i13_LC_10_17_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i13_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i13_LC_10_17_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i13_LC_10_17_3  (
            .in0(N__50137),
            .in1(N__50305),
            .in2(N__28085),
            .in3(N__28121),
            .lcout(\SIG_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i6_LC_10_17_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i6_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i6_LC_10_17_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i6_LC_10_17_4  (
            .in0(N__50308),
            .in1(N__50140),
            .in2(N__28451),
            .in3(N__31301),
            .lcout(\SIG_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i12_LC_10_17_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i12_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i12_LC_10_17_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \SIG_DDS.tmp_buf_i12_LC_10_17_5  (
            .in0(N__40333),
            .in1(N__28091),
            .in2(N__50157),
            .in3(N__50304),
            .lcout(\SIG_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i15_LC_10_17_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i15_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i15_LC_10_17_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i15_LC_10_17_6  (
            .in0(N__50307),
            .in1(N__50139),
            .in2(N__28073),
            .in3(N__28056),
            .lcout(tmp_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i9_LC_10_17_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i9_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i9_LC_10_17_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i9_LC_10_17_7  (
            .in0(N__50141),
            .in1(N__50309),
            .in2(N__28352),
            .in3(N__28034),
            .lcout(\SIG_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57939),
            .ce(N__31400),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i7_LC_10_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i7_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i7_LC_10_18_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i7_LC_10_18_1  (
            .in0(N__50184),
            .in1(N__50300),
            .in2(N__27998),
            .in3(N__44567),
            .lcout(\SIG_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i5_LC_10_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i5_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i5_LC_10_18_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i5_LC_10_18_2  (
            .in0(N__50299),
            .in1(N__50183),
            .in2(N__28391),
            .in3(N__36548),
            .lcout(\SIG_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i2_LC_10_18_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i2_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i2_LC_10_18_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i2_LC_10_18_3  (
            .in0(N__50180),
            .in1(N__50296),
            .in2(N__28316),
            .in3(N__28441),
            .lcout(\SIG_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i4_LC_10_18_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i4_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i4_LC_10_18_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \SIG_DDS.tmp_buf_i4_LC_10_18_4  (
            .in0(N__50298),
            .in1(N__50182),
            .in2(N__28421),
            .in3(N__28271),
            .lcout(\SIG_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i8_LC_10_18_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i8_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i8_LC_10_18_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i8_LC_10_18_5  (
            .in0(N__50185),
            .in1(N__50301),
            .in2(N__28382),
            .in3(N__28373),
            .lcout(\SIG_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i1_LC_10_18_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i1_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i1_LC_10_18_6 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \SIG_DDS.tmp_buf_i1_LC_10_18_6  (
            .in0(N__50295),
            .in1(N__28340),
            .in2(N__31409),
            .in3(N__50179),
            .lcout(\SIG_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i3_LC_10_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i3_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i3_LC_10_18_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i3_LC_10_18_7  (
            .in0(N__50181),
            .in1(N__50297),
            .in2(N__28307),
            .in3(N__28298),
            .lcout(\SIG_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57950),
            .ce(N__31390),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_9_i15_4_lut_LC_10_19_6.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_9_i15_4_lut_LC_10_19_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_9_i15_4_lut_LC_10_19_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_365_Mux_9_i15_4_lut_LC_10_19_6 (
            .in0(N__54982),
            .in1(N__28265),
            .in2(N__49829),
            .in3(N__28256),
            .lcout(data_index_9_N_216_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i2_LC_11_3_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i2_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i2_LC_11_3_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i2_LC_11_3_1  (
            .in0(N__34652),
            .in1(N__35410),
            .in2(N__28541),
            .in3(N__28606),
            .lcout(buf_adcdata_vac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57805),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_LC_11_3_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_11_3_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_LC_11_3_2  (
            .in0(N__31324),
            .in1(N__31429),
            .in2(N__31472),
            .in3(N__31447),
            .lcout(\ADC_VDC.genclk.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_2_i19_3_lut_LC_11_3_3.C_ON=1'b0;
    defparam mux_136_Mux_2_i19_3_lut_LC_11_3_3.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_2_i19_3_lut_LC_11_3_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_136_Mux_2_i19_3_lut_LC_11_3_3 (
            .in0(N__28643),
            .in1(N__28605),
            .in2(_gnd_net_),
            .in3(N__56341),
            .lcout(),
            .ltout(n19_adj_1646_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_2_i22_3_lut_LC_11_3_4.C_ON=1'b0;
    defparam mux_136_Mux_2_i22_3_lut_LC_11_3_4.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_2_i22_3_lut_LC_11_3_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_136_Mux_2_i22_3_lut_LC_11_3_4 (
            .in0(_gnd_net_),
            .in1(N__28581),
            .in2(N__28565),
            .in3(N__49098),
            .lcout(),
            .ltout(n22_adj_1647_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_2_i30_3_lut_LC_11_3_5.C_ON=1'b0;
    defparam mux_136_Mux_2_i30_3_lut_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_2_i30_3_lut_LC_11_3_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_136_Mux_2_i30_3_lut_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(N__28562),
            .in2(N__28544),
            .in3(N__48719),
            .lcout(n30_adj_1648),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_11_3_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_11_3_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i11_LC_11_3_6  (
            .in0(N__35409),
            .in1(N__28537),
            .in2(N__28824),
            .in3(N__34453),
            .lcout(cmd_rdadctmp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57805),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19102_2_lut_LC_11_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19102_2_lut_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19102_2_lut_LC_11_4_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ADC_VDC.genclk.i19102_2_lut_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__33677),
            .in2(_gnd_net_),
            .in3(N__40171),
            .lcout(\ADC_VDC.genclk.n11751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_3_i19_3_lut_LC_11_5_0.C_ON=1'b0;
    defparam mux_136_Mux_3_i19_3_lut_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_3_i19_3_lut_LC_11_5_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_136_Mux_3_i19_3_lut_LC_11_5_0 (
            .in0(N__28514),
            .in1(N__28794),
            .in2(_gnd_net_),
            .in3(N__56291),
            .lcout(),
            .ltout(n19_adj_1642_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_3_i22_3_lut_LC_11_5_1.C_ON=1'b0;
    defparam mux_136_Mux_3_i22_3_lut_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_3_i22_3_lut_LC_11_5_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_136_Mux_3_i22_3_lut_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(N__28464),
            .in2(N__28493),
            .in3(N__49052),
            .lcout(),
            .ltout(n22_adj_1643_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_3_i30_3_lut_LC_11_5_2.C_ON=1'b0;
    defparam mux_136_Mux_3_i30_3_lut_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_3_i30_3_lut_LC_11_5_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_136_Mux_3_i30_3_lut_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(N__28490),
            .in2(N__28475),
            .in3(N__48681),
            .lcout(n30_adj_1644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_5_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i3_LC_11_5_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i3_LC_11_5_3  (
            .in0(N__53200),
            .in1(N__52999),
            .in2(N__28781),
            .in3(N__28465),
            .lcout(buf_adcdata_iac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_5_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i3_LC_11_5_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i3_LC_11_5_4  (
            .in0(N__34621),
            .in1(N__35412),
            .in2(N__28834),
            .in3(N__28795),
            .lcout(buf_adcdata_vac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_11_5_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_11_5_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i11_LC_11_5_5  (
            .in0(N__52077),
            .in1(N__28669),
            .in2(N__28780),
            .in3(N__53000),
            .lcout(cmd_rdadctmp_11_adj_1439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_11_5_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_11_5_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i12_LC_11_5_6  (
            .in0(N__52998),
            .in1(N__28776),
            .in2(N__28755),
            .in3(N__52078),
            .lcout(cmd_rdadctmp_12_adj_1438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57811),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_11_5_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_11_5_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i17_LC_11_5_7  (
            .in0(N__35411),
            .in1(N__30580),
            .in2(N__30430),
            .in3(N__34452),
            .lcout(cmd_rdadctmp_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57811),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i7_LC_11_6_0.C_ON=1'b0;
    defparam comm_buf_5__i7_LC_11_6_0.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i7_LC_11_6_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i7_LC_11_6_0 (
            .in0(N__51406),
            .in1(N__28724),
            .in2(_gnd_net_),
            .in3(N__54138),
            .lcout(comm_buf_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57816),
            .ce(N__31493),
            .sr(N__31673));
    defparam comm_buf_5__i6_LC_11_6_1.C_ON=1'b0;
    defparam comm_buf_5__i6_LC_11_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i6_LC_11_6_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i6_LC_11_6_1 (
            .in0(N__54136),
            .in1(N__40245),
            .in2(_gnd_net_),
            .in3(N__28706),
            .lcout(comm_buf_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57816),
            .ce(N__31493),
            .sr(N__31673));
    defparam comm_buf_5__i5_LC_11_6_2.C_ON=1'b0;
    defparam comm_buf_5__i5_LC_11_6_2.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i5_LC_11_6_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i5_LC_11_6_2 (
            .in0(N__51055),
            .in1(N__28691),
            .in2(_gnd_net_),
            .in3(N__54137),
            .lcout(comm_buf_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57816),
            .ce(N__31493),
            .sr(N__31673));
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i10_LC_11_7_0  (
            .in0(N__29365),
            .in1(N__52958),
            .in2(N__28668),
            .in3(N__52090),
            .lcout(cmd_rdadctmp_10_adj_1440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57819),
            .ce(),
            .sr(_gnd_net_));
    defparam i36_4_lut_4_lut_LC_11_7_2.C_ON=1'b0;
    defparam i36_4_lut_4_lut_LC_11_7_2.SEQ_MODE=4'b0000;
    defparam i36_4_lut_4_lut_LC_11_7_2.LUT_INIT=16'b0010010011110100;
    LogicCell40 i36_4_lut_4_lut_LC_11_7_2 (
            .in0(N__56252),
            .in1(N__48195),
            .in2(N__48718),
            .in3(N__48997),
            .lcout(),
            .ltout(n30_adj_1480_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_96_LC_11_7_3.C_ON=1'b0;
    defparam i1_4_lut_adj_96_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_96_LC_11_7_3.LUT_INIT=16'b1111000100000000;
    LogicCell40 i1_4_lut_adj_96_LC_11_7_3 (
            .in0(N__48998),
            .in1(N__48266),
            .in2(N__28940),
            .in3(N__45187),
            .lcout(comm_state_3_N_420_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_1_i19_3_lut_LC_11_7_4.C_ON=1'b0;
    defparam mux_136_Mux_1_i19_3_lut_LC_11_7_4.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_1_i19_3_lut_LC_11_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_136_Mux_1_i19_3_lut_LC_11_7_4 (
            .in0(N__56253),
            .in1(N__28937),
            .in2(_gnd_net_),
            .in3(N__34741),
            .lcout(),
            .ltout(n19_adj_1491_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_1_i22_3_lut_LC_11_7_5.C_ON=1'b0;
    defparam mux_136_Mux_1_i22_3_lut_LC_11_7_5.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_1_i22_3_lut_LC_11_7_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_136_Mux_1_i22_3_lut_LC_11_7_5 (
            .in0(N__48999),
            .in1(_gnd_net_),
            .in2(N__28916),
            .in3(N__28905),
            .lcout(n22_adj_1489),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i1_LC_11_7_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i1_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i1_LC_11_7_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i1_LC_11_7_6  (
            .in0(N__28906),
            .in1(N__53183),
            .in2(N__29369),
            .in3(N__52959),
            .lcout(buf_adcdata_iac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57819),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19528_LC_11_7_7.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19528_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19528_LC_11_7_7.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19528_LC_11_7_7 (
            .in0(N__48194),
            .in1(N__29495),
            .in2(N__28892),
            .in3(N__56251),
            .lcout(n22160),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i15_LC_11_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i15_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i15_LC_11_8_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i15_LC_11_8_0  (
            .in0(N__29165),
            .in1(N__33366),
            .in2(N__29341),
            .in3(N__28871),
            .lcout(buf_adcdata_vdc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i14_LC_11_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i14_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i14_LC_11_8_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i14_LC_11_8_1  (
            .in0(N__33363),
            .in1(N__29169),
            .in2(N__38101),
            .in3(N__28859),
            .lcout(buf_adcdata_vdc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i13_LC_11_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i13_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i13_LC_11_8_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i13_LC_11_8_2  (
            .in0(N__29164),
            .in1(N__33365),
            .in2(N__46666),
            .in3(N__28847),
            .lcout(buf_adcdata_vdc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_37_LC_11_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_37_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_37_LC_11_8_3 .LUT_INIT=16'b1011000011100000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_37_LC_11_8_3  (
            .in0(N__33125),
            .in1(N__32868),
            .in2(N__33373),
            .in3(N__33522),
            .lcout(\ADC_VDC.n12915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i16_LC_11_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i16_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i16_LC_11_8_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i16_LC_11_8_4  (
            .in0(N__29166),
            .in1(N__33367),
            .in2(N__29278),
            .in3(N__29216),
            .lcout(buf_adcdata_vdc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i0_LC_11_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i0_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i0_LC_11_8_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i0_LC_11_8_5  (
            .in0(N__33362),
            .in1(N__29168),
            .in2(N__33982),
            .in3(N__29204),
            .lcout(buf_adcdata_vdc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i22_LC_11_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i22_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i22_LC_11_8_6 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \ADC_VDC.ADC_DATA_i22_LC_11_8_6  (
            .in0(N__29167),
            .in1(N__29189),
            .in2(N__33374),
            .in3(N__31924),
            .lcout(buf_adcdata_vdc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i9_LC_11_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i9_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i9_LC_11_8_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i9_LC_11_8_7  (
            .in0(N__33364),
            .in1(N__29170),
            .in2(N__30850),
            .in3(N__29045),
            .lcout(buf_adcdata_vdc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40107),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_166_LC_11_9_0.C_ON=1'b0;
    defparam i1_4_lut_adj_166_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_166_LC_11_9_0.LUT_INIT=16'b1101000011000000;
    LogicCell40 i1_4_lut_adj_166_LC_11_9_0 (
            .in0(N__52432),
            .in1(N__54902),
            .in2(N__51569),
            .in3(N__40496),
            .lcout(n11918),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i18_LC_11_9_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i18_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i18_LC_11_9_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i18_LC_11_9_1  (
            .in0(N__34583),
            .in1(N__35392),
            .in2(N__34244),
            .in3(N__29028),
            .lcout(buf_adcdata_vac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57831),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i2_LC_11_9_2.C_ON=1'b0;
    defparam comm_buf_6__i2_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i2_LC_11_9_2.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i2_LC_11_9_2 (
            .in0(N__43303),
            .in1(N__54903),
            .in2(N__47248),
            .in3(N__51319),
            .lcout(comm_buf_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57831),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i6_LC_11_9_3.C_ON=1'b0;
    defparam comm_buf_6__i6_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i6_LC_11_9_3.LUT_INIT=16'b0100111001000100;
    LogicCell40 comm_buf_6__i6_LC_11_9_3 (
            .in0(N__51320),
            .in1(N__43201),
            .in2(N__54961),
            .in3(N__40246),
            .lcout(comm_buf_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57831),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_11_9_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_11_9_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i27_LC_11_9_4  (
            .in0(N__35391),
            .in1(N__34240),
            .in2(N__29451),
            .in3(N__34432),
            .lcout(cmd_rdadctmp_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57831),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i6_LC_11_9_5.C_ON=1'b0;
    defparam buf_cfgRTD_i6_LC_11_9_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i6_LC_11_9_5.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_cfgRTD_i6_LC_11_9_5 (
            .in0(N__29005),
            .in1(N__49628),
            .in2(N__43175),
            .in3(N__29488),
            .lcout(buf_cfgRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57831),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i19_LC_11_9_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i19_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i19_LC_11_9_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i19_LC_11_9_6  (
            .in0(N__35390),
            .in1(N__34584),
            .in2(N__29452),
            .in3(N__29421),
            .lcout(buf_adcdata_vac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57831),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_11_10_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_11_10_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i9_LC_11_10_0  (
            .in0(N__29399),
            .in1(N__52991),
            .in2(N__29364),
            .in3(N__52094),
            .lcout(cmd_rdadctmp_9_adj_1441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57841),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i15_LC_11_10_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i15_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i15_LC_11_10_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i15_LC_11_10_1  (
            .in0(N__29311),
            .in1(N__34595),
            .in2(N__29261),
            .in3(N__35342),
            .lcout(buf_adcdata_vac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57841),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_7_i19_3_lut_LC_11_10_2.C_ON=1'b0;
    defparam mux_135_Mux_7_i19_3_lut_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_7_i19_3_lut_LC_11_10_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_7_i19_3_lut_LC_11_10_2 (
            .in0(N__29345),
            .in1(N__29310),
            .in2(_gnd_net_),
            .in3(N__55943),
            .lcout(n19_adj_1502),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22016_bdd_4_lut_LC_11_10_3.C_ON=1'b0;
    defparam n22016_bdd_4_lut_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam n22016_bdd_4_lut_LC_11_10_3.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22016_bdd_4_lut_LC_11_10_3 (
            .in0(N__30396),
            .in1(N__29297),
            .in2(N__29285),
            .in3(N__48098),
            .lcout(n22019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_11_10_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_11_10_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i23_LC_11_10_4  (
            .in0(N__35341),
            .in1(N__32002),
            .in2(N__29260),
            .in3(N__34425),
            .lcout(cmd_rdadctmp_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57841),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_11_10_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_11_10_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i24_LC_11_10_5  (
            .in0(N__34426),
            .in1(N__35343),
            .in2(N__29240),
            .in3(N__29256),
            .lcout(cmd_rdadctmp_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57841),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_303_LC_11_10_6.C_ON=1'b0;
    defparam i1_2_lut_adj_303_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_303_LC_11_10_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_303_LC_11_10_6 (
            .in0(_gnd_net_),
            .in1(N__34960),
            .in2(_gnd_net_),
            .in3(N__35044),
            .lcout(n20590),
            .ltout(n20590_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i16_LC_11_10_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i16_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i16_LC_11_10_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i16_LC_11_10_7  (
            .in0(N__30397),
            .in1(N__29238),
            .in2(N__30413),
            .in3(N__35344),
            .lcout(buf_adcdata_vac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57841),
            .ce(),
            .sr(_gnd_net_));
    defparam data_count_i0_i0_LC_11_11_0.C_ON=1'b1;
    defparam data_count_i0_i0_LC_11_11_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i0_LC_11_11_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i0_LC_11_11_0 (
            .in0(_gnd_net_),
            .in1(N__41437),
            .in2(N__30303),
            .in3(_gnd_net_),
            .lcout(data_count_0),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(n19345),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i1_LC_11_11_1.C_ON=1'b1;
    defparam data_count_i0_i1_LC_11_11_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i1_LC_11_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i1_LC_11_11_1 (
            .in0(_gnd_net_),
            .in1(N__30189),
            .in2(_gnd_net_),
            .in3(N__30170),
            .lcout(data_count_1),
            .ltout(),
            .carryin(n19345),
            .carryout(n19346),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i2_LC_11_11_2.C_ON=1'b1;
    defparam data_count_i0_i2_LC_11_11_2.SEQ_MODE=4'b1000;
    defparam data_count_i0_i2_LC_11_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i2_LC_11_11_2 (
            .in0(_gnd_net_),
            .in1(N__30075),
            .in2(_gnd_net_),
            .in3(N__30056),
            .lcout(data_count_2),
            .ltout(),
            .carryin(n19346),
            .carryout(n19347),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i3_LC_11_11_3.C_ON=1'b1;
    defparam data_count_i0_i3_LC_11_11_3.SEQ_MODE=4'b1000;
    defparam data_count_i0_i3_LC_11_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i3_LC_11_11_3 (
            .in0(_gnd_net_),
            .in1(N__29973),
            .in2(_gnd_net_),
            .in3(N__29951),
            .lcout(data_count_3),
            .ltout(),
            .carryin(n19347),
            .carryout(n19348),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i4_LC_11_11_4.C_ON=1'b1;
    defparam data_count_i0_i4_LC_11_11_4.SEQ_MODE=4'b1000;
    defparam data_count_i0_i4_LC_11_11_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i4_LC_11_11_4 (
            .in0(_gnd_net_),
            .in1(N__29859),
            .in2(_gnd_net_),
            .in3(N__29837),
            .lcout(data_count_4),
            .ltout(),
            .carryin(n19348),
            .carryout(n19349),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i5_LC_11_11_5.C_ON=1'b1;
    defparam data_count_i0_i5_LC_11_11_5.SEQ_MODE=4'b1000;
    defparam data_count_i0_i5_LC_11_11_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i5_LC_11_11_5 (
            .in0(_gnd_net_),
            .in1(N__29757),
            .in2(_gnd_net_),
            .in3(N__29735),
            .lcout(data_count_5),
            .ltout(),
            .carryin(n19349),
            .carryout(n19350),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i6_LC_11_11_6.C_ON=1'b1;
    defparam data_count_i0_i6_LC_11_11_6.SEQ_MODE=4'b1000;
    defparam data_count_i0_i6_LC_11_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i6_LC_11_11_6 (
            .in0(_gnd_net_),
            .in1(N__29649),
            .in2(_gnd_net_),
            .in3(N__29627),
            .lcout(data_count_6),
            .ltout(),
            .carryin(n19350),
            .carryout(n19351),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i7_LC_11_11_7.C_ON=1'b1;
    defparam data_count_i0_i7_LC_11_11_7.SEQ_MODE=4'b1000;
    defparam data_count_i0_i7_LC_11_11_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i7_LC_11_11_7 (
            .in0(_gnd_net_),
            .in1(N__29538),
            .in2(_gnd_net_),
            .in3(N__29519),
            .lcout(data_count_7),
            .ltout(),
            .carryin(n19351),
            .carryout(n19352),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__41886),
            .sr(N__41839));
    defparam data_count_i0_i8_LC_11_12_0.C_ON=1'b1;
    defparam data_count_i0_i8_LC_11_12_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i8_LC_11_12_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i8_LC_11_12_0 (
            .in0(_gnd_net_),
            .in1(N__30720),
            .in2(_gnd_net_),
            .in3(N__30698),
            .lcout(data_count_8),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(n19353),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__41875),
            .sr(N__41840));
    defparam data_count_i0_i9_LC_11_12_1.C_ON=1'b0;
    defparam data_count_i0_i9_LC_11_12_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i9_LC_11_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i9_LC_11_12_1 (
            .in0(_gnd_net_),
            .in1(N__30606),
            .in2(_gnd_net_),
            .in3(N__30695),
            .lcout(data_count_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__41875),
            .sr(N__41840));
    defparam \ADC_VAC.ADC_DATA_i8_LC_11_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i8_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i8_LC_11_13_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i8_LC_11_13_0  (
            .in0(N__30511),
            .in1(N__34624),
            .in2(N__35422),
            .in3(N__30584),
            .lcout(buf_adcdata_vac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57871),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_0_i19_3_lut_LC_11_13_1.C_ON=1'b0;
    defparam mux_135_Mux_0_i19_3_lut_LC_11_13_1.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_0_i19_3_lut_LC_11_13_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_135_Mux_0_i19_3_lut_LC_11_13_1 (
            .in0(N__56072),
            .in1(N__30545),
            .in2(_gnd_net_),
            .in3(N__30510),
            .lcout(n19_adj_1487),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i9_LC_11_13_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i9_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i9_LC_11_13_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i9_LC_11_13_2  (
            .in0(N__34622),
            .in1(N__35394),
            .in2(N__30446),
            .in3(N__30823),
            .lcout(buf_adcdata_vac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_11_13_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_11_13_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i21_LC_11_13_3  (
            .in0(N__30909),
            .in1(N__52990),
            .in2(N__51094),
            .in3(N__52076),
            .lcout(cmd_rdadctmp_21_adj_1429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i10_LC_11_13_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i10_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i10_LC_11_13_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i10_LC_11_13_4  (
            .in0(N__30460),
            .in1(N__34623),
            .in2(N__30971),
            .in3(N__35395),
            .lcout(buf_adcdata_vac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57871),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_2_i19_3_lut_LC_11_13_5.C_ON=1'b0;
    defparam mux_135_Mux_2_i19_3_lut_LC_11_13_5.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_2_i19_3_lut_LC_11_13_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_135_Mux_2_i19_3_lut_LC_11_13_5 (
            .in0(N__56071),
            .in1(N__30497),
            .in2(_gnd_net_),
            .in3(N__30459),
            .lcout(n19_adj_1516),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_11_13_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_11_13_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i18_LC_11_13_6  (
            .in0(N__30966),
            .in1(N__34430),
            .in2(N__30445),
            .in3(N__35396),
            .lcout(cmd_rdadctmp_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_11_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_11_13_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i19_LC_11_13_7  (
            .in0(N__35393),
            .in1(N__30967),
            .in2(N__34518),
            .in3(N__34431),
            .lcout(cmd_rdadctmp_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i12_LC_11_14_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i12_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i12_LC_11_14_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i12_LC_11_14_0  (
            .in0(N__38148),
            .in1(N__51095),
            .in2(N__53156),
            .in3(N__52936),
            .lcout(buf_adcdata_iac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57884),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i13_LC_11_14_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i13_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i13_LC_11_14_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i13_LC_11_14_1  (
            .in0(N__52933),
            .in1(N__53116),
            .in2(N__43578),
            .in3(N__30911),
            .lcout(buf_adcdata_iac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57884),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_5_i23_3_lut_LC_11_14_2.C_ON=1'b0;
    defparam mux_134_Mux_5_i23_3_lut_LC_11_14_2.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_5_i23_3_lut_LC_11_14_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_134_Mux_5_i23_3_lut_LC_11_14_2 (
            .in0(N__30946),
            .in1(N__56236),
            .in2(_gnd_net_),
            .in3(N__38843),
            .lcout(n23_adj_1536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_11_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_11_14_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i22_LC_11_14_3  (
            .in0(N__52935),
            .in1(N__30910),
            .in2(N__30876),
            .in3(N__52075),
            .lcout(cmd_rdadctmp_22_adj_1428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57884),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i0_LC_11_14_4.C_ON=1'b0;
    defparam data_index_i0_LC_11_14_4.SEQ_MODE=4'b1000;
    defparam data_index_i0_LC_11_14_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i0_LC_11_14_4 (
            .in0(N__54947),
            .in1(N__31009),
            .in2(N__49827),
            .in3(N__30895),
            .lcout(data_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57884),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i14_LC_11_14_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i14_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i14_LC_11_14_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i14_LC_11_14_5  (
            .in0(N__52934),
            .in1(N__53117),
            .in2(N__30877),
            .in3(N__38352),
            .lcout(buf_adcdata_iac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57884),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i12_LC_11_14_6.C_ON=1'b0;
    defparam buf_dds0_i12_LC_11_14_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i12_LC_11_14_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i12_LC_11_14_6 (
            .in0(N__49750),
            .in1(N__38972),
            .in2(N__44169),
            .in3(N__40326),
            .lcout(buf_dds0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57884),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_1_i19_3_lut_LC_11_14_7.C_ON=1'b0;
    defparam mux_135_Mux_1_i19_3_lut_LC_11_14_7.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_1_i19_3_lut_LC_11_14_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_135_Mux_1_i19_3_lut_LC_11_14_7 (
            .in0(N__56237),
            .in1(N__30854),
            .in2(_gnd_net_),
            .in3(N__30813),
            .lcout(n19_adj_1520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15012_3_lut_LC_11_15_0.C_ON=1'b0;
    defparam i15012_3_lut_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam i15012_3_lut_LC_11_15_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 i15012_3_lut_LC_11_15_0 (
            .in0(N__45916),
            .in1(N__31052),
            .in2(_gnd_net_),
            .in3(N__41728),
            .lcout(n17411),
            .ltout(n17411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15014_4_lut_LC_11_15_1.C_ON=1'b0;
    defparam i15014_4_lut_LC_11_15_1.SEQ_MODE=4'b0000;
    defparam i15014_4_lut_LC_11_15_1.LUT_INIT=16'b0111010100100000;
    LogicCell40 i15014_4_lut_LC_11_15_1 (
            .in0(N__54888),
            .in1(N__49663),
            .in2(N__31169),
            .in3(N__31066),
            .lcout(data_index_9_N_216_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i5_LC_11_15_2.C_ON=1'b0;
    defparam data_index_i5_LC_11_15_2.SEQ_MODE=4'b1000;
    defparam data_index_i5_LC_11_15_2.LUT_INIT=16'b0000110010101010;
    LogicCell40 data_index_i5_LC_11_15_2 (
            .in0(N__31067),
            .in1(N__31058),
            .in2(N__49758),
            .in3(N__54891),
            .lcout(data_index_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57896),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_11_15_3.C_ON=1'b0;
    defparam i3_4_lut_LC_11_15_3.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_11_15_3.LUT_INIT=16'b1111111011111111;
    LogicCell40 i3_4_lut_LC_11_15_3 (
            .in0(N__53586),
            .in1(N__48232),
            .in2(N__34864),
            .in3(N__49003),
            .lcout(n8828),
            .ltout(n8828_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4419_3_lut_LC_11_15_4.C_ON=1'b0;
    defparam i4419_3_lut_LC_11_15_4.SEQ_MODE=4'b0000;
    defparam i4419_3_lut_LC_11_15_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 i4419_3_lut_LC_11_15_4 (
            .in0(_gnd_net_),
            .in1(N__41158),
            .in2(N__31034),
            .in3(N__31030),
            .lcout(n8_adj_1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i11_LC_11_15_5.C_ON=1'b0;
    defparam buf_dds1_i11_LC_11_15_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i11_LC_11_15_5.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i11_LC_11_15_5 (
            .in0(N__38555),
            .in1(N__40479),
            .in2(N__44309),
            .in3(N__38454),
            .lcout(buf_dds1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57896),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i13_LC_11_15_6.C_ON=1'b0;
    defparam buf_dds1_i13_LC_11_15_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i13_LC_11_15_6.LUT_INIT=16'b1110001011101110;
    LogicCell40 buf_dds1_i13_LC_11_15_6 (
            .in0(N__30993),
            .in1(N__38556),
            .in2(N__47591),
            .in3(N__54890),
            .lcout(buf_dds1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57896),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i2_LC_11_15_7.C_ON=1'b0;
    defparam data_index_i2_LC_11_15_7.SEQ_MODE=4'b1000;
    defparam data_index_i2_LC_11_15_7.LUT_INIT=16'b0100010011100100;
    LogicCell40 data_index_i2_LC_11_15_7 (
            .in0(N__54889),
            .in1(N__39427),
            .in2(N__39449),
            .in3(N__49664),
            .lcout(data_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57896),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_6_i16_3_lut_LC_11_16_0.C_ON=1'b0;
    defparam mux_135_Mux_6_i16_3_lut_LC_11_16_0.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_6_i16_3_lut_LC_11_16_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_6_i16_3_lut_LC_11_16_0 (
            .in0(N__31275),
            .in1(N__31299),
            .in2(_gnd_net_),
            .in3(N__56244),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9341_1_lut_LC_11_16_1.C_ON=1'b0;
    defparam i9341_1_lut_LC_11_16_1.SEQ_MODE=4'b0000;
    defparam i9341_1_lut_LC_11_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i9341_1_lut_LC_11_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50002),
            .lcout(n11757),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i7_LC_11_16_2.C_ON=1'b0;
    defparam buf_dds1_i7_LC_11_16_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i7_LC_11_16_2.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i7_LC_11_16_2 (
            .in0(N__44586),
            .in1(N__38561),
            .in2(N__47681),
            .in3(N__38453),
            .lcout(buf_dds1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57913),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i6_LC_11_16_3.C_ON=1'b0;
    defparam buf_dds0_i6_LC_11_16_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i6_LC_11_16_3.LUT_INIT=16'b0000110010101010;
    LogicCell40 buf_dds0_i6_LC_11_16_3 (
            .in0(N__31300),
            .in1(N__52507),
            .in2(N__49832),
            .in3(N__38954),
            .lcout(buf_dds0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57913),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i6_LC_11_16_4.C_ON=1'b0;
    defparam buf_dds1_i6_LC_11_16_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i6_LC_11_16_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i6_LC_11_16_4 (
            .in0(N__31276),
            .in1(N__38560),
            .in2(N__52511),
            .in3(N__38452),
            .lcout(buf_dds1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57913),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i14_LC_11_16_7.C_ON=1'b0;
    defparam acadc_skipCount_i14_LC_11_16_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i14_LC_11_16_7.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i14_LC_11_16_7 (
            .in0(N__49767),
            .in1(N__49373),
            .in2(N__32371),
            .in3(N__43155),
            .lcout(acadc_skipCount_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57913),
            .ce(),
            .sr(_gnd_net_));
    defparam wdtick_cnt_3774_3775__i1_LC_11_17_0.C_ON=1'b0;
    defparam wdtick_cnt_3774_3775__i1_LC_11_17_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3774_3775__i1_LC_11_17_0.LUT_INIT=16'b0011001100010001;
    LogicCell40 wdtick_cnt_3774_3775__i1_LC_11_17_0 (
            .in0(N__31206),
            .in1(N__31245),
            .in2(_gnd_net_),
            .in3(N__31226),
            .lcout(wdtick_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32734),
            .ce(N__31262),
            .sr(N__40696));
    defparam wdtick_cnt_3774_3775__i3_LC_11_17_1.C_ON=1'b0;
    defparam wdtick_cnt_3774_3775__i3_LC_11_17_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3774_3775__i3_LC_11_17_1.LUT_INIT=16'b0101101010100000;
    LogicCell40 wdtick_cnt_3774_3775__i3_LC_11_17_1 (
            .in0(N__31228),
            .in1(_gnd_net_),
            .in2(N__31250),
            .in3(N__31207),
            .lcout(wdtick_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32734),
            .ce(N__31262),
            .sr(N__40696));
    defparam wdtick_cnt_3774_3775__i2_LC_11_17_2.C_ON=1'b0;
    defparam wdtick_cnt_3774_3775__i2_LC_11_17_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3774_3775__i2_LC_11_17_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 wdtick_cnt_3774_3775__i2_LC_11_17_2 (
            .in0(_gnd_net_),
            .in1(N__31244),
            .in2(_gnd_net_),
            .in3(N__31227),
            .lcout(wdtick_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32734),
            .ce(N__31262),
            .sr(N__40696));
    defparam wdtick_flag_299_LC_11_18_0.C_ON=1'b0;
    defparam wdtick_flag_299_LC_11_18_0.SEQ_MODE=4'b1010;
    defparam wdtick_flag_299_LC_11_18_0.LUT_INIT=16'b1111111100010000;
    LogicCell40 wdtick_flag_299_LC_11_18_0 (
            .in0(N__31249),
            .in1(N__31229),
            .in2(N__31211),
            .in3(N__49998),
            .lcout(wdtick_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32733),
            .ce(),
            .sr(N__40697));
    defparam \SIG_DDS.tmp_buf_i0_LC_11_19_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i0_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i0_LC_11_19_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i0_LC_11_19_0  (
            .in0(N__50178),
            .in1(N__50249),
            .in2(N__44728),
            .in3(N__31193),
            .lcout(\SIG_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57951),
            .ce(N__31389),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19098_4_lut_LC_11_19_3 .C_ON=1'b0;
    defparam \SIG_DDS.i19098_4_lut_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19098_4_lut_LC_11_19_3 .LUT_INIT=16'b1010101000100110;
    LogicCell40 \SIG_DDS.i19098_4_lut_LC_11_19_3  (
            .in0(N__50248),
            .in1(N__50366),
            .in2(N__44811),
            .in3(N__50177),
            .lcout(\SIG_DDS.n12738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15029_2_lut_LC_12_1_7.C_ON=1'b0;
    defparam i15029_2_lut_LC_12_1_7.SEQ_MODE=4'b0000;
    defparam i15029_2_lut_LC_12_1_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i15029_2_lut_LC_12_1_7 (
            .in0(N__35716),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31369),
            .lcout(OUT_SYNCCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0off_i0_LC_12_3_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i0_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i0_LC_12_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i0_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(N__32609),
            .in2(_gnd_net_),
            .in3(N__31334),
            .lcout(\ADC_VDC.genclk.t0off_0 ),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(\ADC_VDC.genclk.n19468 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i1_LC_12_3_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i1_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i1_LC_12_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i1_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__32579),
            .in2(N__57324),
            .in3(N__31331),
            .lcout(\ADC_VDC.genclk.t0off_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19468 ),
            .carryout(\ADC_VDC.genclk.n19469 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i2_LC_12_3_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i2_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i2_LC_12_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i2_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(N__57251),
            .in2(N__31328),
            .in3(N__31313),
            .lcout(\ADC_VDC.genclk.t0off_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19469 ),
            .carryout(\ADC_VDC.genclk.n19470 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i3_LC_12_3_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i3_LC_12_3_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0off_i3_LC_12_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i3_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__32678),
            .in2(N__57325),
            .in3(N__31310),
            .lcout(\ADC_VDC.genclk.t0off_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19470 ),
            .carryout(\ADC_VDC.genclk.n19471 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i4_LC_12_3_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i4_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i4_LC_12_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i4_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__57255),
            .in2(N__32597),
            .in3(N__31307),
            .lcout(\ADC_VDC.genclk.t0off_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19471 ),
            .carryout(\ADC_VDC.genclk.n19472 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i5_LC_12_3_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i5_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i5_LC_12_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i5_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__32665),
            .in2(N__57326),
            .in3(N__31304),
            .lcout(\ADC_VDC.genclk.t0off_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19472 ),
            .carryout(\ADC_VDC.genclk.n19473 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i6_LC_12_3_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i6_LC_12_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i6_LC_12_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i6_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__57259),
            .in2(N__32624),
            .in3(N__31475),
            .lcout(\ADC_VDC.genclk.t0off_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19473 ),
            .carryout(\ADC_VDC.genclk.n19474 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i7_LC_12_3_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i7_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i7_LC_12_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i7_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(N__31471),
            .in2(N__57327),
            .in3(N__31457),
            .lcout(\ADC_VDC.genclk.t0off_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19474 ),
            .carryout(\ADC_VDC.genclk.n19475 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__31601),
            .sr(N__33880));
    defparam \ADC_VDC.genclk.t0off_i8_LC_12_4_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i8_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i8_LC_12_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i8_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(N__32651),
            .in2(N__57384),
            .in3(N__31454),
            .lcout(\ADC_VDC.genclk.t0off_8 ),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(\ADC_VDC.genclk.n19476 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i9_LC_12_4_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i9_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i9_LC_12_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i9_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(N__57346),
            .in2(N__32549),
            .in3(N__31451),
            .lcout(\ADC_VDC.genclk.t0off_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19476 ),
            .carryout(\ADC_VDC.genclk.n19477 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i10_LC_12_4_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i10_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i10_LC_12_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i10_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(N__31448),
            .in2(N__57381),
            .in3(N__31436),
            .lcout(\ADC_VDC.genclk.t0off_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19477 ),
            .carryout(\ADC_VDC.genclk.n19478 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i11_LC_12_4_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i11_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i11_LC_12_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i11_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(N__57334),
            .in2(N__32519),
            .in3(N__31433),
            .lcout(\ADC_VDC.genclk.t0off_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19478 ),
            .carryout(\ADC_VDC.genclk.n19479 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i12_LC_12_4_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i12_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i12_LC_12_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i12_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(N__31430),
            .in2(N__57382),
            .in3(N__31418),
            .lcout(\ADC_VDC.genclk.t0off_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19479 ),
            .carryout(\ADC_VDC.genclk.n19480 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i13_LC_12_4_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i13_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i13_LC_12_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i13_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(N__57338),
            .in2(N__32693),
            .in3(N__31415),
            .lcout(\ADC_VDC.genclk.t0off_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19480 ),
            .carryout(\ADC_VDC.genclk.n19481 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i14_LC_12_4_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i14_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i14_LC_12_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i14_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(N__32561),
            .in2(N__57383),
            .in3(N__31412),
            .lcout(\ADC_VDC.genclk.t0off_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19481 ),
            .carryout(\ADC_VDC.genclk.n19482 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam \ADC_VDC.genclk.t0off_i15_LC_12_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0off_i15_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i15_LC_12_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0off_i15_LC_12_4_7  (
            .in0(N__32533),
            .in1(N__57342),
            .in2(_gnd_net_),
            .in3(N__31604),
            .lcout(\ADC_VDC.genclk.t0off_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__31597),
            .sr(N__33872));
    defparam i19_4_lut_adj_249_LC_12_5_0.C_ON=1'b0;
    defparam i19_4_lut_adj_249_LC_12_5_0.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_249_LC_12_5_0.LUT_INIT=16'b1011000100010001;
    LogicCell40 i19_4_lut_adj_249_LC_12_5_0 (
            .in0(N__54174),
            .in1(N__37516),
            .in2(N__54383),
            .in3(N__31625),
            .lcout(),
            .ltout(n12_adj_1615_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_250_LC_12_5_1.C_ON=1'b0;
    defparam i1_3_lut_adj_250_LC_12_5_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_250_LC_12_5_1.LUT_INIT=16'b1100110011000000;
    LogicCell40 i1_3_lut_adj_250_LC_12_5_1 (
            .in0(_gnd_net_),
            .in1(N__42785),
            .in2(N__31577),
            .in3(N__50926),
            .lcout(n12236),
            .ltout(n12236_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12388_2_lut_LC_12_5_2.C_ON=1'b0;
    defparam i12388_2_lut_LC_12_5_2.SEQ_MODE=4'b0000;
    defparam i12388_2_lut_LC_12_5_2.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12388_2_lut_LC_12_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31574),
            .in3(N__54911),
            .lcout(n14801),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i0_LC_12_5_3.C_ON=1'b0;
    defparam comm_buf_5__i0_LC_12_5_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i0_LC_12_5_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i0_LC_12_5_3 (
            .in0(N__50776),
            .in1(N__31571),
            .in2(_gnd_net_),
            .in3(N__54177),
            .lcout(comm_buf_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57806),
            .ce(N__31489),
            .sr(N__31669));
    defparam comm_buf_5__i1_LC_12_5_4.C_ON=1'b0;
    defparam comm_buf_5__i1_LC_12_5_4.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i1_LC_12_5_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i1_LC_12_5_4 (
            .in0(N__54175),
            .in1(N__45365),
            .in2(_gnd_net_),
            .in3(N__31556),
            .lcout(comm_buf_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57806),
            .ce(N__31489),
            .sr(N__31669));
    defparam comm_buf_5__i2_LC_12_5_5.C_ON=1'b0;
    defparam comm_buf_5__i2_LC_12_5_5.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i2_LC_12_5_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i2_LC_12_5_5 (
            .in0(N__47241),
            .in1(N__31538),
            .in2(_gnd_net_),
            .in3(N__54178),
            .lcout(comm_buf_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57806),
            .ce(N__31489),
            .sr(N__31669));
    defparam comm_buf_5__i3_LC_12_5_6.C_ON=1'b0;
    defparam comm_buf_5__i3_LC_12_5_6.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i3_LC_12_5_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i3_LC_12_5_6 (
            .in0(N__54176),
            .in1(N__40776),
            .in2(_gnd_net_),
            .in3(N__31523),
            .lcout(comm_buf_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57806),
            .ce(N__31489),
            .sr(N__31669));
    defparam comm_buf_5__i4_LC_12_5_7.C_ON=1'b0;
    defparam comm_buf_5__i4_LC_12_5_7.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i4_LC_12_5_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i4_LC_12_5_7 (
            .in0(N__40645),
            .in1(N__31508),
            .in2(_gnd_net_),
            .in3(N__54179),
            .lcout(comm_buf_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57806),
            .ce(N__31489),
            .sr(N__31669));
    defparam mux_143_Mux_4_i2_3_lut_LC_12_6_0.C_ON=1'b0;
    defparam mux_143_Mux_4_i2_3_lut_LC_12_6_0.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_4_i2_3_lut_LC_12_6_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_143_Mux_4_i2_3_lut_LC_12_6_0 (
            .in0(N__36986),
            .in1(N__31823),
            .in2(_gnd_net_),
            .in3(N__54382),
            .lcout(),
            .ltout(n2_adj_1587_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i4_LC_12_6_1.C_ON=1'b0;
    defparam comm_tx_buf_i4_LC_12_6_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i4_LC_12_6_1.LUT_INIT=16'b1111101001000100;
    LogicCell40 comm_tx_buf_i4_LC_12_6_1 (
            .in0(N__50687),
            .in1(N__31631),
            .in2(N__31655),
            .in3(N__31637),
            .lcout(comm_tx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57808),
            .ce(N__46223),
            .sr(N__46140));
    defparam i18721_2_lut_LC_12_6_2.C_ON=1'b0;
    defparam i18721_2_lut_LC_12_6_2.SEQ_MODE=4'b0000;
    defparam i18721_2_lut_LC_12_6_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18721_2_lut_LC_12_6_2 (
            .in0(_gnd_net_),
            .in1(N__31904),
            .in2(_gnd_net_),
            .in3(N__54379),
            .lcout(n21324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_4_i4_3_lut_LC_12_6_3.C_ON=1'b0;
    defparam mux_143_Mux_4_i4_3_lut_LC_12_6_3.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_4_i4_3_lut_LC_12_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_143_Mux_4_i4_3_lut_LC_12_6_3 (
            .in0(N__54380),
            .in1(N__31652),
            .in2(_gnd_net_),
            .in3(N__37721),
            .lcout(),
            .ltout(n4_adj_1588_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19504_LC_12_6_4.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19504_LC_12_6_4.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19504_LC_12_6_4.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_index_1__bdd_4_lut_19504_LC_12_6_4 (
            .in0(N__31646),
            .in1(N__50554),
            .in2(N__31640),
            .in3(N__50686),
            .lcout(n22136),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_4_i1_3_lut_LC_12_6_5.C_ON=1'b0;
    defparam mux_143_Mux_4_i1_3_lut_LC_12_6_5.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_4_i1_3_lut_LC_12_6_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_143_Mux_4_i1_3_lut_LC_12_6_5 (
            .in0(N__54381),
            .in1(N__51182),
            .in2(_gnd_net_),
            .in3(N__44120),
            .lcout(n1_adj_1586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_12_6_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_12_6_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_12_6_6.LUT_INIT=16'b0011000000000000;
    LogicCell40 i1_2_lut_3_lut_LC_12_6_6 (
            .in0(_gnd_net_),
            .in1(N__50553),
            .in2(N__43070),
            .in3(N__50685),
            .lcout(n19006),
            .ltout(n19006_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_246_LC_12_6_7.C_ON=1'b0;
    defparam i19_4_lut_adj_246_LC_12_6_7.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_246_LC_12_6_7.LUT_INIT=16'b0100000001110011;
    LogicCell40 i19_4_lut_adj_246_LC_12_6_7 (
            .in0(N__54378),
            .in1(N__54150),
            .in2(N__31619),
            .in3(N__37517),
            .lcout(n12_adj_1639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i7_LC_12_7_0.C_ON=1'b0;
    defparam comm_buf_2__i7_LC_12_7_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i7_LC_12_7_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i7_LC_12_7_0 (
            .in0(N__54166),
            .in1(N__51393),
            .in2(_gnd_net_),
            .in3(N__31616),
            .lcout(comm_buf_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57813),
            .ce(N__34217),
            .sr(N__34190));
    defparam comm_buf_2__i6_LC_12_7_1.C_ON=1'b0;
    defparam comm_buf_2__i6_LC_12_7_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i6_LC_12_7_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i6_LC_12_7_1 (
            .in0(N__40234),
            .in1(N__31862),
            .in2(_gnd_net_),
            .in3(N__54168),
            .lcout(comm_buf_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57813),
            .ce(N__34217),
            .sr(N__34190));
    defparam comm_buf_2__i5_LC_12_7_2.C_ON=1'b0;
    defparam comm_buf_2__i5_LC_12_7_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i5_LC_12_7_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i5_LC_12_7_2 (
            .in0(N__54165),
            .in1(N__51043),
            .in2(_gnd_net_),
            .in3(N__31850),
            .lcout(comm_buf_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57813),
            .ce(N__34217),
            .sr(N__34190));
    defparam comm_buf_2__i4_LC_12_7_3.C_ON=1'b0;
    defparam comm_buf_2__i4_LC_12_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i4_LC_12_7_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_2__i4_LC_12_7_3 (
            .in0(N__54139),
            .in1(N__31838),
            .in2(_gnd_net_),
            .in3(N__40646),
            .lcout(comm_buf_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57813),
            .ce(N__34217),
            .sr(N__34190));
    defparam comm_buf_2__i3_LC_12_7_4.C_ON=1'b0;
    defparam comm_buf_2__i3_LC_12_7_4.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i3_LC_12_7_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i3_LC_12_7_4 (
            .in0(N__54164),
            .in1(N__40793),
            .in2(_gnd_net_),
            .in3(N__31817),
            .lcout(comm_buf_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57813),
            .ce(N__34217),
            .sr(N__34190));
    defparam comm_buf_2__i2_LC_12_7_5.C_ON=1'b0;
    defparam comm_buf_2__i2_LC_12_7_5.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i2_LC_12_7_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i2_LC_12_7_5 (
            .in0(N__47242),
            .in1(N__31805),
            .in2(_gnd_net_),
            .in3(N__54167),
            .lcout(comm_buf_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57813),
            .ce(N__34217),
            .sr(N__34190));
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_12_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_12_8_0 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i23_LC_12_8_0  (
            .in0(N__31793),
            .in1(N__31763),
            .in2(N__31744),
            .in3(N__32869),
            .lcout(\ADC_VDC.cmd_rdadctmp_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40131),
            .ce(N__31724),
            .sr(N__31718));
    defparam \RTD.i2_3_lut_LC_12_8_1 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_LC_12_8_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \RTD.i2_3_lut_LC_12_8_1  (
            .in0(N__33766),
            .in1(N__33789),
            .in2(_gnd_net_),
            .in3(N__33806),
            .lcout(\RTD.n17720 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_6_i23_3_lut_LC_12_8_6.C_ON=1'b0;
    defparam mux_134_Mux_6_i23_3_lut_LC_12_8_6.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_6_i23_3_lut_LC_12_8_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_134_Mux_6_i23_3_lut_LC_12_8_6 (
            .in0(N__45017),
            .in1(N__56106),
            .in2(_gnd_net_),
            .in3(N__32372),
            .lcout(n23_adj_1534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i7_LC_12_9_1.C_ON=1'b0;
    defparam comm_cmd_i7_LC_12_9_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i7_LC_12_9_1.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i7_LC_12_9_1 (
            .in0(N__32100),
            .in1(N__32027),
            .in2(N__40569),
            .in3(N__51405),
            .lcout(comm_cmd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57821),
            .ce(),
            .sr(_gnd_net_));
    defparam n22160_bdd_4_lut_LC_12_9_2.C_ON=1'b0;
    defparam n22160_bdd_4_lut_LC_12_9_2.SEQ_MODE=4'b0000;
    defparam n22160_bdd_4_lut_LC_12_9_2.LUT_INIT=16'b1111110000100010;
    LogicCell40 n22160_bdd_4_lut_LC_12_9_2 (
            .in0(N__31966),
            .in1(N__48094),
            .in2(N__31928),
            .in3(N__31913),
            .lcout(n22163),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_12_9_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_12_9_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i20_LC_12_9_3  (
            .in0(N__34519),
            .in1(N__34410),
            .in2(N__34686),
            .in3(N__35376),
            .lcout(cmd_rdadctmp_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57821),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i3_LC_12_9_4.C_ON=1'b0;
    defparam comm_buf_6__i3_LC_12_9_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i3_LC_12_9_4.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i3_LC_12_9_4 (
            .in0(N__37618),
            .in1(N__54907),
            .in2(N__40801),
            .in3(N__51312),
            .lcout(comm_buf_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57821),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i4_LC_12_9_5.C_ON=1'b0;
    defparam comm_buf_6__i4_LC_12_9_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i4_LC_12_9_5.LUT_INIT=16'b0100111001000100;
    LogicCell40 comm_buf_6__i4_LC_12_9_5 (
            .in0(N__51313),
            .in1(N__31903),
            .in2(N__54962),
            .in3(N__40654),
            .lcout(comm_buf_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57821),
            .ce(),
            .sr(_gnd_net_));
    defparam i18755_2_lut_LC_12_9_6.C_ON=1'b0;
    defparam i18755_2_lut_LC_12_9_6.SEQ_MODE=4'b0000;
    defparam i18755_2_lut_LC_12_9_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18755_2_lut_LC_12_9_6 (
            .in0(_gnd_net_),
            .in1(N__53561),
            .in2(_gnd_net_),
            .in3(N__31889),
            .lcout(n20962),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i2_LC_12_10_0.C_ON=1'b0;
    defparam comm_cmd_i2_LC_12_10_0.SEQ_MODE=4'b1000;
    defparam comm_cmd_i2_LC_12_10_0.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i2_LC_12_10_0 (
            .in0(N__48816),
            .in1(N__32121),
            .in2(N__47252),
            .in3(N__32032),
            .lcout(comm_cmd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i1_LC_12_10_1.C_ON=1'b0;
    defparam comm_cmd_i1_LC_12_10_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i1_LC_12_10_1.LUT_INIT=16'b1100101000001010;
    LogicCell40 comm_cmd_i1_LC_12_10_1 (
            .in0(N__47998),
            .in1(N__45377),
            .in2(N__32044),
            .in3(N__32120),
            .lcout(comm_cmd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_12_10_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_12_10_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i22_LC_12_10_2  (
            .in0(N__35406),
            .in1(N__34702),
            .in2(N__32003),
            .in3(N__34428),
            .lcout(cmd_rdadctmp_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_12_10_3.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_12_10_3.LUT_INIT=16'b1101110111111111;
    LogicCell40 i2_2_lut_3_lut_LC_12_10_3 (
            .in0(N__47997),
            .in1(N__55816),
            .in2(_gnd_net_),
            .in3(N__48815),
            .lcout(n10733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_12_10_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_12_10_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i21_LC_12_10_4  (
            .in0(N__35405),
            .in1(N__34701),
            .in2(N__34687),
            .in3(N__34427),
            .lcout(cmd_rdadctmp_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i17_LC_12_10_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i17_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i17_LC_12_10_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i17_LC_12_10_5  (
            .in0(N__34594),
            .in1(N__35408),
            .in2(N__34487),
            .in3(N__43947),
            .lcout(buf_adcdata_vac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i0_LC_12_10_6.C_ON=1'b0;
    defparam comm_cmd_i0_LC_12_10_6.SEQ_MODE=4'b1000;
    defparam comm_cmd_i0_LC_12_10_6.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i0_LC_12_10_6 (
            .in0(N__55817),
            .in1(N__50783),
            .in2(N__32123),
            .in3(N__32028),
            .lcout(comm_cmd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i14_LC_12_10_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i14_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i14_LC_12_10_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i14_LC_12_10_7  (
            .in0(N__34593),
            .in1(N__35407),
            .in2(N__38077),
            .in3(N__32001),
            .lcout(buf_adcdata_vac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57829),
            .ce(),
            .sr(_gnd_net_));
    defparam data_idxvec_i0_LC_12_11_0.C_ON=1'b1;
    defparam data_idxvec_i0_LC_12_11_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i0_LC_12_11_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i0_LC_12_11_0 (
            .in0(N__46547),
            .in1(N__54803),
            .in2(N__41234),
            .in3(N__31985),
            .lcout(data_idxvec_0),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(n19393),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i1_LC_12_11_1.C_ON=1'b1;
    defparam data_idxvec_i1_LC_12_11_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i1_LC_12_11_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i1_LC_12_11_1 (
            .in0(N__46816),
            .in1(N__54807),
            .in2(N__43421),
            .in3(N__31982),
            .lcout(data_idxvec_1),
            .ltout(),
            .carryin(n19393),
            .carryout(n19394),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i2_LC_12_11_2.C_ON=1'b1;
    defparam data_idxvec_i2_LC_12_11_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i2_LC_12_11_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i2_LC_12_11_2 (
            .in0(N__44054),
            .in1(N__54804),
            .in2(N__46870),
            .in3(N__31979),
            .lcout(data_idxvec_2),
            .ltout(),
            .carryin(n19394),
            .carryout(n19395),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i3_LC_12_11_3.C_ON=1'b1;
    defparam data_idxvec_i3_LC_12_11_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i3_LC_12_11_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i3_LC_12_11_3 (
            .in0(N__47843),
            .in1(N__54808),
            .in2(N__37880),
            .in3(N__31976),
            .lcout(data_idxvec_3),
            .ltout(),
            .carryin(n19395),
            .carryout(n19396),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i4_LC_12_11_4.C_ON=1'b1;
    defparam data_idxvec_i4_LC_12_11_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i4_LC_12_11_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i4_LC_12_11_4 (
            .in0(N__51119),
            .in1(N__54805),
            .in2(N__38218),
            .in3(N__31973),
            .lcout(data_idxvec_4),
            .ltout(),
            .carryin(n19396),
            .carryout(n19397),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i5_LC_12_11_5.C_ON=1'b1;
    defparam data_idxvec_i5_LC_12_11_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i5_LC_12_11_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i5_LC_12_11_5 (
            .in0(N__47322),
            .in1(N__54809),
            .in2(N__43489),
            .in3(N__31970),
            .lcout(data_idxvec_5),
            .ltout(),
            .carryin(n19397),
            .carryout(n19398),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i6_LC_12_11_6.C_ON=1'b1;
    defparam data_idxvec_i6_LC_12_11_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i6_LC_12_11_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i6_LC_12_11_6 (
            .in0(N__52175),
            .in1(N__54806),
            .in2(N__37786),
            .in3(N__32174),
            .lcout(data_idxvec_6),
            .ltout(),
            .carryin(n19398),
            .carryout(n19399),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i7_LC_12_11_7.C_ON=1'b1;
    defparam data_idxvec_i7_LC_12_11_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i7_LC_12_11_7.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i7_LC_12_11_7 (
            .in0(N__47606),
            .in1(N__54810),
            .in2(N__49249),
            .in3(N__32171),
            .lcout(data_idxvec_7),
            .ltout(),
            .carryin(n19399),
            .carryout(n19400),
            .clk(N__57839),
            .ce(N__39061),
            .sr(_gnd_net_));
    defparam data_idxvec_i8_LC_12_12_0.C_ON=1'b1;
    defparam data_idxvec_i8_LC_12_12_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i8_LC_12_12_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i8_LC_12_12_0 (
            .in0(N__44478),
            .in1(N__54892),
            .in2(N__41584),
            .in3(N__32168),
            .lcout(data_idxvec_8),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(n19401),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i9_LC_12_12_1.C_ON=1'b1;
    defparam data_idxvec_i9_LC_12_12_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i9_LC_12_12_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i9_LC_12_12_1 (
            .in0(N__47462),
            .in1(N__54899),
            .in2(N__44347),
            .in3(N__32165),
            .lcout(data_idxvec_9),
            .ltout(),
            .carryin(n19401),
            .carryout(n19402),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i10_LC_12_12_2.C_ON=1'b1;
    defparam data_idxvec_i10_LC_12_12_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i10_LC_12_12_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i10_LC_12_12_2 (
            .in0(N__39313),
            .in1(N__54893),
            .in2(N__34165),
            .in3(N__32162),
            .lcout(data_idxvec_10),
            .ltout(),
            .carryin(n19402),
            .carryout(n19403),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i11_LC_12_12_3.C_ON=1'b1;
    defparam data_idxvec_i11_LC_12_12_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i11_LC_12_12_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i11_LC_12_12_3 (
            .in0(N__39274),
            .in1(N__54900),
            .in2(N__40864),
            .in3(N__32159),
            .lcout(data_idxvec_11),
            .ltout(),
            .carryin(n19403),
            .carryout(n19404),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i12_LC_12_12_4.C_ON=1'b1;
    defparam data_idxvec_i12_LC_12_12_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i12_LC_12_12_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i12_LC_12_12_4 (
            .in0(N__44077),
            .in1(N__54894),
            .in2(N__40945),
            .in3(N__32156),
            .lcout(data_idxvec_12),
            .ltout(),
            .carryin(n19404),
            .carryout(n19405),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i13_LC_12_12_5.C_ON=1'b1;
    defparam data_idxvec_i13_LC_12_12_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i13_LC_12_12_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i13_LC_12_12_5 (
            .in0(N__47587),
            .in1(N__54901),
            .in2(N__32149),
            .in3(N__32129),
            .lcout(data_idxvec_13),
            .ltout(),
            .carryin(n19405),
            .carryout(n19406),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i14_LC_12_12_6.C_ON=1'b1;
    defparam data_idxvec_i14_LC_12_12_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i14_LC_12_12_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i14_LC_12_12_6 (
            .in0(N__39190),
            .in1(N__54895),
            .in2(N__36274),
            .in3(N__32126),
            .lcout(data_idxvec_14),
            .ltout(),
            .carryin(n19406),
            .carryout(n19407),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam data_idxvec_i15_LC_12_12_7.C_ON=1'b0;
    defparam data_idxvec_i15_LC_12_12_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i15_LC_12_12_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i15_LC_12_12_7 (
            .in0(N__46795),
            .in1(N__32267),
            .in2(N__54960),
            .in3(N__32291),
            .lcout(data_idxvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57849),
            .ce(N__39065),
            .sr(_gnd_net_));
    defparam i18129_4_lut_LC_12_13_0.C_ON=1'b0;
    defparam i18129_4_lut_LC_12_13_0.SEQ_MODE=4'b0000;
    defparam i18129_4_lut_LC_12_13_0.LUT_INIT=16'b1111111111001010;
    LogicCell40 i18129_4_lut_LC_12_13_0 (
            .in0(N__36715),
            .in1(N__36418),
            .in2(N__41050),
            .in3(N__36335),
            .lcout(n20742),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22166_bdd_4_lut_LC_12_13_1.C_ON=1'b0;
    defparam n22166_bdd_4_lut_LC_12_13_1.SEQ_MODE=4'b0000;
    defparam n22166_bdd_4_lut_LC_12_13_1.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22166_bdd_4_lut_LC_12_13_1 (
            .in0(N__49011),
            .in1(N__41303),
            .in2(N__47765),
            .in3(N__32240),
            .lcout(),
            .ltout(n22169_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1545458_i1_3_lut_LC_12_13_2.C_ON=1'b0;
    defparam i1545458_i1_3_lut_LC_12_13_2.SEQ_MODE=4'b0000;
    defparam i1545458_i1_3_lut_LC_12_13_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 i1545458_i1_3_lut_LC_12_13_2 (
            .in0(N__48714),
            .in1(_gnd_net_),
            .in2(N__32288),
            .in3(N__32285),
            .lcout(n30_adj_1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19099_4_lut_LC_12_13_3.C_ON=1'b0;
    defparam i19099_4_lut_LC_12_13_3.SEQ_MODE=4'b0000;
    defparam i19099_4_lut_LC_12_13_3.LUT_INIT=16'b0101000100110011;
    LogicCell40 i19099_4_lut_LC_12_13_3 (
            .in0(N__36419),
            .in1(N__36716),
            .in2(N__36062),
            .in3(N__41035),
            .lcout(),
            .ltout(n20568_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_309_LC_12_13_4.C_ON=1'b0;
    defparam eis_end_309_LC_12_13_4.SEQ_MODE=4'b1000;
    defparam eis_end_309_LC_12_13_4.LUT_INIT=16'b1100110010101100;
    LogicCell40 eis_end_309_LC_12_13_4 (
            .in0(N__36717),
            .in1(N__32255),
            .in2(N__32270),
            .in3(N__36336),
            .lcout(eis_end),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_end_309C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_7_i26_3_lut_LC_12_13_5.C_ON=1'b0;
    defparam mux_134_Mux_7_i26_3_lut_LC_12_13_5.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i26_3_lut_LC_12_13_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_134_Mux_7_i26_3_lut_LC_12_13_5 (
            .in0(N__32266),
            .in1(N__56073),
            .in2(_gnd_net_),
            .in3(N__32254),
            .lcout(),
            .ltout(n26_adj_1528_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19523_LC_12_13_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19523_LC_12_13_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19523_LC_12_13_6.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19523_LC_12_13_6 (
            .in0(N__55586),
            .in1(N__48228),
            .in2(N__32243),
            .in3(N__49010),
            .lcout(n22166),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_trig_310_LC_12_13_7.C_ON=1'b0;
    defparam acadc_trig_310_LC_12_13_7.SEQ_MODE=4'b1000;
    defparam acadc_trig_310_LC_12_13_7.LUT_INIT=16'b1111000000100010;
    LogicCell40 acadc_trig_310_LC_12_13_7 (
            .in0(N__41036),
            .in1(N__36718),
            .in2(N__32217),
            .in3(N__32234),
            .lcout(acadc_trig),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_end_309C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i14176_4_lut_LC_12_14_0.C_ON=1'b0;
    defparam i14176_4_lut_LC_12_14_0.SEQ_MODE=4'b0000;
    defparam i14176_4_lut_LC_12_14_0.LUT_INIT=16'b1100010111001111;
    LogicCell40 i14176_4_lut_LC_12_14_0 (
            .in0(N__41626),
            .in1(N__43925),
            .in2(N__36725),
            .in3(N__36191),
            .lcout(),
            .ltout(n16594_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i0_LC_12_14_1.C_ON=1'b0;
    defparam eis_state_i0_LC_12_14_1.SEQ_MODE=4'b1010;
    defparam eis_state_i0_LC_12_14_1.LUT_INIT=16'b1111101000010001;
    LogicCell40 eis_state_i0_LC_12_14_1 (
            .in0(N__36416),
            .in1(N__36724),
            .in2(N__32309),
            .in3(N__32306),
            .lcout(eis_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__36146),
            .sr(N__36352));
    defparam eis_state_1__bdd_4_lut_LC_12_14_2.C_ON=1'b0;
    defparam eis_state_1__bdd_4_lut_LC_12_14_2.SEQ_MODE=4'b0000;
    defparam eis_state_1__bdd_4_lut_LC_12_14_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 eis_state_1__bdd_4_lut_LC_12_14_2 (
            .in0(N__35885),
            .in1(N__36415),
            .in2(N__35897),
            .in3(N__41021),
            .lcout(n22196),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_197_LC_12_14_4.C_ON=1'b0;
    defparam i1_2_lut_adj_197_LC_12_14_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_197_LC_12_14_4.LUT_INIT=16'b1111111101010101;
    LogicCell40 i1_2_lut_adj_197_LC_12_14_4 (
            .in0(N__41625),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36190),
            .lcout(n16602),
            .ltout(n16602_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i1_LC_12_14_5.C_ON=1'b0;
    defparam eis_state_i1_LC_12_14_5.SEQ_MODE=4'b1010;
    defparam eis_state_i1_LC_12_14_5.LUT_INIT=16'b1111111100000100;
    LogicCell40 eis_state_i1_LC_12_14_5 (
            .in0(N__36417),
            .in1(N__41023),
            .in2(N__32300),
            .in3(N__35432),
            .lcout(eis_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__36146),
            .sr(N__36352));
    defparam i34_3_lut_LC_12_14_7.C_ON=1'b0;
    defparam i34_3_lut_LC_12_14_7.SEQ_MODE=4'b0000;
    defparam i34_3_lut_LC_12_14_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i34_3_lut_LC_12_14_7 (
            .in0(N__36414),
            .in1(N__41433),
            .in2(_gnd_net_),
            .in3(N__32297),
            .lcout(n13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_168_LC_12_15_0.C_ON=1'b0;
    defparam i5_4_lut_adj_168_LC_12_15_0.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_168_LC_12_15_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i5_4_lut_adj_168_LC_12_15_0 (
            .in0(N__32447),
            .in1(N__32483),
            .in2(N__38995),
            .in3(N__32337),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i0_LC_12_15_1.C_ON=1'b0;
    defparam acadc_skipCount_i0_LC_12_15_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i0_LC_12_15_1.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i0_LC_12_15_1 (
            .in0(N__41284),
            .in1(N__49691),
            .in2(N__41167),
            .in3(N__49371),
            .lcout(acadc_skipCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57880),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i12_LC_12_15_2.C_ON=1'b0;
    defparam acadc_skipCount_i12_LC_12_15_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i12_LC_12_15_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i12_LC_12_15_2 (
            .in0(N__49368),
            .in1(N__44155),
            .in2(N__49775),
            .in3(N__38994),
            .lcout(acadc_skipCount_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57880),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_12_15_3.C_ON=1'b0;
    defparam i7_4_lut_LC_12_15_3.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_12_15_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_LC_12_15_3 (
            .in0(N__32426),
            .in1(N__32465),
            .in2(N__42438),
            .in3(N__32361),
            .lcout(n23_adj_1624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i10_LC_12_15_4.C_ON=1'b0;
    defparam acadc_skipCount_i10_LC_12_15_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i10_LC_12_15_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i10_LC_12_15_4 (
            .in0(N__49367),
            .in1(N__42987),
            .in2(N__49774),
            .in3(N__32338),
            .lcout(acadc_skipCount_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57880),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i11_LC_12_15_5.C_ON=1'b0;
    defparam acadc_skipCount_i11_LC_12_15_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i11_LC_12_15_5.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i11_LC_12_15_5 (
            .in0(N__44308),
            .in1(N__49369),
            .in2(N__42439),
            .in3(N__49698),
            .lcout(acadc_skipCount_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57880),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_176_LC_12_15_6.C_ON=1'b0;
    defparam i1_4_lut_adj_176_LC_12_15_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_176_LC_12_15_6.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_176_LC_12_15_6 (
            .in0(N__38014),
            .in1(N__32320),
            .in2(N__32393),
            .in3(N__41283),
            .lcout(n17_adj_1612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i5_LC_12_15_7.C_ON=1'b0;
    defparam acadc_skipCount_i5_LC_12_15_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i5_LC_12_15_7.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i5_LC_12_15_7 (
            .in0(N__45911),
            .in1(N__49370),
            .in2(N__43528),
            .in3(N__49699),
            .lcout(acadc_skipCount_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57880),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i0_LC_12_16_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i0_LC_12_16_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i0_LC_12_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i0_LC_12_16_0 (
            .in0(_gnd_net_),
            .in1(N__41432),
            .in2(N__32324),
            .in3(_gnd_net_),
            .lcout(acadc_skipcnt_0),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(n19369),
            .clk(INVacadc_skipcnt_i0_i0C_net),
            .ce(N__36627),
            .sr(N__36446));
    defparam add_79_2_THRU_CRY_0_LC_12_16_1.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_0_LC_12_16_1.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_0_LC_12_16_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_0_LC_12_16_1 (
            .in0(_gnd_net_),
            .in1(N__57410),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369),
            .carryout(n19369_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_79_2_THRU_CRY_1_LC_12_16_2.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_1_LC_12_16_2.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_1_LC_12_16_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_1_LC_12_16_2 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__57423),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369_THRU_CRY_0_THRU_CO),
            .carryout(n19369_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_79_2_THRU_CRY_2_LC_12_16_3.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_2_LC_12_16_3.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_2_LC_12_16_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_2_LC_12_16_3 (
            .in0(_gnd_net_),
            .in1(N__57414),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369_THRU_CRY_1_THRU_CO),
            .carryout(n19369_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_79_2_THRU_CRY_3_LC_12_16_4.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_3_LC_12_16_4.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_3_LC_12_16_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_3_LC_12_16_4 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__57424),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369_THRU_CRY_2_THRU_CO),
            .carryout(n19369_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_79_2_THRU_CRY_4_LC_12_16_5.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_4_LC_12_16_5.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_4_LC_12_16_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_4_LC_12_16_5 (
            .in0(_gnd_net_),
            .in1(N__57418),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369_THRU_CRY_3_THRU_CO),
            .carryout(n19369_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_79_2_THRU_CRY_5_LC_12_16_6.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_5_LC_12_16_6.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_5_LC_12_16_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_5_LC_12_16_6 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__57425),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369_THRU_CRY_4_THRU_CO),
            .carryout(n19369_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_79_2_THRU_CRY_6_LC_12_16_7.C_ON=1'b1;
    defparam add_79_2_THRU_CRY_6_LC_12_16_7.SEQ_MODE=4'b0000;
    defparam add_79_2_THRU_CRY_6_LC_12_16_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_79_2_THRU_CRY_6_LC_12_16_7 (
            .in0(_gnd_net_),
            .in1(N__57422),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19369_THRU_CRY_5_THRU_CO),
            .carryout(n19369_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i1_LC_12_17_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i1_LC_12_17_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i1_LC_12_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i1_LC_12_17_0 (
            .in0(_gnd_net_),
            .in1(N__38809),
            .in2(_gnd_net_),
            .in3(N__32408),
            .lcout(acadc_skipcnt_1),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(n19370),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i2_LC_12_17_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i2_LC_12_17_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i2_LC_12_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i2_LC_12_17_1 (
            .in0(_gnd_net_),
            .in1(N__39235),
            .in2(_gnd_net_),
            .in3(N__32405),
            .lcout(acadc_skipcnt_2),
            .ltout(),
            .carryin(n19370),
            .carryout(n19371),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i3_LC_12_17_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i3_LC_12_17_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i3_LC_12_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i3_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(N__36235),
            .in2(_gnd_net_),
            .in3(N__32402),
            .lcout(acadc_skipcnt_3),
            .ltout(),
            .carryin(n19371),
            .carryout(n19372),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i4_LC_12_17_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i4_LC_12_17_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i4_LC_12_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i4_LC_12_17_3 (
            .in0(_gnd_net_),
            .in1(N__38788),
            .in2(_gnd_net_),
            .in3(N__32399),
            .lcout(acadc_skipcnt_4),
            .ltout(),
            .carryin(n19372),
            .carryout(n19373),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i5_LC_12_17_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i5_LC_12_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i5_LC_12_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i5_LC_12_17_4 (
            .in0(_gnd_net_),
            .in1(N__36253),
            .in2(_gnd_net_),
            .in3(N__32396),
            .lcout(acadc_skipcnt_5),
            .ltout(),
            .carryin(n19373),
            .carryout(n19374),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i6_LC_12_17_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i6_LC_12_17_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i6_LC_12_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i6_LC_12_17_5 (
            .in0(_gnd_net_),
            .in1(N__32389),
            .in2(_gnd_net_),
            .in3(N__32375),
            .lcout(acadc_skipcnt_6),
            .ltout(),
            .carryin(n19374),
            .carryout(n19375),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i7_LC_12_17_6.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i7_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i7_LC_12_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i7_LC_12_17_6 (
            .in0(_gnd_net_),
            .in1(N__39253),
            .in2(_gnd_net_),
            .in3(N__32492),
            .lcout(acadc_skipcnt_7),
            .ltout(),
            .carryin(n19375),
            .carryout(n19376),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i8_LC_12_17_7.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i8_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i8_LC_12_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i8_LC_12_17_7 (
            .in0(_gnd_net_),
            .in1(N__36217),
            .in2(_gnd_net_),
            .in3(N__32489),
            .lcout(acadc_skipcnt_8),
            .ltout(),
            .carryin(n19376),
            .carryout(n19377),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__36635),
            .sr(N__36598));
    defparam acadc_skipcnt_i0_i9_LC_12_18_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i9_LC_12_18_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i9_LC_12_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i9_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(N__36481),
            .in2(_gnd_net_),
            .in3(N__32486),
            .lcout(acadc_skipcnt_9),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(n19378),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam acadc_skipcnt_i0_i10_LC_12_18_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i10_LC_12_18_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i10_LC_12_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i10_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(N__32482),
            .in2(_gnd_net_),
            .in3(N__32468),
            .lcout(acadc_skipcnt_10),
            .ltout(),
            .carryin(n19378),
            .carryout(n19379),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam acadc_skipcnt_i0_i11_LC_12_18_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i11_LC_12_18_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i11_LC_12_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i11_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(N__32464),
            .in2(_gnd_net_),
            .in3(N__32450),
            .lcout(acadc_skipcnt_11),
            .ltout(),
            .carryin(n19379),
            .carryout(n19380),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam acadc_skipcnt_i0_i12_LC_12_18_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i12_LC_12_18_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i12_LC_12_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i12_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(N__32446),
            .in2(_gnd_net_),
            .in3(N__32432),
            .lcout(acadc_skipcnt_12),
            .ltout(),
            .carryin(n19380),
            .carryout(n19381),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam acadc_skipcnt_i0_i13_LC_12_18_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i13_LC_12_18_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i13_LC_12_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i13_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(N__38857),
            .in2(_gnd_net_),
            .in3(N__32429),
            .lcout(acadc_skipcnt_13),
            .ltout(),
            .carryin(n19381),
            .carryout(n19382),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam acadc_skipcnt_i0_i14_LC_12_18_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i14_LC_12_18_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i14_LC_12_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i14_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(N__32425),
            .in2(_gnd_net_),
            .in3(N__32411),
            .lcout(acadc_skipcnt_14),
            .ltout(),
            .carryin(n19382),
            .carryout(n19383),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam acadc_skipcnt_i0_i15_LC_12_18_6.C_ON=1'b0;
    defparam acadc_skipcnt_i0_i15_LC_12_18_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i15_LC_12_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i15_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(N__36496),
            .in2(_gnd_net_),
            .in3(N__32744),
            .lcout(acadc_skipcnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__36634),
            .sr(N__36599));
    defparam SecClk_302_LC_12_19_7.C_ON=1'b0;
    defparam SecClk_302_LC_12_19_7.SEQ_MODE=4'b1000;
    defparam SecClk_302_LC_12_19_7.LUT_INIT=16'b0101010110101010;
    LogicCell40 SecClk_302_LC_12_19_7 (
            .in0(N__32714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39746),
            .lcout(TEST_LED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45081),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_LC_13_3_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_13_3_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_LC_13_3_0  (
            .in0(N__32689),
            .in1(N__32677),
            .in2(N__32666),
            .in3(N__32650),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i18779_4_lut_LC_13_3_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i18779_4_lut_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i18779_4_lut_LC_13_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i18779_4_lut_LC_13_3_1  (
            .in0(N__32504),
            .in1(N__32639),
            .in2(N__32630),
            .in3(N__32567),
            .lcout(\ADC_VDC.genclk.n21206 ),
            .ltout(\ADC_VDC.genclk.n21206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i0_LC_13_3_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i0_LC_13_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i0_LC_13_3_2 .LUT_INIT=16'b1111011111010101;
    LogicCell40 \ADC_VDC.genclk.div_state_i0_LC_13_3_2  (
            .in0(N__33673),
            .in1(N__40170),
            .in2(N__32627),
            .in3(N__37216),
            .lcout(\ADC_VDC.genclk.div_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19076_4_lut_LC_13_3_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19076_4_lut_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19076_4_lut_LC_13_3_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \ADC_VDC.genclk.i19076_4_lut_LC_13_3_3  (
            .in0(N__32620),
            .in1(N__32608),
            .in2(N__32596),
            .in3(N__32578),
            .lcout(\ADC_VDC.genclk.n21208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_LC_13_3_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_13_3_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_LC_13_3_4  (
            .in0(N__32560),
            .in1(N__32545),
            .in2(N__32534),
            .in3(N__32515),
            .lcout(\ADC_VDC.genclk.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19182_2_lut_4_lut_LC_13_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19182_2_lut_4_lut_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19182_2_lut_4_lut_LC_13_4_0 .LUT_INIT=16'b0010011111111111;
    LogicCell40 \ADC_VDC.genclk.i19182_2_lut_4_lut_LC_13_4_0  (
            .in0(N__40162),
            .in1(N__32498),
            .in2(N__37217),
            .in3(N__33668),
            .lcout(\ADC_VDC.genclk.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i1_LC_13_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i1_LC_13_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i1_LC_13_4_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ADC_VDC.genclk.div_state_i1_LC_13_4_1  (
            .in0(N__33669),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40163),
            .lcout(\ADC_VDC.genclk.div_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i1C_net ),
            .ce(N__33686),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12662_2_lut_2_lut_LC_13_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12662_2_lut_2_lut_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12662_2_lut_2_lut_LC_13_4_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \ADC_VDC.genclk.i12662_2_lut_2_lut_LC_13_4_2  (
            .in0(N__40160),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33667),
            .lcout(\ADC_VDC.genclk.n15067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_4_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_4_4  (
            .in0(N__40161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.genclk.div_state_1__N_1275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16075_4_lut_LC_13_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i16075_4_lut_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16075_4_lut_LC_13_4_5 .LUT_INIT=16'b1001100010111010;
    LogicCell40 \ADC_VDC.i16075_4_lut_LC_13_4_5  (
            .in0(N__33300),
            .in1(N__33097),
            .in2(N__33383),
            .in3(N__32895),
            .lcout(\ADC_VDC.n11766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_39_LC_13_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_39_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_39_LC_13_4_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_39_LC_13_4_6  (
            .in0(N__33630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33524),
            .lcout(\ADC_VDC.n62 ),
            .ltout(\ADC_VDC.n62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i24_4_lut_LC_13_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i24_4_lut_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i24_4_lut_LC_13_4_7 .LUT_INIT=16'b1001100010111010;
    LogicCell40 \ADC_VDC.i24_4_lut_LC_13_4_7  (
            .in0(N__33299),
            .in1(N__33096),
            .in2(N__32909),
            .in3(N__32894),
            .lcout(\ADC_VDC.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0on_i0_LC_13_5_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i0_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i0_LC_13_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i0_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__37232),
            .in2(_gnd_net_),
            .in3(N__32753),
            .lcout(\ADC_VDC.genclk.t0on_0 ),
            .ltout(),
            .carryin(bfn_13_5_0_),
            .carryout(\ADC_VDC.genclk.n19483 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i1_LC_13_5_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i1_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i1_LC_13_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i1_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(N__37265),
            .in2(N__57388),
            .in3(N__32750),
            .lcout(\ADC_VDC.genclk.t0on_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19483 ),
            .carryout(\ADC_VDC.genclk.n19484 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i2_LC_13_5_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i2_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i2_LC_13_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i2_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(N__57353),
            .in2(N__37064),
            .in3(N__32747),
            .lcout(\ADC_VDC.genclk.t0on_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19484 ),
            .carryout(\ADC_VDC.genclk.n19485 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i3_LC_13_5_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i3_LC_13_5_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0on_i3_LC_13_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i3_LC_13_5_3  (
            .in0(_gnd_net_),
            .in1(N__37187),
            .in2(N__57389),
            .in3(N__33713),
            .lcout(\ADC_VDC.genclk.t0on_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19485 ),
            .carryout(\ADC_VDC.genclk.n19486 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i4_LC_13_5_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i4_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i4_LC_13_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i4_LC_13_5_4  (
            .in0(_gnd_net_),
            .in1(N__57357),
            .in2(N__37252),
            .in3(N__33710),
            .lcout(\ADC_VDC.genclk.t0on_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19486 ),
            .carryout(\ADC_VDC.genclk.n19487 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i5_LC_13_5_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i5_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i5_LC_13_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i5_LC_13_5_5  (
            .in0(_gnd_net_),
            .in1(N__37174),
            .in2(N__57390),
            .in3(N__33707),
            .lcout(\ADC_VDC.genclk.t0on_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19487 ),
            .carryout(\ADC_VDC.genclk.n19488 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i6_LC_13_5_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i6_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i6_LC_13_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i6_LC_13_5_6  (
            .in0(_gnd_net_),
            .in1(N__57361),
            .in2(N__37280),
            .in3(N__33704),
            .lcout(\ADC_VDC.genclk.t0on_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19488 ),
            .carryout(\ADC_VDC.genclk.n19489 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i7_LC_13_5_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i7_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i7_LC_13_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i7_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__37048),
            .in2(N__57391),
            .in3(N__33701),
            .lcout(\ADC_VDC.genclk.t0on_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19489 ),
            .carryout(\ADC_VDC.genclk.n19490 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__33908),
            .sr(N__33881));
    defparam \ADC_VDC.genclk.t0on_i8_LC_13_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i8_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i8_LC_13_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i8_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__57375),
            .in2(N__37160),
            .in3(N__33698),
            .lcout(\ADC_VDC.genclk.t0on_8 ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\ADC_VDC.genclk.n19491 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i9_LC_13_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i9_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i9_LC_13_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i9_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__37124),
            .in2(N__57394),
            .in3(N__33695),
            .lcout(\ADC_VDC.genclk.t0on_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19491 ),
            .carryout(\ADC_VDC.genclk.n19492 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i10_LC_13_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i10_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i10_LC_13_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i10_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__57365),
            .in2(N__37034),
            .in3(N__33692),
            .lcout(\ADC_VDC.genclk.t0on_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19492 ),
            .carryout(\ADC_VDC.genclk.n19493 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i11_LC_13_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i11_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i11_LC_13_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i11_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__37097),
            .in2(N__57392),
            .in3(N__33689),
            .lcout(\ADC_VDC.genclk.t0on_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19493 ),
            .carryout(\ADC_VDC.genclk.n19494 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i12_LC_13_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i12_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i12_LC_13_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i12_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__57369),
            .in2(N__37079),
            .in3(N__33920),
            .lcout(\ADC_VDC.genclk.t0on_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19494 ),
            .carryout(\ADC_VDC.genclk.n19495 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i13_LC_13_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i13_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i13_LC_13_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i13_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__37199),
            .in2(N__57393),
            .in3(N__33917),
            .lcout(\ADC_VDC.genclk.t0on_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19495 ),
            .carryout(\ADC_VDC.genclk.n19496 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i14_LC_13_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i14_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i14_LC_13_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i14_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__57373),
            .in2(N__37139),
            .in3(N__33914),
            .lcout(\ADC_VDC.genclk.t0on_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19496 ),
            .carryout(\ADC_VDC.genclk.n19497 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \ADC_VDC.genclk.t0on_i15_LC_13_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0on_i15_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i15_LC_13_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0on_i15_LC_13_6_7  (
            .in0(N__57374),
            .in1(N__37111),
            .in2(_gnd_net_),
            .in3(N__33911),
            .lcout(\ADC_VDC.genclk.t0on_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__33907),
            .sr(N__33873));
    defparam \RTD.bit_cnt_3782__i3_LC_13_7_0 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3782__i3_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3782__i3_LC_13_7_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \RTD.bit_cnt_3782__i3_LC_13_7_0  (
            .in0(N__33809),
            .in1(N__33823),
            .in2(N__33776),
            .in3(N__33791),
            .lcout(\RTD.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43735),
            .ce(N__33749),
            .sr(N__33731));
    defparam \RTD.bit_cnt_3782__i1_LC_13_7_1 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3782__i1_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3782__i1_LC_13_7_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RTD.bit_cnt_3782__i1_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__33768),
            .in2(_gnd_net_),
            .in3(N__33807),
            .lcout(\RTD.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43735),
            .ce(N__33749),
            .sr(N__33731));
    defparam \RTD.bit_cnt_3782__i2_LC_13_7_2 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3782__i2_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3782__i2_LC_13_7_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \RTD.bit_cnt_3782__i2_LC_13_7_2  (
            .in0(N__33808),
            .in1(_gnd_net_),
            .in2(N__33775),
            .in3(N__33790),
            .lcout(\RTD.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43735),
            .ce(N__33749),
            .sr(N__33731));
    defparam \RTD.bit_cnt_3782__i0_LC_13_7_3 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3782__i0_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3782__i0_LC_13_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \RTD.bit_cnt_3782__i0_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33767),
            .lcout(\RTD.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__43735),
            .ce(N__33749),
            .sr(N__33731));
    defparam i1_3_lut_adj_245_LC_13_7_4.C_ON=1'b0;
    defparam i1_3_lut_adj_245_LC_13_7_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_245_LC_13_7_4.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_3_lut_adj_245_LC_13_7_4 (
            .in0(N__42783),
            .in1(N__50931),
            .in2(_gnd_net_),
            .in3(N__37478),
            .lcout(n12152),
            .ltout(n12152_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12374_2_lut_LC_13_7_5.C_ON=1'b0;
    defparam i12374_2_lut_LC_13_7_5.SEQ_MODE=4'b0000;
    defparam i12374_2_lut_LC_13_7_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12374_2_lut_LC_13_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34085),
            .in3(N__54829),
            .lcout(n14787),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_247_LC_13_7_6.C_ON=1'b0;
    defparam i1_3_lut_adj_247_LC_13_7_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_247_LC_13_7_6.LUT_INIT=16'b1010101010100000;
    LogicCell40 i1_3_lut_adj_247_LC_13_7_6 (
            .in0(N__42784),
            .in1(_gnd_net_),
            .in2(N__34082),
            .in3(N__50930),
            .lcout(n12194),
            .ltout(n12194_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12381_2_lut_LC_13_7_7.C_ON=1'b0;
    defparam i12381_2_lut_LC_13_7_7.SEQ_MODE=4'b0000;
    defparam i12381_2_lut_LC_13_7_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12381_2_lut_LC_13_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34073),
            .in3(N__54828),
            .lcout(n14794),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_0_i22_3_lut_LC_13_8_0.C_ON=1'b0;
    defparam mux_136_Mux_0_i22_3_lut_LC_13_8_0.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_0_i22_3_lut_LC_13_8_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_136_Mux_0_i22_3_lut_LC_13_8_0 (
            .in0(N__34063),
            .in1(N__33926),
            .in2(_gnd_net_),
            .in3(N__49074),
            .lcout(),
            .ltout(n22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_136_Mux_0_i30_3_lut_LC_13_8_1.C_ON=1'b0;
    defparam mux_136_Mux_0_i30_3_lut_LC_13_8_1.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_0_i30_3_lut_LC_13_8_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_136_Mux_0_i30_3_lut_LC_13_8_1 (
            .in0(N__48738),
            .in1(_gnd_net_),
            .in2(N__34037),
            .in3(N__34034),
            .lcout(),
            .ltout(n30_adj_1484_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i0_LC_13_8_2.C_ON=1'b0;
    defparam comm_buf_2__i0_LC_13_8_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i0_LC_13_8_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_2__i0_LC_13_8_2 (
            .in0(_gnd_net_),
            .in1(N__50778),
            .in2(N__34022),
            .in3(N__53842),
            .lcout(comm_buf_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57823),
            .ce(N__34216),
            .sr(N__34189));
    defparam mux_136_Mux_1_i30_3_lut_LC_13_8_3.C_ON=1'b0;
    defparam mux_136_Mux_1_i30_3_lut_LC_13_8_3.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_1_i30_3_lut_LC_13_8_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_136_Mux_1_i30_3_lut_LC_13_8_3 (
            .in0(N__48739),
            .in1(_gnd_net_),
            .in2(N__34019),
            .in3(N__34004),
            .lcout(),
            .ltout(n30_adj_1504_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i1_LC_13_8_4.C_ON=1'b0;
    defparam comm_buf_2__i1_LC_13_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i1_LC_13_8_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_2__i1_LC_13_8_4 (
            .in0(N__45364),
            .in1(_gnd_net_),
            .in2(N__33989),
            .in3(N__53843),
            .lcout(comm_buf_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57823),
            .ce(N__34216),
            .sr(N__34189));
    defparam mux_136_Mux_0_i19_3_lut_LC_13_8_5.C_ON=1'b0;
    defparam mux_136_Mux_0_i19_3_lut_LC_13_8_5.SEQ_MODE=4'b0000;
    defparam mux_136_Mux_0_i19_3_lut_LC_13_8_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_136_Mux_0_i19_3_lut_LC_13_8_5 (
            .in0(N__33986),
            .in1(N__33965),
            .in2(_gnd_net_),
            .in3(N__56143),
            .lcout(n19_adj_1485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_242_LC_13_8_6.C_ON=1'b0;
    defparam i1_4_lut_adj_242_LC_13_8_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_242_LC_13_8_6.LUT_INIT=16'b1100010011000000;
    LogicCell40 i1_4_lut_adj_242_LC_13_8_6 (
            .in0(N__53566),
            .in1(N__42782),
            .in2(N__50933),
            .in3(N__37793),
            .lcout(n12110),
            .ltout(n12110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12367_2_lut_LC_13_8_7.C_ON=1'b0;
    defparam i12367_2_lut_LC_13_8_7.SEQ_MODE=4'b0000;
    defparam i12367_2_lut_LC_13_8_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12367_2_lut_LC_13_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34193),
            .in3(N__54735),
            .lcout(n14780),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18291_3_lut_LC_13_9_0.C_ON=1'b0;
    defparam i18291_3_lut_LC_13_9_0.SEQ_MODE=4'b0000;
    defparam i18291_3_lut_LC_13_9_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18291_3_lut_LC_13_9_0 (
            .in0(N__55948),
            .in1(N__34166),
            .in2(_gnd_net_),
            .in3(N__42068),
            .lcout(),
            .ltout(n20905_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19514_LC_13_9_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19514_LC_13_9_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19514_LC_13_9_1.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19514_LC_13_9_1 (
            .in0(N__48217),
            .in1(N__34091),
            .in2(N__34145),
            .in3(N__48875),
            .lcout(),
            .ltout(n22148_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22148_bdd_4_lut_LC_13_9_2.C_ON=1'b0;
    defparam n22148_bdd_4_lut_LC_13_9_2.SEQ_MODE=4'b0000;
    defparam n22148_bdd_4_lut_LC_13_9_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22148_bdd_4_lut_LC_13_9_2 (
            .in0(N__48876),
            .in1(N__34142),
            .in2(N__34127),
            .in3(N__34715),
            .lcout(),
            .ltout(n22151_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18275_3_lut_LC_13_9_3.C_ON=1'b0;
    defparam i18275_3_lut_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam i18275_3_lut_LC_13_9_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i18275_3_lut_LC_13_9_3 (
            .in0(_gnd_net_),
            .in1(N__34124),
            .in2(N__34112),
            .in3(N__48619),
            .lcout(),
            .ltout(n20889_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i2_LC_13_9_4.C_ON=1'b0;
    defparam comm_buf_0__i2_LC_13_9_4.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i2_LC_13_9_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_0__i2_LC_13_9_4 (
            .in0(_gnd_net_),
            .in1(N__47247),
            .in2(N__34109),
            .in3(N__54089),
            .lcout(comm_buf_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57832),
            .ce(N__42725),
            .sr(N__42856));
    defparam i18735_2_lut_LC_13_9_5.C_ON=1'b0;
    defparam i18735_2_lut_LC_13_9_5.SEQ_MODE=4'b0000;
    defparam i18735_2_lut_LC_13_9_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18735_2_lut_LC_13_9_5 (
            .in0(_gnd_net_),
            .in1(N__34106),
            .in2(_gnd_net_),
            .in3(N__55947),
            .lcout(n20906),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_i8_2_lut_LC_13_9_6.C_ON=1'b0;
    defparam comm_cmd_6__I_0_i8_2_lut_LC_13_9_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_i8_2_lut_LC_13_9_6.LUT_INIT=16'b1010101011111111;
    LogicCell40 comm_cmd_6__I_0_i8_2_lut_LC_13_9_6 (
            .in0(N__48874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48216),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_278_LC_13_9_7.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_278_LC_13_9_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_278_LC_13_9_7.LUT_INIT=16'b1111111111111011;
    LogicCell40 i1_2_lut_4_lut_adj_278_LC_13_9_7 (
            .in0(N__48215),
            .in1(N__55946),
            .in2(N__34838),
            .in3(N__48873),
            .lcout(n20672),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i1_LC_13_10_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i1_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i1_LC_13_10_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i1_LC_13_10_0  (
            .in0(N__34650),
            .in1(N__35404),
            .in2(N__34772),
            .in3(N__34734),
            .lcout(buf_adcdata_vac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57842),
            .ce(),
            .sr(_gnd_net_));
    defparam i18226_3_lut_LC_13_10_1.C_ON=1'b0;
    defparam i18226_3_lut_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam i18226_3_lut_LC_13_10_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18226_3_lut_LC_13_10_1 (
            .in0(N__55945),
            .in1(N__35678),
            .in2(_gnd_net_),
            .in3(N__42017),
            .lcout(n20840),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i13_LC_13_10_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i13_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i13_LC_13_10_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i13_LC_13_10_2  (
            .in0(N__34649),
            .in1(N__35403),
            .in2(N__34706),
            .in3(N__46635),
            .lcout(buf_adcdata_vac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57842),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i12_LC_13_10_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i12_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i12_LC_13_10_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i12_LC_13_10_3  (
            .in0(N__35400),
            .in1(N__34651),
            .in2(N__34688),
            .in3(N__35593),
            .lcout(buf_adcdata_vac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57842),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i11_LC_13_10_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i11_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i11_LC_13_10_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i11_LC_13_10_4  (
            .in0(N__34648),
            .in1(N__35402),
            .in2(N__38290),
            .in3(N__34520),
            .lcout(buf_adcdata_vac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57842),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_13_10_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_13_10_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i26_LC_13_10_5  (
            .in0(N__35401),
            .in1(N__34483),
            .in2(N__34234),
            .in3(N__34429),
            .lcout(cmd_rdadctmp_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57842),
            .ce(),
            .sr(_gnd_net_));
    defparam i39_3_lut_LC_13_10_6.C_ON=1'b0;
    defparam i39_3_lut_LC_13_10_6.SEQ_MODE=4'b0000;
    defparam i39_3_lut_LC_13_10_6.LUT_INIT=16'b0101010110001000;
    LogicCell40 i39_3_lut_LC_13_10_6 (
            .in0(N__48090),
            .in1(N__55944),
            .in2(_gnd_net_),
            .in3(N__48856),
            .lcout(),
            .ltout(n24_adj_1622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i41_3_lut_LC_13_10_7.C_ON=1'b0;
    defparam i41_3_lut_LC_13_10_7.SEQ_MODE=4'b0000;
    defparam i41_3_lut_LC_13_10_7.LUT_INIT=16'b0011000011111100;
    LogicCell40 i41_3_lut_LC_13_10_7 (
            .in0(_gnd_net_),
            .in1(N__48703),
            .in2(N__35630),
            .in3(N__36572),
            .lcout(n21_adj_1618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_4_i19_3_lut_LC_13_11_0.C_ON=1'b0;
    defparam mux_135_Mux_4_i19_3_lut_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_4_i19_3_lut_LC_13_11_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_4_i19_3_lut_LC_13_11_0 (
            .in0(N__35627),
            .in1(N__35589),
            .in2(_gnd_net_),
            .in3(N__55949),
            .lcout(n19_adj_1509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_214_LC_13_11_1.C_ON=1'b0;
    defparam i1_2_lut_adj_214_LC_13_11_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_214_LC_13_11_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_214_LC_13_11_1 (
            .in0(_gnd_net_),
            .in1(N__41051),
            .in2(_gnd_net_),
            .in3(N__36432),
            .lcout(),
            .ltout(n35_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3798_3_lut_3_lut_4_lut_LC_13_11_2.C_ON=1'b0;
    defparam i3798_3_lut_3_lut_4_lut_LC_13_11_2.SEQ_MODE=4'b0000;
    defparam i3798_3_lut_3_lut_4_lut_LC_13_11_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 i3798_3_lut_3_lut_4_lut_LC_13_11_2 (
            .in0(N__41418),
            .in1(N__36719),
            .in2(N__35573),
            .in3(N__36337),
            .lcout(iac_raw_buf_N_735),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_13_11_3.C_ON=1'b0;
    defparam i24_4_lut_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_13_11_3.LUT_INIT=16'b0111101001011000;
    LogicCell40 i24_4_lut_LC_13_11_3 (
            .in0(N__36720),
            .in1(N__41052),
            .in2(N__36437),
            .in3(N__41419),
            .lcout(n17_adj_1645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.DTRIG_39_LC_13_11_4 .C_ON=1'b0;
    defparam \ADC_VAC.DTRIG_39_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.DTRIG_39_LC_13_11_4 .LUT_INIT=16'b1111111001000000;
    LogicCell40 \ADC_VAC.DTRIG_39_LC_13_11_4  (
            .in0(N__35416),
            .in1(N__35048),
            .in2(N__34967),
            .in3(N__36118),
            .lcout(acadc_dtrig_v),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57852),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_start_340_LC_13_11_5.C_ON=1'b0;
    defparam eis_start_340_LC_13_11_5.SEQ_MODE=4'b1000;
    defparam eis_start_340_LC_13_11_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 eis_start_340_LC_13_11_5 (
            .in0(N__41623),
            .in1(N__43878),
            .in2(_gnd_net_),
            .in3(N__41493),
            .lcout(eis_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57852),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_13_11_6.C_ON=1'b0;
    defparam i2_4_lut_LC_13_11_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_13_11_6.LUT_INIT=16'b0000000000000010;
    LogicCell40 i2_4_lut_LC_13_11_6 (
            .in0(N__54823),
            .in1(N__53567),
            .in2(N__34877),
            .in3(N__34865),
            .lcout(n10534),
            .ltout(n10534_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam auxmode_337_LC_13_11_7.C_ON=1'b0;
    defparam auxmode_337_LC_13_11_7.SEQ_MODE=4'b1000;
    defparam auxmode_337_LC_13_11_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 auxmode_337_LC_13_11_7 (
            .in0(N__44281),
            .in1(_gnd_net_),
            .in2(N__34841),
            .in3(N__35698),
            .lcout(auxmode),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57852),
            .ce(),
            .sr(_gnd_net_));
    defparam i14180_1_lut_2_lut_3_lut_LC_13_12_0.C_ON=1'b0;
    defparam i14180_1_lut_2_lut_3_lut_LC_13_12_0.SEQ_MODE=4'b0000;
    defparam i14180_1_lut_2_lut_3_lut_LC_13_12_0.LUT_INIT=16'b1111111101011111;
    LogicCell40 i14180_1_lut_2_lut_3_lut_LC_13_12_0 (
            .in0(N__36085),
            .in1(_gnd_net_),
            .in2(N__36122),
            .in3(N__36675),
            .lcout(n16598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_LC_13_12_1 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_LC_13_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VAC.i1_2_lut_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__36111),
            .in2(_gnd_net_),
            .in3(N__36083),
            .lcout(iac_raw_buf_N_737),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18743_2_lut_3_lut_LC_13_12_2.C_ON=1'b0;
    defparam i18743_2_lut_3_lut_LC_13_12_2.SEQ_MODE=4'b0000;
    defparam i18743_2_lut_3_lut_LC_13_12_2.LUT_INIT=16'b0101111100000000;
    LogicCell40 i18743_2_lut_3_lut_LC_13_12_2 (
            .in0(N__36084),
            .in1(_gnd_net_),
            .in2(N__36121),
            .in3(N__36676),
            .lcout(n20957),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.DTRIG_39_LC_13_12_3 .C_ON=1'b0;
    defparam \ADC_IAC.DTRIG_39_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.DTRIG_39_LC_13_12_3 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \ADC_IAC.DTRIG_39_LC_13_12_3  (
            .in0(N__35876),
            .in1(N__35804),
            .in2(N__53001),
            .in3(N__36086),
            .lcout(acadc_dtrig_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57862),
            .ce(),
            .sr(_gnd_net_));
    defparam ICE_GPMO_0_I_0_3_lut_LC_13_12_4.C_ON=1'b0;
    defparam ICE_GPMO_0_I_0_3_lut_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam ICE_GPMO_0_I_0_3_lut_LC_13_12_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 ICE_GPMO_0_I_0_3_lut_LC_13_12_4 (
            .in0(N__35741),
            .in1(N__35697),
            .in2(_gnd_net_),
            .in3(N__35673),
            .lcout(acadc_rst),
            .ltout(acadc_rst_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_4_lut_LC_13_12_5.C_ON=1'b0;
    defparam i2_4_lut_4_lut_4_lut_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_4_lut_LC_13_12_5.LUT_INIT=16'b0000010100000001;
    LogicCell40 i2_4_lut_4_lut_4_lut_LC_13_12_5 (
            .in0(N__36674),
            .in1(N__41045),
            .in2(N__35681),
            .in3(N__36421),
            .lcout(n13473),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam tacadc_rst_338_LC_13_12_6.C_ON=1'b0;
    defparam tacadc_rst_338_LC_13_12_6.SEQ_MODE=4'b1000;
    defparam tacadc_rst_338_LC_13_12_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 tacadc_rst_338_LC_13_12_6 (
            .in0(N__42970),
            .in1(N__43879),
            .in2(_gnd_net_),
            .in3(N__35674),
            .lcout(tacadc_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57862),
            .ce(),
            .sr(_gnd_net_));
    defparam i18184_3_lut_LC_13_12_7.C_ON=1'b0;
    defparam i18184_3_lut_LC_13_12_7.SEQ_MODE=4'b0000;
    defparam i18184_3_lut_LC_13_12_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18184_3_lut_LC_13_12_7 (
            .in0(N__35660),
            .in1(N__35642),
            .in2(_gnd_net_),
            .in3(N__48335),
            .lcout(n20798),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_201_LC_13_13_0.C_ON=1'b0;
    defparam i24_4_lut_adj_201_LC_13_13_0.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_201_LC_13_13_0.LUT_INIT=16'b1111110010101100;
    LogicCell40 i24_4_lut_adj_201_LC_13_13_0 (
            .in0(N__41624),
            .in1(N__36128),
            .in2(N__36431),
            .in3(N__44905),
            .lcout(),
            .ltout(n11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19147_3_lut_LC_13_13_1.C_ON=1'b0;
    defparam i19147_3_lut_LC_13_13_1.SEQ_MODE=4'b0000;
    defparam i19147_3_lut_LC_13_13_1.LUT_INIT=16'b0011111111111111;
    LogicCell40 i19147_3_lut_LC_13_13_1 (
            .in0(_gnd_net_),
            .in1(N__41020),
            .in2(N__36158),
            .in3(N__36685),
            .lcout(n11760),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18865_2_lut_LC_13_13_2.C_ON=1'b0;
    defparam i18865_2_lut_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam i18865_2_lut_LC_13_13_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i18865_2_lut_LC_13_13_2 (
            .in0(N__43920),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36420),
            .lcout(),
            .ltout(n21099_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i2_LC_13_13_3.C_ON=1'b0;
    defparam eis_state_i2_LC_13_13_3.SEQ_MODE=4'b1010;
    defparam eis_state_i2_LC_13_13_3.LUT_INIT=16'b1110011011000100;
    LogicCell40 eis_state_i2_LC_13_13_3 (
            .in0(N__41022),
            .in1(N__36686),
            .in2(N__36155),
            .in3(N__36152),
            .lcout(eis_end_N_725),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i2C_net),
            .ce(N__36142),
            .sr(N__36338));
    defparam i15032_2_lut_LC_13_13_4.C_ON=1'b0;
    defparam i15032_2_lut_LC_13_13_4.SEQ_MODE=4'b0000;
    defparam i15032_2_lut_LC_13_13_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i15032_2_lut_LC_13_13_4 (
            .in0(_gnd_net_),
            .in1(N__36119),
            .in2(_gnd_net_),
            .in3(N__36081),
            .lcout(n17430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_263_LC_13_13_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_263_LC_13_13_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_263_LC_13_13_6.LUT_INIT=16'b0000000000110000;
    LogicCell40 i1_2_lut_3_lut_adj_263_LC_13_13_6 (
            .in0(_gnd_net_),
            .in1(N__36120),
            .in2(N__43924),
            .in3(N__36082),
            .lcout(n4_adj_1569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i3_LC_13_14_0.C_ON=1'b0;
    defparam data_index_i3_LC_13_14_0.SEQ_MODE=4'b1000;
    defparam data_index_i3_LC_13_14_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i3_LC_13_14_0 (
            .in0(N__36023),
            .in1(N__54967),
            .in2(N__49780),
            .in3(N__36014),
            .lcout(data_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57885),
            .ce(),
            .sr(_gnd_net_));
    defparam i6444_3_lut_LC_13_14_1.C_ON=1'b0;
    defparam i6444_3_lut_LC_13_14_1.SEQ_MODE=4'b0000;
    defparam i6444_3_lut_LC_13_14_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 i6444_3_lut_LC_13_14_1 (
            .in0(N__41747),
            .in1(N__37970),
            .in2(_gnd_net_),
            .in3(N__36039),
            .lcout(n8_adj_1563),
            .ltout(n8_adj_1563_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_3_i15_4_lut_LC_13_14_2.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_3_i15_4_lut_LC_13_14_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_3_i15_4_lut_LC_13_14_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_365_Mux_3_i15_4_lut_LC_13_14_2 (
            .in0(N__49708),
            .in1(N__54966),
            .in2(N__36017),
            .in3(N__36013),
            .lcout(data_index_9_N_216_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i3_LC_13_14_3.C_ON=1'b0;
    defparam acadc_skipCount_i3_LC_13_14_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i3_LC_13_14_3.LUT_INIT=16'b0111001001010000;
    LogicCell40 acadc_skipCount_i3_LC_13_14_3 (
            .in0(N__49343),
            .in1(N__49709),
            .in2(N__37930),
            .in3(N__37971),
            .lcout(acadc_skipCount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57885),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i8_LC_13_14_4.C_ON=1'b0;
    defparam acadc_skipCount_i8_LC_13_14_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i8_LC_13_14_4.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i8_LC_13_14_4 (
            .in0(N__49710),
            .in1(N__49342),
            .in2(N__41656),
            .in3(N__41494),
            .lcout(acadc_skipCount_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57885),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_13_14_5.C_ON=1'b0;
    defparam i4_4_lut_LC_13_14_5.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_13_14_5.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_LC_13_14_5 (
            .in0(N__36254),
            .in1(N__36239),
            .in2(N__37929),
            .in3(N__43524),
            .lcout(),
            .ltout(n20_adj_1617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_13_14_6.C_ON=1'b0;
    defparam i10_4_lut_LC_13_14_6.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_13_14_6.LUT_INIT=16'b1111111111110110;
    LogicCell40 i10_4_lut_LC_13_14_6 (
            .in0(N__36221),
            .in1(N__41646),
            .in2(N__36203),
            .in3(N__38819),
            .lcout(),
            .ltout(n26_adj_1640_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_179_LC_13_14_7.C_ON=1'b0;
    defparam i15_4_lut_adj_179_LC_13_14_7.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_179_LC_13_14_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_179_LC_13_14_7 (
            .in0(N__38774),
            .in1(N__36200),
            .in2(N__36194),
            .in3(N__36452),
            .lcout(n31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6434_3_lut_LC_13_15_1.C_ON=1'b0;
    defparam i6434_3_lut_LC_13_15_1.SEQ_MODE=4'b0000;
    defparam i6434_3_lut_LC_13_15_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6434_3_lut_LC_13_15_1 (
            .in0(N__51168),
            .in1(N__38755),
            .in2(_gnd_net_),
            .in3(N__41729),
            .lcout(n8_adj_1561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i6_LC_13_15_2.C_ON=1'b0;
    defparam acadc_skipCount_i6_LC_13_15_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i6_LC_13_15_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 acadc_skipCount_i6_LC_13_15_2 (
            .in0(N__49357),
            .in1(N__49686),
            .in2(N__52506),
            .in3(N__38013),
            .lcout(acadc_skipCount_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57897),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i9_LC_13_15_3.C_ON=1'b0;
    defparam acadc_skipCount_i9_LC_13_15_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i9_LC_13_15_3.LUT_INIT=16'b0000110010101010;
    LogicCell40 acadc_skipCount_i9_LC_13_15_3 (
            .in0(N__44608),
            .in1(N__45556),
            .in2(N__49773),
            .in3(N__49359),
            .lcout(acadc_skipCount_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57897),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i7_LC_13_15_4.C_ON=1'b0;
    defparam acadc_skipCount_i7_LC_13_15_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i7_LC_13_15_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 acadc_skipCount_i7_LC_13_15_4 (
            .in0(N__49358),
            .in1(N__49687),
            .in2(N__47673),
            .in3(N__49176),
            .lcout(acadc_skipCount_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57897),
            .ce(),
            .sr(_gnd_net_));
    defparam i6454_3_lut_LC_13_15_5.C_ON=1'b0;
    defparam i6454_3_lut_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam i6454_3_lut_LC_13_15_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i6454_3_lut_LC_13_15_5 (
            .in0(N__36180),
            .in1(N__47139),
            .in2(_gnd_net_),
            .in3(N__41730),
            .lcout(n8_adj_1565),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_13_15_6.C_ON=1'b0;
    defparam i8_4_lut_LC_13_15_6.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_13_15_6.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_LC_13_15_6 (
            .in0(N__36500),
            .in1(N__36482),
            .in2(N__47787),
            .in3(N__44607),
            .lcout(),
            .ltout(n24_adj_1537_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_13_15_7.C_ON=1'b0;
    defparam i14_4_lut_LC_13_15_7.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_13_15_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_13_15_7 (
            .in0(N__39221),
            .in1(N__36467),
            .in2(N__36461),
            .in3(N__36458),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19175_2_lut_3_lut_LC_13_16_0.C_ON=1'b0;
    defparam i19175_2_lut_3_lut_LC_13_16_0.SEQ_MODE=4'b0000;
    defparam i19175_2_lut_3_lut_LC_13_16_0.LUT_INIT=16'b0000000000010001;
    LogicCell40 i19175_2_lut_3_lut_LC_13_16_0 (
            .in0(N__36345),
            .in1(N__41049),
            .in2(_gnd_net_),
            .in3(N__36708),
            .lcout(n20789),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i5_LC_13_16_1.C_ON=1'b0;
    defparam buf_dds1_i5_LC_13_16_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i5_LC_13_16_1.LUT_INIT=16'b1110001011101110;
    LogicCell40 buf_dds1_i5_LC_13_16_1 (
            .in0(N__36295),
            .in1(N__38567),
            .in2(N__47327),
            .in3(N__54847),
            .lcout(buf_dds1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57914),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i7_LC_13_16_3.C_ON=1'b0;
    defparam buf_dds0_i7_LC_13_16_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i7_LC_13_16_3.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i7_LC_13_16_3 (
            .in0(N__38950),
            .in1(N__49720),
            .in2(N__47680),
            .in3(N__44562),
            .lcout(buf_dds0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57914),
            .ce(),
            .sr(_gnd_net_));
    defparam i19179_3_lut_4_lut_LC_13_16_5.C_ON=1'b0;
    defparam i19179_3_lut_4_lut_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam i19179_3_lut_4_lut_LC_13_16_5.LUT_INIT=16'b0000000000000111;
    LogicCell40 i19179_3_lut_4_lut_LC_13_16_5 (
            .in0(N__36707),
            .in1(N__36433),
            .in2(N__41054),
            .in3(N__36344),
            .lcout(n11670),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_5_i16_3_lut_LC_13_16_6.C_ON=1'b0;
    defparam mux_135_Mux_5_i16_3_lut_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_5_i16_3_lut_LC_13_16_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_5_i16_3_lut_LC_13_16_6 (
            .in0(N__36291),
            .in1(N__36547),
            .in2(_gnd_net_),
            .in3(N__56298),
            .lcout(n16_adj_1496),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_12224_12225_set_LC_13_17_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12224_12225_set_LC_13_17_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i3_12224_12225_set_LC_13_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12224_12225_set_LC_13_17_0  (
            .in0(N__55400),
            .in1(N__55373),
            .in2(_gnd_net_),
            .in3(N__55349),
            .lcout(\comm_spi.n14642 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57035),
            .ce(),
            .sr(N__41930));
    defparam i19065_2_lut_LC_13_17_3.C_ON=1'b0;
    defparam i19065_2_lut_LC_13_17_3.SEQ_MODE=4'b0000;
    defparam i19065_2_lut_LC_13_17_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19065_2_lut_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(N__36275),
            .in2(_gnd_net_),
            .in3(N__56340),
            .lcout(n21037),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19118_2_lut_LC_13_17_5.C_ON=1'b0;
    defparam i19118_2_lut_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam i19118_2_lut_LC_13_17_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19118_2_lut_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(N__36709),
            .in2(_gnd_net_),
            .in3(N__36617),
            .lcout(n14687),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_237_LC_13_17_6.C_ON=1'b0;
    defparam i1_2_lut_adj_237_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_237_LC_13_17_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_237_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__36586),
            .in2(_gnd_net_),
            .in3(N__46581),
            .lcout(n10713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_13_18_3.C_ON=1'b0;
    defparam i9_4_lut_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_13_18_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_13_18_3 (
            .in0(N__39886),
            .in1(N__39709),
            .in2(N__39575),
            .in3(N__39511),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i5_LC_13_18_4.C_ON=1'b0;
    defparam buf_dds0_i5_LC_13_18_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i5_LC_13_18_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i5_LC_13_18_4 (
            .in0(N__49781),
            .in1(N__36543),
            .in2(N__45917),
            .in3(N__38966),
            .lcout(buf_dds0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57940),
            .ce(),
            .sr(_gnd_net_));
    defparam i18827_2_lut_LC_13_18_7.C_ON=1'b0;
    defparam i18827_2_lut_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam i18827_2_lut_LC_13_18_7.LUT_INIT=16'b0000000010101010;
    LogicCell40 i18827_2_lut_LC_13_18_7 (
            .in0(N__42041),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56363),
            .lcout(n21067),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_174_LC_13_19_0.C_ON=1'b0;
    defparam i11_4_lut_adj_174_LC_13_19_0.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_174_LC_13_19_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_174_LC_13_19_0 (
            .in0(N__39496),
            .in1(N__39610),
            .in2(N__39680),
            .in3(N__39541),
            .lcout(),
            .ltout(n27_adj_1551_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_13_19_1.C_ON=1'b0;
    defparam i15_4_lut_LC_13_19_1.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_13_19_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_LC_13_19_1 (
            .in0(N__36977),
            .in1(N__36506),
            .in2(N__36524),
            .in3(N__36521),
            .lcout(),
            .ltout(n19608_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_187_LC_13_19_2.C_ON=1'b0;
    defparam i7_4_lut_adj_187_LC_13_19_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_187_LC_13_19_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 i7_4_lut_adj_187_LC_13_19_2 (
            .in0(N__39808),
            .in1(N__36971),
            .in2(N__36515),
            .in3(N__36512),
            .lcout(n14731),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_175_LC_13_19_3.C_ON=1'b0;
    defparam i2_2_lut_adj_175_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_175_LC_13_19_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i2_2_lut_adj_175_LC_13_19_3 (
            .in0(N__39694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39856),
            .lcout(n10_adj_1594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_173_LC_13_19_4.C_ON=1'b0;
    defparam i10_4_lut_adj_173_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_173_LC_13_19_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_173_LC_13_19_4 (
            .in0(N__39871),
            .in1(N__39724),
            .in2(N__39629),
            .in3(N__39556),
            .lcout(n26_adj_1543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_172_LC_13_19_5.C_ON=1'b0;
    defparam i12_4_lut_adj_172_LC_13_19_5.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_172_LC_13_19_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_172_LC_13_19_5 (
            .in0(N__39526),
            .in1(N__39589),
            .in2(N__39842),
            .in3(N__39661),
            .lcout(n28_adj_1621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_177_LC_13_20_1.C_ON=1'b0;
    defparam i6_4_lut_adj_177_LC_13_20_1.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_177_LC_13_20_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_adj_177_LC_13_20_1 (
            .in0(N__39793),
            .in1(N__39823),
            .in2(N__39647),
            .in3(N__39775),
            .lcout(n14_adj_1592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22112_bdd_4_lut_LC_14_4_0.C_ON=1'b0;
    defparam n22112_bdd_4_lut_LC_14_4_0.SEQ_MODE=4'b0000;
    defparam n22112_bdd_4_lut_LC_14_4_0.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22112_bdd_4_lut_LC_14_4_0 (
            .in0(N__48362),
            .in1(N__36965),
            .in2(N__36926),
            .in3(N__36779),
            .lcout(),
            .ltout(n22115_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18242_3_lut_LC_14_4_1.C_ON=1'b0;
    defparam i18242_3_lut_LC_14_4_1.SEQ_MODE=4'b0000;
    defparam i18242_3_lut_LC_14_4_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 i18242_3_lut_LC_14_4_1 (
            .in0(_gnd_net_),
            .in1(N__49118),
            .in2(N__36887),
            .in3(N__36884),
            .lcout(n20856),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19509_LC_14_4_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19509_LC_14_4_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19509_LC_14_4_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19509_LC_14_4_3 (
            .in0(N__36865),
            .in1(N__48361),
            .in2(N__36824),
            .in3(N__56299),
            .lcout(n22112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19439_LC_14_4_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19439_LC_14_4_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19439_LC_14_4_4.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19439_LC_14_4_4 (
            .in0(N__48363),
            .in1(N__42629),
            .in2(N__36773),
            .in3(N__49119),
            .lcout(),
            .ltout(n22070_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22070_bdd_4_lut_LC_14_4_5.C_ON=1'b0;
    defparam n22070_bdd_4_lut_LC_14_4_5.SEQ_MODE=4'b0000;
    defparam n22070_bdd_4_lut_LC_14_4_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22070_bdd_4_lut_LC_14_4_5 (
            .in0(N__49120),
            .in1(N__36752),
            .in2(N__36737),
            .in3(N__39170),
            .lcout(),
            .ltout(n22073_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1544855_i1_3_lut_LC_14_4_6.C_ON=1'b0;
    defparam i1544855_i1_3_lut_LC_14_4_6.SEQ_MODE=4'b0000;
    defparam i1544855_i1_3_lut_LC_14_4_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1544855_i1_3_lut_LC_14_4_6 (
            .in0(_gnd_net_),
            .in1(N__36734),
            .in2(N__36728),
            .in3(N__48729),
            .lcout(),
            .ltout(n30_adj_1535_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i6_LC_14_4_7.C_ON=1'b0;
    defparam comm_buf_0__i6_LC_14_4_7.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i6_LC_14_4_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i6_LC_14_4_7 (
            .in0(N__40198),
            .in1(_gnd_net_),
            .in2(N__37283),
            .in3(N__54077),
            .lcout(comm_buf_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57812),
            .ce(N__42723),
            .sr(N__42851));
    defparam \ADC_VDC.genclk.i18784_4_lut_LC_14_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i18784_4_lut_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i18784_4_lut_LC_14_5_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i18784_4_lut_LC_14_5_0  (
            .in0(N__37276),
            .in1(N__37264),
            .in2(N__37253),
            .in3(N__37231),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n21211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i18825_4_lut_LC_14_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i18825_4_lut_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i18825_4_lut_LC_14_5_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i18825_4_lut_LC_14_5_1  (
            .in0(N__37085),
            .in1(N__37145),
            .in2(N__37220),
            .in3(N__37019),
            .lcout(\ADC_VDC.genclk.n21205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_adj_25_LC_14_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_25_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_25_LC_14_5_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_adj_25_LC_14_5_2  (
            .in0(N__37198),
            .in1(N__37186),
            .in2(N__37175),
            .in3(N__37156),
            .lcout(\ADC_VDC.genclk.n26_adj_1408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_adj_24_LC_14_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_24_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_24_LC_14_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_adj_24_LC_14_5_3  (
            .in0(N__37135),
            .in1(N__37123),
            .in2(N__37112),
            .in3(N__37096),
            .lcout(\ADC_VDC.genclk.n28_adj_1407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_adj_26_LC_14_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_26_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_26_LC_14_5_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_adj_26_LC_14_5_4  (
            .in0(N__37075),
            .in1(N__37060),
            .in2(N__37049),
            .in3(N__37030),
            .lcout(\ADC_VDC.genclk.n27_adj_1409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i0_LC_14_6_0.C_ON=1'b0;
    defparam comm_buf_3__i0_LC_14_6_0.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i0_LC_14_6_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_3__i0_LC_14_6_0 (
            .in0(N__37013),
            .in1(N__54082),
            .in2(_gnd_net_),
            .in3(N__50761),
            .lcout(comm_buf_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i4_LC_14_6_1.C_ON=1'b0;
    defparam comm_buf_3__i4_LC_14_6_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i4_LC_14_6_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i4_LC_14_6_1 (
            .in0(N__54080),
            .in1(N__40620),
            .in2(_gnd_net_),
            .in3(N__37001),
            .lcout(comm_buf_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i7_LC_14_6_2.C_ON=1'b0;
    defparam comm_buf_3__i7_LC_14_6_2.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i7_LC_14_6_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i7_LC_14_6_2 (
            .in0(N__51383),
            .in1(N__37403),
            .in2(_gnd_net_),
            .in3(N__54085),
            .lcout(comm_buf_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i6_LC_14_6_3.C_ON=1'b0;
    defparam comm_buf_3__i6_LC_14_6_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i6_LC_14_6_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i6_LC_14_6_3 (
            .in0(N__54081),
            .in1(N__40215),
            .in2(_gnd_net_),
            .in3(N__37385),
            .lcout(comm_buf_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i5_LC_14_6_4.C_ON=1'b0;
    defparam comm_buf_3__i5_LC_14_6_4.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i5_LC_14_6_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i5_LC_14_6_4 (
            .in0(N__51032),
            .in1(N__37370),
            .in2(_gnd_net_),
            .in3(N__54084),
            .lcout(comm_buf_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i3_LC_14_6_5.C_ON=1'b0;
    defparam comm_buf_3__i3_LC_14_6_5.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i3_LC_14_6_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i3_LC_14_6_5 (
            .in0(N__54079),
            .in1(N__40757),
            .in2(_gnd_net_),
            .in3(N__37355),
            .lcout(comm_buf_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i2_LC_14_6_6.C_ON=1'b0;
    defparam comm_buf_3__i2_LC_14_6_6.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i2_LC_14_6_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i2_LC_14_6_6 (
            .in0(N__47221),
            .in1(N__37340),
            .in2(_gnd_net_),
            .in3(N__54083),
            .lcout(comm_buf_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam comm_buf_3__i1_LC_14_6_7.C_ON=1'b0;
    defparam comm_buf_3__i1_LC_14_6_7.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i1_LC_14_6_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i1_LC_14_6_7 (
            .in0(N__54078),
            .in1(N__45362),
            .in2(_gnd_net_),
            .in3(N__37322),
            .lcout(comm_buf_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57820),
            .ce(N__37304),
            .sr(N__37292));
    defparam mux_143_Mux_0_i1_3_lut_LC_14_7_0.C_ON=1'b0;
    defparam mux_143_Mux_0_i1_3_lut_LC_14_7_0.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_0_i1_3_lut_LC_14_7_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_143_Mux_0_i1_3_lut_LC_14_7_0 (
            .in0(N__41500),
            .in1(N__41157),
            .in2(_gnd_net_),
            .in3(N__54373),
            .lcout(),
            .ltout(n1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i0_LC_14_7_1.C_ON=1'b0;
    defparam comm_tx_buf_i0_LC_14_7_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i0_LC_14_7_1.LUT_INIT=16'b1110111001010000;
    LogicCell40 comm_tx_buf_i0_LC_14_7_1 (
            .in0(N__50680),
            .in1(N__37553),
            .in2(N__37286),
            .in3(N__37526),
            .lcout(comm_tx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57824),
            .ce(N__46218),
            .sr(N__46115));
    defparam i18722_2_lut_LC_14_7_2.C_ON=1'b0;
    defparam i18722_2_lut_LC_14_7_2.SEQ_MODE=4'b0000;
    defparam i18722_2_lut_LC_14_7_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18722_2_lut_LC_14_7_2 (
            .in0(_gnd_net_),
            .in1(N__50702),
            .in2(_gnd_net_),
            .in3(N__54370),
            .lcout(n20970),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_0_i2_3_lut_LC_14_7_3.C_ON=1'b0;
    defparam mux_143_Mux_0_i2_3_lut_LC_14_7_3.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_0_i2_3_lut_LC_14_7_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_143_Mux_0_i2_3_lut_LC_14_7_3 (
            .in0(N__54372),
            .in1(_gnd_net_),
            .in2(N__37571),
            .in3(N__37562),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_0_i4_3_lut_LC_14_7_4.C_ON=1'b0;
    defparam mux_143_Mux_0_i4_3_lut_LC_14_7_4.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_0_i4_3_lut_LC_14_7_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_143_Mux_0_i4_3_lut_LC_14_7_4 (
            .in0(N__37547),
            .in1(N__37457),
            .in2(_gnd_net_),
            .in3(N__54371),
            .lcout(),
            .ltout(n4_adj_1507_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19366_LC_14_7_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19366_LC_14_7_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19366_LC_14_7_5.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_index_1__bdd_4_lut_19366_LC_14_7_5 (
            .in0(N__50679),
            .in1(N__37535),
            .in2(N__37529),
            .in3(N__50545),
            .lcout(n21980),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19011_2_lut_3_lut_LC_14_7_6.C_ON=1'b0;
    defparam i19011_2_lut_3_lut_LC_14_7_6.SEQ_MODE=4'b0000;
    defparam i19011_2_lut_3_lut_LC_14_7_6.LUT_INIT=16'b0010001000000000;
    LogicCell40 i19011_2_lut_3_lut_LC_14_7_6 (
            .in0(N__50544),
            .in1(N__50678),
            .in2(_gnd_net_),
            .in3(N__43059),
            .lcout(),
            .ltout(n21116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_LC_14_7_7.C_ON=1'b0;
    defparam i19_4_lut_LC_14_7_7.SEQ_MODE=4'b0000;
    defparam i19_4_lut_LC_14_7_7.LUT_INIT=16'b1000000010110011;
    LogicCell40 i19_4_lut_LC_14_7_7 (
            .in0(N__54369),
            .in1(N__54075),
            .in2(N__37520),
            .in3(N__37512),
            .lcout(n12_adj_1602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i0_LC_14_8_0.C_ON=1'b0;
    defparam comm_buf_4__i0_LC_14_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i0_LC_14_8_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i0_LC_14_8_0 (
            .in0(N__37472),
            .in1(N__54071),
            .in2(_gnd_net_),
            .in3(N__50777),
            .lcout(comm_buf_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i7_LC_14_8_1.C_ON=1'b0;
    defparam comm_buf_4__i7_LC_14_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i7_LC_14_8_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_4__i7_LC_14_8_1 (
            .in0(N__54070),
            .in1(_gnd_net_),
            .in2(N__51398),
            .in3(N__37451),
            .lcout(comm_buf_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i6_LC_14_8_2.C_ON=1'b0;
    defparam comm_buf_4__i6_LC_14_8_2.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i6_LC_14_8_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_4__i6_LC_14_8_2 (
            .in0(N__40233),
            .in1(N__54074),
            .in2(_gnd_net_),
            .in3(N__37433),
            .lcout(comm_buf_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i5_LC_14_8_3.C_ON=1'b0;
    defparam comm_buf_4__i5_LC_14_8_3.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i5_LC_14_8_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_4__i5_LC_14_8_3 (
            .in0(N__54069),
            .in1(_gnd_net_),
            .in2(N__51047),
            .in3(N__37421),
            .lcout(comm_buf_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i4_LC_14_8_4.C_ON=1'b0;
    defparam comm_buf_4__i4_LC_14_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i4_LC_14_8_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_4__i4_LC_14_8_4 (
            .in0(N__40638),
            .in1(N__54073),
            .in2(_gnd_net_),
            .in3(N__37739),
            .lcout(comm_buf_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i3_LC_14_8_5.C_ON=1'b0;
    defparam comm_buf_4__i3_LC_14_8_5.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i3_LC_14_8_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i3_LC_14_8_5 (
            .in0(N__54068),
            .in1(N__40792),
            .in2(_gnd_net_),
            .in3(N__37709),
            .lcout(comm_buf_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i2_LC_14_8_6.C_ON=1'b0;
    defparam comm_buf_4__i2_LC_14_8_6.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i2_LC_14_8_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_4__i2_LC_14_8_6 (
            .in0(N__47234),
            .in1(N__54072),
            .in2(_gnd_net_),
            .in3(N__37688),
            .lcout(comm_buf_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam comm_buf_4__i1_LC_14_8_7.C_ON=1'b0;
    defparam comm_buf_4__i1_LC_14_8_7.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i1_LC_14_8_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i1_LC_14_8_7 (
            .in0(N__54067),
            .in1(N__45363),
            .in2(_gnd_net_),
            .in3(N__37667),
            .lcout(comm_buf_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57833),
            .ce(N__37646),
            .sr(N__37634));
    defparam mux_143_Mux_3_i1_3_lut_LC_14_9_0.C_ON=1'b0;
    defparam mux_143_Mux_3_i1_3_lut_LC_14_9_0.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_3_i1_3_lut_LC_14_9_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_143_Mux_3_i1_3_lut_LC_14_9_0 (
            .in0(N__37969),
            .in1(N__54331),
            .in2(_gnd_net_),
            .in3(N__44259),
            .lcout(),
            .ltout(n1_adj_1589_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i3_LC_14_9_1.C_ON=1'b0;
    defparam comm_tx_buf_i3_LC_14_9_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i3_LC_14_9_1.LUT_INIT=16'b1100110010111000;
    LogicCell40 comm_tx_buf_i3_LC_14_9_1 (
            .in0(N__37808),
            .in1(N__37601),
            .in2(N__37622),
            .in3(N__50667),
            .lcout(comm_tx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57843),
            .ce(N__46212),
            .sr(N__46141));
    defparam i19059_2_lut_LC_14_9_2.C_ON=1'b0;
    defparam i19059_2_lut_LC_14_9_2.SEQ_MODE=4'b0000;
    defparam i19059_2_lut_LC_14_9_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19059_2_lut_LC_14_9_2 (
            .in0(_gnd_net_),
            .in1(N__54329),
            .in2(_gnd_net_),
            .in3(N__37619),
            .lcout(),
            .ltout(n21296_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_LC_14_9_3.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_LC_14_9_3.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_LC_14_9_3.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_1__bdd_4_lut_LC_14_9_3 (
            .in0(N__50533),
            .in1(N__37577),
            .in2(N__37604),
            .in3(N__50666),
            .lcout(n22154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_3_i4_3_lut_LC_14_9_4.C_ON=1'b0;
    defparam mux_143_Mux_3_i4_3_lut_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_3_i4_3_lut_LC_14_9_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_143_Mux_3_i4_3_lut_LC_14_9_4 (
            .in0(N__37595),
            .in1(N__54328),
            .in2(_gnd_net_),
            .in3(N__37589),
            .lcout(n4_adj_1591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_3_i2_3_lut_LC_14_9_5.C_ON=1'b0;
    defparam mux_143_Mux_3_i2_3_lut_LC_14_9_5.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_3_i2_3_lut_LC_14_9_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_143_Mux_3_i2_3_lut_LC_14_9_5 (
            .in0(N__54330),
            .in1(N__37832),
            .in2(_gnd_net_),
            .in3(N__37823),
            .lcout(n2_adj_1590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18879_3_lut_LC_14_9_6.C_ON=1'b0;
    defparam i18879_3_lut_LC_14_9_6.SEQ_MODE=4'b0000;
    defparam i18879_3_lut_LC_14_9_6.LUT_INIT=16'b0011000000000000;
    LogicCell40 i18879_3_lut_LC_14_9_6 (
            .in0(_gnd_net_),
            .in1(N__54327),
            .in2(N__43271),
            .in3(N__50532),
            .lcout(),
            .ltout(n21102_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i40_4_lut_LC_14_9_7.C_ON=1'b0;
    defparam i40_4_lut_LC_14_9_7.SEQ_MODE=4'b0000;
    defparam i40_4_lut_LC_14_9_7.LUT_INIT=16'b1110001011000000;
    LogicCell40 i40_4_lut_LC_14_9_7 (
            .in0(N__45193),
            .in1(N__54022),
            .in2(N__37802),
            .in3(N__37799),
            .lcout(n16_adj_1599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_6_i26_3_lut_LC_14_10_0.C_ON=1'b0;
    defparam mux_135_Mux_6_i26_3_lut_LC_14_10_0.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_6_i26_3_lut_LC_14_10_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_135_Mux_6_i26_3_lut_LC_14_10_0 (
            .in0(N__56007),
            .in1(N__37787),
            .in2(_gnd_net_),
            .in3(N__46522),
            .lcout(),
            .ltout(n26_adj_1505_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18316_4_lut_LC_14_10_1.C_ON=1'b0;
    defparam i18316_4_lut_LC_14_10_1.SEQ_MODE=4'b0000;
    defparam i18316_4_lut_LC_14_10_1.LUT_INIT=16'b1111101011011000;
    LogicCell40 i18316_4_lut_LC_14_10_1 (
            .in0(N__48153),
            .in1(N__37766),
            .in2(N__37751),
            .in3(N__56008),
            .lcout(),
            .ltout(n20930_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19424_LC_14_10_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19424_LC_14_10_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19424_LC_14_10_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19424_LC_14_10_2 (
            .in0(N__37991),
            .in1(N__48685),
            .in2(N__37748),
            .in3(N__48954),
            .lcout(),
            .ltout(n21962_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21962_bdd_4_lut_LC_14_10_3.C_ON=1'b0;
    defparam n21962_bdd_4_lut_LC_14_10_3.SEQ_MODE=4'b0000;
    defparam n21962_bdd_4_lut_LC_14_10_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n21962_bdd_4_lut_LC_14_10_3 (
            .in0(N__48686),
            .in1(N__38030),
            .in2(N__37745),
            .in3(N__38324),
            .lcout(),
            .ltout(n21965_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i6_LC_14_10_4.C_ON=1'b0;
    defparam comm_buf_1__i6_LC_14_10_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i6_LC_14_10_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_1__i6_LC_14_10_4 (
            .in0(N__54086),
            .in1(_gnd_net_),
            .in2(N__37742),
            .in3(N__40244),
            .lcout(comm_buf_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57853),
            .ce(N__47054),
            .sr(N__46969));
    defparam mux_135_Mux_6_i19_3_lut_LC_14_10_5.C_ON=1'b0;
    defparam mux_135_Mux_6_i19_3_lut_LC_14_10_5.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_6_i19_3_lut_LC_14_10_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_6_i19_3_lut_LC_14_10_5 (
            .in0(N__38108),
            .in1(N__38076),
            .in2(_gnd_net_),
            .in3(N__56006),
            .lcout(),
            .ltout(n19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18340_3_lut_LC_14_10_6.C_ON=1'b0;
    defparam i18340_3_lut_LC_14_10_6.SEQ_MODE=4'b0000;
    defparam i18340_3_lut_LC_14_10_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i18340_3_lut_LC_14_10_6 (
            .in0(_gnd_net_),
            .in1(N__38051),
            .in2(N__38033),
            .in3(N__48152),
            .lcout(n20954),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18315_3_lut_LC_14_10_7.C_ON=1'b0;
    defparam i18315_3_lut_LC_14_10_7.SEQ_MODE=4'b0000;
    defparam i18315_3_lut_LC_14_10_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 i18315_3_lut_LC_14_10_7 (
            .in0(N__48151),
            .in1(_gnd_net_),
            .in2(N__38021),
            .in3(N__46331),
            .lcout(n20929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i3_LC_14_11_0.C_ON=1'b0;
    defparam comm_buf_1__i3_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i3_LC_14_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i3_LC_14_11_0 (
            .in0(N__40797),
            .in1(N__54087),
            .in2(_gnd_net_),
            .in3(N__37886),
            .lcout(comm_buf_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57863),
            .ce(N__47069),
            .sr(N__47000));
    defparam i18270_3_lut_LC_14_11_1.C_ON=1'b0;
    defparam i18270_3_lut_LC_14_11_1.SEQ_MODE=4'b0000;
    defparam i18270_3_lut_LC_14_11_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18270_3_lut_LC_14_11_1 (
            .in0(N__48312),
            .in1(N__47708),
            .in2(_gnd_net_),
            .in3(N__37931),
            .lcout(),
            .ltout(n20884_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19557_LC_14_11_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19557_LC_14_11_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19557_LC_14_11_2.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19557_LC_14_11_2 (
            .in0(N__48597),
            .in1(N__49075),
            .in2(N__37907),
            .in3(N__37838),
            .lcout(),
            .ltout(n22124_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22124_bdd_4_lut_LC_14_11_3.C_ON=1'b0;
    defparam n22124_bdd_4_lut_LC_14_11_3.SEQ_MODE=4'b0000;
    defparam n22124_bdd_4_lut_LC_14_11_3.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22124_bdd_4_lut_LC_14_11_3 (
            .in0(N__37904),
            .in1(N__38300),
            .in2(N__37889),
            .in3(N__48598),
            .lcout(n22127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_3_i26_3_lut_LC_14_11_4.C_ON=1'b0;
    defparam mux_135_Mux_3_i26_3_lut_LC_14_11_4.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_3_i26_3_lut_LC_14_11_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_3_i26_3_lut_LC_14_11_4 (
            .in0(N__37876),
            .in1(N__56269),
            .in2(_gnd_net_),
            .in3(N__47731),
            .lcout(),
            .ltout(n26_adj_1514_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18271_4_lut_LC_14_11_5.C_ON=1'b0;
    defparam i18271_4_lut_LC_14_11_5.SEQ_MODE=4'b0000;
    defparam i18271_4_lut_LC_14_11_5.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18271_4_lut_LC_14_11_5 (
            .in0(N__56270),
            .in1(N__37862),
            .in2(N__37841),
            .in3(N__48310),
            .lcout(n20885),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18265_3_lut_LC_14_11_6.C_ON=1'b0;
    defparam i18265_3_lut_LC_14_11_6.SEQ_MODE=4'b0000;
    defparam i18265_3_lut_LC_14_11_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 i18265_3_lut_LC_14_11_6 (
            .in0(N__38237),
            .in1(N__38315),
            .in2(_gnd_net_),
            .in3(N__48311),
            .lcout(n20879),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_3_i19_3_lut_LC_14_11_7.C_ON=1'b0;
    defparam mux_135_Mux_3_i19_3_lut_LC_14_11_7.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_3_i19_3_lut_LC_14_11_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_135_Mux_3_i19_3_lut_LC_14_11_7 (
            .in0(N__56268),
            .in1(N__38286),
            .in2(_gnd_net_),
            .in3(N__38258),
            .lcout(n19_adj_1513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19533_LC_14_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19533_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19533_LC_14_12_0.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19533_LC_14_12_0 (
            .in0(N__48315),
            .in1(N__49050),
            .in2(N__52571),
            .in3(N__38198),
            .lcout(),
            .ltout(n22178_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22178_bdd_4_lut_LC_14_12_1.C_ON=1'b0;
    defparam n22178_bdd_4_lut_LC_14_12_1.SEQ_MODE=4'b0000;
    defparam n22178_bdd_4_lut_LC_14_12_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22178_bdd_4_lut_LC_14_12_1 (
            .in0(N__49051),
            .in1(N__49283),
            .in2(N__38231),
            .in3(N__46724),
            .lcout(),
            .ltout(n22181_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1547870_i1_3_lut_LC_14_12_2.C_ON=1'b0;
    defparam i1547870_i1_3_lut_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam i1547870_i1_3_lut_LC_14_12_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1547870_i1_3_lut_LC_14_12_2 (
            .in0(_gnd_net_),
            .in1(N__38618),
            .in2(N__38228),
            .in3(N__48701),
            .lcout(),
            .ltout(n30_adj_1511_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i4_LC_14_12_3.C_ON=1'b0;
    defparam comm_buf_1__i4_LC_14_12_3.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i4_LC_14_12_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i4_LC_14_12_3 (
            .in0(N__40650),
            .in1(_gnd_net_),
            .in2(N__38225),
            .in3(N__54088),
            .lcout(comm_buf_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57873),
            .ce(N__47071),
            .sr(N__46995));
    defparam mux_135_Mux_4_i26_3_lut_LC_14_12_5.C_ON=1'b0;
    defparam mux_135_Mux_4_i26_3_lut_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_4_i26_3_lut_LC_14_12_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_4_i26_3_lut_LC_14_12_5 (
            .in0(N__38222),
            .in1(N__56184),
            .in2(_gnd_net_),
            .in3(N__46740),
            .lcout(n26_adj_1510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19400_LC_14_12_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19400_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19400_LC_14_12_6.LUT_INIT=16'b1110110000101100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19400_LC_14_12_6 (
            .in0(N__38192),
            .in1(N__48314),
            .in2(N__49127),
            .in3(N__38186),
            .lcout(),
            .ltout(n22010_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22010_bdd_4_lut_LC_14_12_7.C_ON=1'b0;
    defparam n22010_bdd_4_lut_LC_14_12_7.SEQ_MODE=4'b0000;
    defparam n22010_bdd_4_lut_LC_14_12_7.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22010_bdd_4_lut_LC_14_12_7 (
            .in0(N__49049),
            .in1(N__38161),
            .in2(N__38126),
            .in3(N__38123),
            .lcout(n22013),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_228_LC_14_13_0.C_ON=1'b0;
    defparam i1_4_lut_adj_228_LC_14_13_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_228_LC_14_13_0.LUT_INIT=16'b1000100010001010;
    LogicCell40 i1_4_lut_adj_228_LC_14_13_0 (
            .in0(N__54764),
            .in1(N__49593),
            .in2(N__39215),
            .in3(N__46585),
            .lcout(n12441),
            .ltout(n12441_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i1_LC_14_13_1.C_ON=1'b0;
    defparam acadc_skipCount_i1_LC_14_13_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i1_LC_14_13_1.LUT_INIT=16'b0010111100100000;
    LogicCell40 acadc_skipCount_i1_LC_14_13_1 (
            .in0(N__45456),
            .in1(N__49630),
            .in2(N__38612),
            .in3(N__43395),
            .lcout(acadc_skipCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57886),
            .ce(),
            .sr(_gnd_net_));
    defparam i6464_3_lut_LC_14_13_3.C_ON=1'b0;
    defparam i6464_3_lut_LC_14_13_3.SEQ_MODE=4'b0000;
    defparam i6464_3_lut_LC_14_13_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6464_3_lut_LC_14_13_3 (
            .in0(N__45454),
            .in1(N__38593),
            .in2(_gnd_net_),
            .in3(N__41746),
            .lcout(n8_adj_1567),
            .ltout(n8_adj_1567_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i1_LC_14_13_4.C_ON=1'b0;
    defparam data_index_i1_LC_14_13_4.SEQ_MODE=4'b1000;
    defparam data_index_i1_LC_14_13_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 data_index_i1_LC_14_13_4 (
            .in0(N__54765),
            .in1(N__49595),
            .in2(N__38609),
            .in3(N__42200),
            .lcout(data_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57886),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i13_LC_14_13_5.C_ON=1'b0;
    defparam acadc_skipCount_i13_LC_14_13_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i13_LC_14_13_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i13_LC_14_13_5 (
            .in0(N__49594),
            .in1(N__49344),
            .in2(N__46410),
            .in3(N__38839),
            .lcout(acadc_skipCount_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57886),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i1_LC_14_13_6.C_ON=1'b0;
    defparam buf_dds1_i1_LC_14_13_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i1_LC_14_13_6.LUT_INIT=16'b1100101000000000;
    LogicCell40 buf_dds1_i1_LC_14_13_6 (
            .in0(N__38388),
            .in1(N__45457),
            .in2(N__38579),
            .in3(N__38480),
            .lcout(buf_dds1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57886),
            .ce(),
            .sr(_gnd_net_));
    defparam i15262_2_lut_3_lut_LC_14_13_7.C_ON=1'b0;
    defparam i15262_2_lut_3_lut_LC_14_13_7.SEQ_MODE=4'b0000;
    defparam i15262_2_lut_3_lut_LC_14_13_7.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15262_2_lut_3_lut_LC_14_13_7 (
            .in0(N__45455),
            .in1(N__54124),
            .in2(_gnd_net_),
            .in3(N__52434),
            .lcout(n14_adj_1550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i4_LC_14_14_0.C_ON=1'b0;
    defparam buf_control_i4_LC_14_14_0.SEQ_MODE=4'b1000;
    defparam buf_control_i4_LC_14_14_0.LUT_INIT=16'b0100111101000000;
    LogicCell40 buf_control_i4_LC_14_14_0 (
            .in0(N__49592),
            .in1(N__44173),
            .in2(N__44440),
            .in3(N__39016),
            .lcout(VDC_RNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57898),
            .ce(),
            .sr(_gnd_net_));
    defparam i18339_3_lut_LC_14_14_1.C_ON=1'b0;
    defparam i18339_3_lut_LC_14_14_1.SEQ_MODE=4'b0000;
    defparam i18339_3_lut_LC_14_14_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18339_3_lut_LC_14_14_1 (
            .in0(N__38359),
            .in1(N__38336),
            .in2(_gnd_net_),
            .in3(N__48313),
            .lcout(n20953),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_239_LC_14_14_2.C_ON=1'b0;
    defparam i15_4_lut_adj_239_LC_14_14_2.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_239_LC_14_14_2.LUT_INIT=16'b1100010011110111;
    LogicCell40 i15_4_lut_adj_239_LC_14_14_2 (
            .in0(N__41748),
            .in1(N__54763),
            .in2(N__49700),
            .in3(N__39157),
            .lcout(n12312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i6_LC_14_14_3.C_ON=1'b0;
    defparam buf_control_i6_LC_14_14_3.SEQ_MODE=4'b1000;
    defparam buf_control_i6_LC_14_14_3.LUT_INIT=16'b0011000010111000;
    LogicCell40 buf_control_i6_LC_14_14_3 (
            .in0(N__43154),
            .in1(N__44434),
            .in2(N__45012),
            .in3(N__49590),
            .lcout(buf_control_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57898),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_4_i23_3_lut_LC_14_14_4.C_ON=1'b0;
    defparam mux_134_Mux_4_i23_3_lut_LC_14_14_4.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_4_i23_3_lut_LC_14_14_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_134_Mux_4_i23_3_lut_LC_14_14_4 (
            .in0(N__39015),
            .in1(N__56183),
            .in2(_gnd_net_),
            .in3(N__38999),
            .lcout(n23_adj_1538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i11_LC_14_14_6.C_ON=1'b0;
    defparam buf_dds0_i11_LC_14_14_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i11_LC_14_14_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i11_LC_14_14_6 (
            .in0(N__49591),
            .in1(N__40449),
            .in2(N__44301),
            .in3(N__38968),
            .lcout(buf_dds0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57898),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_67_i14_2_lut_LC_14_14_7.C_ON=1'b0;
    defparam equal_67_i14_2_lut_LC_14_14_7.SEQ_MODE=4'b0000;
    defparam equal_67_i14_2_lut_LC_14_14_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_67_i14_2_lut_LC_14_14_7 (
            .in0(_gnd_net_),
            .in1(N__38861),
            .in2(_gnd_net_),
            .in3(N__38835),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_170_LC_14_15_0.C_ON=1'b0;
    defparam i2_4_lut_adj_170_LC_14_15_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_170_LC_14_15_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_170_LC_14_15_0 (
            .in0(N__38813),
            .in1(N__49282),
            .in2(N__38795),
            .in3(N__43396),
            .lcout(n18_adj_1611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i4_LC_14_15_1.C_ON=1'b0;
    defparam data_index_i4_LC_14_15_1.SEQ_MODE=4'b1000;
    defparam data_index_i4_LC_14_15_1.LUT_INIT=16'b0010111000100010;
    LogicCell40 data_index_i4_LC_14_15_1 (
            .in0(N__38741),
            .in1(N__54871),
            .in2(N__49772),
            .in3(N__38725),
            .lcout(data_index_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57915),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_4_i15_4_lut_LC_14_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_4_i15_4_lut_LC_14_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_4_i15_4_lut_LC_14_15_2.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_state_3__I_0_365_Mux_4_i15_4_lut_LC_14_15_2 (
            .in0(N__54870),
            .in1(N__38740),
            .in2(N__38726),
            .in3(N__49682),
            .lcout(data_index_9_N_216_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_2_i15_4_lut_LC_14_15_3.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_2_i15_4_lut_LC_14_15_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_2_i15_4_lut_LC_14_15_3.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_365_Mux_2_i15_4_lut_LC_14_15_3 (
            .in0(N__54887),
            .in1(N__39442),
            .in2(N__49771),
            .in3(N__39431),
            .lcout(data_index_9_N_216_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i10_LC_14_15_4.C_ON=1'b0;
    defparam req_data_cnt_i10_LC_14_15_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i10_LC_14_15_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i10_LC_14_15_4 (
            .in0(N__39317),
            .in1(N__47413),
            .in2(_gnd_net_),
            .in3(N__42013),
            .lcout(req_data_cnt_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57915),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i15_LC_14_15_5.C_ON=1'b0;
    defparam acadc_skipCount_i15_LC_14_15_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i15_LC_14_15_5.LUT_INIT=16'b0111001001010000;
    LogicCell40 acadc_skipCount_i15_LC_14_15_5 (
            .in0(N__49356),
            .in1(N__49638),
            .in2(N__47795),
            .in3(N__46048),
            .lcout(acadc_skipCount_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57915),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i11_LC_14_15_6.C_ON=1'b0;
    defparam req_data_cnt_i11_LC_14_15_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i11_LC_14_15_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i11_LC_14_15_6 (
            .in0(N__39284),
            .in1(N__47414),
            .in2(_gnd_net_),
            .in3(N__44529),
            .lcout(req_data_cnt_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57915),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_14_15_7.C_ON=1'b0;
    defparam i6_4_lut_LC_14_15_7.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_14_15_7.LUT_INIT=16'b0111101111011110;
    LogicCell40 i6_4_lut_LC_14_15_7 (
            .in0(N__39257),
            .in1(N__39239),
            .in2(N__49181),
            .in3(N__46278),
            .lcout(n22_adj_1620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15172_2_lut_LC_14_16_0.C_ON=1'b0;
    defparam i15172_2_lut_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam i15172_2_lut_LC_14_16_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i15172_2_lut_LC_14_16_0 (
            .in0(N__42316),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42326),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_193_i9_2_lut_3_lut_LC_14_16_2.C_ON=1'b0;
    defparam equal_193_i9_2_lut_3_lut_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam equal_193_i9_2_lut_3_lut_LC_14_16_2.LUT_INIT=16'b1111111110111011;
    LogicCell40 equal_193_i9_2_lut_3_lut_LC_14_16_2 (
            .in0(N__48359),
            .in1(N__56296),
            .in2(_gnd_net_),
            .in3(N__49099),
            .lcout(n9_adj_1415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i14_LC_14_16_3.C_ON=1'b0;
    defparam req_data_cnt_i14_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i14_LC_14_16_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 req_data_cnt_i14_LC_14_16_3 (
            .in0(N__41765),
            .in1(_gnd_net_),
            .in2(N__39200),
            .in3(N__47412),
            .lcout(req_data_cnt_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57927),
            .ce(),
            .sr(_gnd_net_));
    defparam i18828_2_lut_LC_14_16_4.C_ON=1'b0;
    defparam i18828_2_lut_LC_14_16_4.SEQ_MODE=4'b0000;
    defparam i18828_2_lut_LC_14_16_4.LUT_INIT=16'b0011001100000000;
    LogicCell40 i18828_2_lut_LC_14_16_4 (
            .in0(_gnd_net_),
            .in1(N__56297),
            .in2(_gnd_net_),
            .in3(N__41764),
            .lcout(n21048),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i12_LC_14_16_5.C_ON=1'b0;
    defparam req_data_cnt_i12_LC_14_16_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i12_LC_14_16_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i12_LC_14_16_5 (
            .in0(N__44078),
            .in1(N__47411),
            .in2(_gnd_net_),
            .in3(N__42039),
            .lcout(req_data_cnt_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57927),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i1_LC_14_16_6.C_ON=1'b0;
    defparam buf_control_i1_LC_14_16_6.SEQ_MODE=4'b1000;
    defparam buf_control_i1_LC_14_16_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 buf_control_i1_LC_14_16_6 (
            .in0(N__45566),
            .in1(N__44439),
            .in2(N__44643),
            .in3(N__49776),
            .lcout(DDS_RNG_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57927),
            .ce(),
            .sr(_gnd_net_));
    defparam i17_3_lut_3_lut_LC_14_16_7.C_ON=1'b0;
    defparam i17_3_lut_3_lut_LC_14_16_7.SEQ_MODE=4'b0000;
    defparam i17_3_lut_3_lut_LC_14_16_7.LUT_INIT=16'b0001000110001000;
    LogicCell40 i17_3_lut_3_lut_LC_14_16_7 (
            .in0(N__54169),
            .in1(N__52407),
            .in2(_gnd_net_),
            .in3(N__53581),
            .lcout(n10_adj_1613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i0_LC_14_17_0.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i0_LC_14_17_0.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i0_LC_14_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i0_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(N__42353),
            .in2(_gnd_net_),
            .in3(N__39473),
            .lcout(dds0_mclkcnt_0),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(n19498),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i1_LC_14_17_1.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i1_LC_14_17_1.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i1_LC_14_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i1_LC_14_17_1 (
            .in0(_gnd_net_),
            .in1(N__42391),
            .in2(_gnd_net_),
            .in3(N__39470),
            .lcout(dds0_mclkcnt_1),
            .ltout(),
            .carryin(n19498),
            .carryout(n19499),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i2_LC_14_17_2.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i2_LC_14_17_2.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i2_LC_14_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i2_LC_14_17_2 (
            .in0(_gnd_net_),
            .in1(N__42365),
            .in2(_gnd_net_),
            .in3(N__39467),
            .lcout(dds0_mclkcnt_2),
            .ltout(),
            .carryin(n19499),
            .carryout(n19500),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i3_LC_14_17_3.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i3_LC_14_17_3.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i3_LC_14_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i3_LC_14_17_3 (
            .in0(_gnd_net_),
            .in1(N__42416),
            .in2(_gnd_net_),
            .in3(N__39464),
            .lcout(dds0_mclkcnt_3),
            .ltout(),
            .carryin(n19500),
            .carryout(n19501),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i4_LC_14_17_4.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i4_LC_14_17_4.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i4_LC_14_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i4_LC_14_17_4 (
            .in0(_gnd_net_),
            .in1(N__42377),
            .in2(_gnd_net_),
            .in3(N__39461),
            .lcout(dds0_mclkcnt_4),
            .ltout(),
            .carryin(n19501),
            .carryout(n19502),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i5_LC_14_17_5.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i5_LC_14_17_5.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i5_LC_14_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i5_LC_14_17_5 (
            .in0(_gnd_net_),
            .in1(N__42404),
            .in2(_gnd_net_),
            .in3(N__39458),
            .lcout(dds0_mclkcnt_5),
            .ltout(),
            .carryin(n19502),
            .carryout(n19503),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i6_LC_14_17_6.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3783__i6_LC_14_17_6.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i6_LC_14_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i6_LC_14_17_6 (
            .in0(_gnd_net_),
            .in1(N__39455),
            .in2(_gnd_net_),
            .in3(N__39596),
            .lcout(dds0_mclkcnt_6),
            .ltout(),
            .carryin(n19503),
            .carryout(n19504),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3783__i7_LC_14_17_7.C_ON=1'b0;
    defparam dds0_mclkcnt_i7_3783__i7_LC_14_17_7.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3783__i7_LC_14_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3783__i7_LC_14_17_7 (
            .in0(_gnd_net_),
            .in1(N__42338),
            .in2(_gnd_net_),
            .in3(N__39593),
            .lcout(dds0_mclkcnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclkcnt_i7_3783__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam secclk_cnt_3776_3777__i1_LC_14_18_0.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i1_LC_14_18_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i1_LC_14_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i1_LC_14_18_0 (
            .in0(_gnd_net_),
            .in1(N__39590),
            .in2(_gnd_net_),
            .in3(N__39578),
            .lcout(secclk_cnt_0),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(n19509),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i2_LC_14_18_1.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i2_LC_14_18_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i2_LC_14_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i2_LC_14_18_1 (
            .in0(_gnd_net_),
            .in1(N__39574),
            .in2(_gnd_net_),
            .in3(N__39560),
            .lcout(secclk_cnt_1),
            .ltout(),
            .carryin(n19509),
            .carryout(n19510),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i3_LC_14_18_2.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i3_LC_14_18_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i3_LC_14_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i3_LC_14_18_2 (
            .in0(_gnd_net_),
            .in1(N__39557),
            .in2(_gnd_net_),
            .in3(N__39545),
            .lcout(secclk_cnt_2),
            .ltout(),
            .carryin(n19510),
            .carryout(n19511),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i4_LC_14_18_3.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i4_LC_14_18_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i4_LC_14_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i4_LC_14_18_3 (
            .in0(_gnd_net_),
            .in1(N__39542),
            .in2(_gnd_net_),
            .in3(N__39530),
            .lcout(secclk_cnt_3),
            .ltout(),
            .carryin(n19511),
            .carryout(n19512),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i5_LC_14_18_4.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i5_LC_14_18_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i5_LC_14_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i5_LC_14_18_4 (
            .in0(_gnd_net_),
            .in1(N__39527),
            .in2(_gnd_net_),
            .in3(N__39515),
            .lcout(secclk_cnt_4),
            .ltout(),
            .carryin(n19512),
            .carryout(n19513),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i6_LC_14_18_5.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i6_LC_14_18_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i6_LC_14_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i6_LC_14_18_5 (
            .in0(_gnd_net_),
            .in1(N__39512),
            .in2(_gnd_net_),
            .in3(N__39500),
            .lcout(secclk_cnt_5),
            .ltout(),
            .carryin(n19513),
            .carryout(n19514),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i7_LC_14_18_6.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i7_LC_14_18_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i7_LC_14_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i7_LC_14_18_6 (
            .in0(_gnd_net_),
            .in1(N__39497),
            .in2(_gnd_net_),
            .in3(N__39485),
            .lcout(secclk_cnt_6),
            .ltout(),
            .carryin(n19514),
            .carryout(n19515),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i8_LC_14_18_7.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i8_LC_14_18_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i8_LC_14_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i8_LC_14_18_7 (
            .in0(_gnd_net_),
            .in1(N__39725),
            .in2(_gnd_net_),
            .in3(N__39713),
            .lcout(secclk_cnt_7),
            .ltout(),
            .carryin(n19515),
            .carryout(n19516),
            .clk(N__45084),
            .ce(),
            .sr(N__39763));
    defparam secclk_cnt_3776_3777__i9_LC_14_19_0.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i9_LC_14_19_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i9_LC_14_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i9_LC_14_19_0 (
            .in0(_gnd_net_),
            .in1(N__39710),
            .in2(_gnd_net_),
            .in3(N__39698),
            .lcout(secclk_cnt_8),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(n19517),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i10_LC_14_19_1.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i10_LC_14_19_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i10_LC_14_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i10_LC_14_19_1 (
            .in0(_gnd_net_),
            .in1(N__39695),
            .in2(_gnd_net_),
            .in3(N__39683),
            .lcout(secclk_cnt_9),
            .ltout(),
            .carryin(n19517),
            .carryout(n19518),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i11_LC_14_19_2.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i11_LC_14_19_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i11_LC_14_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i11_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(N__39679),
            .in2(_gnd_net_),
            .in3(N__39665),
            .lcout(secclk_cnt_10),
            .ltout(),
            .carryin(n19518),
            .carryout(n19519),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i12_LC_14_19_3.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i12_LC_14_19_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i12_LC_14_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i12_LC_14_19_3 (
            .in0(_gnd_net_),
            .in1(N__39662),
            .in2(_gnd_net_),
            .in3(N__39650),
            .lcout(secclk_cnt_11),
            .ltout(),
            .carryin(n19519),
            .carryout(n19520),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i13_LC_14_19_4.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i13_LC_14_19_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i13_LC_14_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i13_LC_14_19_4 (
            .in0(_gnd_net_),
            .in1(N__39646),
            .in2(_gnd_net_),
            .in3(N__39632),
            .lcout(secclk_cnt_12),
            .ltout(),
            .carryin(n19520),
            .carryout(n19521),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i14_LC_14_19_5.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i14_LC_14_19_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i14_LC_14_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i14_LC_14_19_5 (
            .in0(_gnd_net_),
            .in1(N__39628),
            .in2(_gnd_net_),
            .in3(N__39614),
            .lcout(secclk_cnt_13),
            .ltout(),
            .carryin(n19521),
            .carryout(n19522),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i15_LC_14_19_6.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i15_LC_14_19_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i15_LC_14_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i15_LC_14_19_6 (
            .in0(_gnd_net_),
            .in1(N__39611),
            .in2(_gnd_net_),
            .in3(N__39599),
            .lcout(secclk_cnt_14),
            .ltout(),
            .carryin(n19522),
            .carryout(n19523),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i16_LC_14_19_7.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i16_LC_14_19_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i16_LC_14_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i16_LC_14_19_7 (
            .in0(_gnd_net_),
            .in1(N__39887),
            .in2(_gnd_net_),
            .in3(N__39875),
            .lcout(secclk_cnt_15),
            .ltout(),
            .carryin(n19523),
            .carryout(n19524),
            .clk(N__45086),
            .ce(),
            .sr(N__39756));
    defparam secclk_cnt_3776_3777__i17_LC_14_20_0.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i17_LC_14_20_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i17_LC_14_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i17_LC_14_20_0 (
            .in0(_gnd_net_),
            .in1(N__39872),
            .in2(_gnd_net_),
            .in3(N__39860),
            .lcout(secclk_cnt_16),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(n19525),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam secclk_cnt_3776_3777__i18_LC_14_20_1.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i18_LC_14_20_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i18_LC_14_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i18_LC_14_20_1 (
            .in0(_gnd_net_),
            .in1(N__39857),
            .in2(_gnd_net_),
            .in3(N__39845),
            .lcout(secclk_cnt_17),
            .ltout(),
            .carryin(n19525),
            .carryout(n19526),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam secclk_cnt_3776_3777__i19_LC_14_20_2.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i19_LC_14_20_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i19_LC_14_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i19_LC_14_20_2 (
            .in0(_gnd_net_),
            .in1(N__39841),
            .in2(_gnd_net_),
            .in3(N__39827),
            .lcout(secclk_cnt_18),
            .ltout(),
            .carryin(n19526),
            .carryout(n19527),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam secclk_cnt_3776_3777__i20_LC_14_20_3.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i20_LC_14_20_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i20_LC_14_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i20_LC_14_20_3 (
            .in0(_gnd_net_),
            .in1(N__39824),
            .in2(_gnd_net_),
            .in3(N__39812),
            .lcout(secclk_cnt_19),
            .ltout(),
            .carryin(n19527),
            .carryout(n19528),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam secclk_cnt_3776_3777__i21_LC_14_20_4.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i21_LC_14_20_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i21_LC_14_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i21_LC_14_20_4 (
            .in0(_gnd_net_),
            .in1(N__39809),
            .in2(_gnd_net_),
            .in3(N__39797),
            .lcout(secclk_cnt_20),
            .ltout(),
            .carryin(n19528),
            .carryout(n19529),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam secclk_cnt_3776_3777__i22_LC_14_20_5.C_ON=1'b1;
    defparam secclk_cnt_3776_3777__i22_LC_14_20_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i22_LC_14_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i22_LC_14_20_5 (
            .in0(_gnd_net_),
            .in1(N__39794),
            .in2(_gnd_net_),
            .in3(N__39782),
            .lcout(secclk_cnt_21),
            .ltout(),
            .carryin(n19529),
            .carryout(n19530),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam secclk_cnt_3776_3777__i23_LC_14_20_6.C_ON=1'b0;
    defparam secclk_cnt_3776_3777__i23_LC_14_20_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3776_3777__i23_LC_14_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3776_3777__i23_LC_14_20_6 (
            .in0(_gnd_net_),
            .in1(N__39776),
            .in2(_gnd_net_),
            .in3(N__39779),
            .lcout(secclk_cnt_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45090),
            .ce(),
            .sr(N__39764));
    defparam \comm_spi.data_rx_i3_LC_15_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i3_LC_15_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i3_LC_15_4_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i3_LC_15_4_0  (
            .in0(N__42605),
            .in1(N__47181),
            .in2(_gnd_net_),
            .in3(N__40523),
            .lcout(comm_rx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \comm_spi.data_rx_i4_LC_15_4_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i4_LC_15_4_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i4_LC_15_4_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i4_LC_15_4_1  (
            .in0(N__40520),
            .in1(N__40736),
            .in2(_gnd_net_),
            .in3(N__42606),
            .lcout(comm_rx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \comm_spi.data_rx_i5_LC_15_4_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i5_LC_15_4_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i5_LC_15_4_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i5_LC_15_4_2  (
            .in0(N__42607),
            .in1(N__40599),
            .in2(_gnd_net_),
            .in3(N__40524),
            .lcout(comm_rx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \comm_spi.data_rx_i6_LC_15_4_3 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i6_LC_15_4_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i6_LC_15_4_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i6_LC_15_4_3  (
            .in0(N__40521),
            .in1(N__50994),
            .in2(_gnd_net_),
            .in3(N__42608),
            .lcout(comm_rx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \comm_spi.data_rx_i7_LC_15_4_4 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i7_LC_15_4_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i7_LC_15_4_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i7_LC_15_4_4  (
            .in0(N__42609),
            .in1(N__40197),
            .in2(_gnd_net_),
            .in3(N__40525),
            .lcout(comm_rx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \comm_spi.data_rx_i2_LC_15_4_5 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i2_LC_15_4_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i2_LC_15_4_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i2_LC_15_4_5  (
            .in0(N__40519),
            .in1(N__45321),
            .in2(_gnd_net_),
            .in3(N__42604),
            .lcout(comm_rx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \comm_spi.data_rx_i1_LC_15_4_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i1_LC_15_4_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i1_LC_15_4_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \comm_spi.data_rx_i1_LC_15_4_6  (
            .in0(N__42603),
            .in1(N__40522),
            .in2(_gnd_net_),
            .in3(N__50775),
            .lcout(comm_rx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57050),
            .ce(),
            .sr(N__56858));
    defparam \ADC_VDC.genclk.t_clk_24_LC_15_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t_clk_24_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t_clk_24_LC_15_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ADC_VDC.genclk.t_clk_24_LC_15_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40175),
            .lcout(VDC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t_clk_24C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i2_3_lut_LC_15_5_3 .C_ON=1'b0;
    defparam \comm_spi.i2_3_lut_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i2_3_lut_LC_15_5_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \comm_spi.i2_3_lut_LC_15_5_3  (
            .in0(N__42535),
            .in1(N__42557),
            .in2(_gnd_net_),
            .in3(N__42573),
            .lcout(\comm_spi.n16869 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12402_3_lut_LC_15_5_4.C_ON=1'b0;
    defparam i12402_3_lut_LC_15_5_4.SEQ_MODE=4'b0000;
    defparam i12402_3_lut_LC_15_5_4.LUT_INIT=16'b1100110001000100;
    LogicCell40 i12402_3_lut_LC_15_5_4 (
            .in0(N__40570),
            .in1(N__46219),
            .in2(_gnd_net_),
            .in3(N__54528),
            .lcout(n14815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18892_3_lut_LC_15_5_5.C_ON=1'b0;
    defparam i18892_3_lut_LC_15_5_5.SEQ_MODE=4'b0000;
    defparam i18892_3_lut_LC_15_5_5.LUT_INIT=16'b1010101010001000;
    LogicCell40 i18892_3_lut_LC_15_5_5 (
            .in0(N__54055),
            .in1(N__41102),
            .in2(_gnd_net_),
            .in3(N__40571),
            .lcout(),
            .ltout(n21506_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18269_4_lut_LC_15_5_6.C_ON=1'b0;
    defparam i18269_4_lut_LC_15_5_6.SEQ_MODE=4'b0000;
    defparam i18269_4_lut_LC_15_5_6.LUT_INIT=16'b1111110010101010;
    LogicCell40 i18269_4_lut_LC_15_5_6 (
            .in0(N__43217),
            .in1(N__45644),
            .in2(N__40424),
            .in3(N__52326),
            .lcout(n20883),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12353_2_lut_LC_15_5_7.C_ON=1'b0;
    defparam i12353_2_lut_LC_15_5_7.SEQ_MODE=4'b0000;
    defparam i12353_2_lut_LC_15_5_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12353_2_lut_LC_15_5_7 (
            .in0(N__54529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42689),
            .lcout(n14766),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22028_bdd_4_lut_LC_15_6_0.C_ON=1'b0;
    defparam n22028_bdd_4_lut_LC_15_6_0.SEQ_MODE=4'b0000;
    defparam n22028_bdd_4_lut_LC_15_6_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22028_bdd_4_lut_LC_15_6_0 (
            .in0(N__40421),
            .in1(N__40388),
            .in2(N__40406),
            .in3(N__49077),
            .lcout(n22031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19429_LC_15_6_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19429_LC_15_6_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19429_LC_15_6_2.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19429_LC_15_6_2 (
            .in0(N__48316),
            .in1(N__45233),
            .in2(N__40925),
            .in3(N__49076),
            .lcout(n22028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19459_LC_15_6_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19459_LC_15_6_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19459_LC_15_6_3.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19459_LC_15_6_3 (
            .in0(N__56368),
            .in1(N__41323),
            .in2(N__40381),
            .in3(N__48317),
            .lcout(),
            .ltout(n22088_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22088_bdd_4_lut_LC_15_6_4.C_ON=1'b0;
    defparam n22088_bdd_4_lut_LC_15_6_4.SEQ_MODE=4'b0000;
    defparam n22088_bdd_4_lut_LC_15_6_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22088_bdd_4_lut_LC_15_6_4 (
            .in0(N__48318),
            .in1(N__40340),
            .in2(N__40307),
            .in3(N__40304),
            .lcout(),
            .ltout(n22091_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18230_3_lut_LC_15_6_5.C_ON=1'b0;
    defparam i18230_3_lut_LC_15_6_5.SEQ_MODE=4'b0000;
    defparam i18230_3_lut_LC_15_6_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 i18230_3_lut_LC_15_6_5 (
            .in0(N__49078),
            .in1(_gnd_net_),
            .in2(N__40274),
            .in3(N__40271),
            .lcout(),
            .ltout(n20844_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1543649_i1_3_lut_LC_15_6_6.C_ON=1'b0;
    defparam i1543649_i1_3_lut_LC_15_6_6.SEQ_MODE=4'b0000;
    defparam i1543649_i1_3_lut_LC_15_6_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i1543649_i1_3_lut_LC_15_6_6 (
            .in0(_gnd_net_),
            .in1(N__40256),
            .in2(N__40250),
            .in3(N__48742),
            .lcout(),
            .ltout(n30_adj_1539_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i4_LC_15_6_7.C_ON=1'b0;
    defparam comm_buf_0__i4_LC_15_6_7.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i4_LC_15_6_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i4_LC_15_6_7 (
            .in0(N__40619),
            .in1(_gnd_net_),
            .in2(N__40574),
            .in3(N__54036),
            .lcout(comm_buf_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57825),
            .ce(N__42717),
            .sr(N__42831));
    defparam i1_2_lut_3_lut_4_lut_LC_15_7_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_15_7_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_15_7_0.LUT_INIT=16'b0000000000010000;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_15_7_0 (
            .in0(N__51828),
            .in1(N__50669),
            .in2(N__51669),
            .in3(N__40562),
            .lcout(n20596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_68_LC_15_7_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_68_LC_15_7_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_68_LC_15_7_1.LUT_INIT=16'b0000000100000000;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_68_LC_15_7_1 (
            .in0(N__40563),
            .in1(N__53549),
            .in2(N__51843),
            .in3(N__51642),
            .lcout(n20621),
            .ltout(n20621_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_248_LC_15_7_2.C_ON=1'b0;
    defparam i1_2_lut_adj_248_LC_15_7_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_248_LC_15_7_2.LUT_INIT=16'b0000000011110000;
    LogicCell40 i1_2_lut_adj_248_LC_15_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40535),
            .in3(N__50538),
            .lcout(),
            .ltout(n25_adj_1619_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_231_LC_15_7_3.C_ON=1'b0;
    defparam i1_4_lut_adj_231_LC_15_7_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_231_LC_15_7_3.LUT_INIT=16'b0001000011111111;
    LogicCell40 i1_4_lut_adj_231_LC_15_7_3 (
            .in0(N__50670),
            .in1(N__54352),
            .in2(N__40532),
            .in3(N__54030),
            .lcout(n4_adj_1616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_valid_85_LC_15_7_4 .C_ON=1'b0;
    defparam \comm_spi.data_valid_85_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_valid_85_LC_15_7_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.data_valid_85_LC_15_7_4  (
            .in0(N__40529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42617),
            .lcout(comm_data_vld),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.data_valid_85C_net ),
            .ce(),
            .sr(N__56854));
    defparam i22_4_lut_4_lut_LC_15_7_5.C_ON=1'b0;
    defparam i22_4_lut_4_lut_LC_15_7_5.SEQ_MODE=4'b0000;
    defparam i22_4_lut_4_lut_LC_15_7_5.LUT_INIT=16'b0010011000100010;
    LogicCell40 i22_4_lut_4_lut_LC_15_7_5 (
            .in0(N__53519),
            .in1(N__54031),
            .in2(N__51844),
            .in3(N__51646),
            .lcout(n7_adj_1609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_LC_15_7_7.C_ON=1'b0;
    defparam i2_4_lut_4_lut_LC_15_7_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_LC_15_7_7.LUT_INIT=16'b0111011111110011;
    LogicCell40 i2_4_lut_4_lut_LC_15_7_7 (
            .in0(N__53520),
            .in1(N__54032),
            .in2(N__51845),
            .in3(N__51647),
            .lcout(n20717),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22082_bdd_4_lut_LC_15_8_0.C_ON=1'b0;
    defparam n22082_bdd_4_lut_LC_15_8_0.SEQ_MODE=4'b0000;
    defparam n22082_bdd_4_lut_LC_15_8_0.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22082_bdd_4_lut_LC_15_8_0 (
            .in0(N__48293),
            .in1(N__40484),
            .in2(N__40456),
            .in3(N__40871),
            .lcout(n22085),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19449_LC_15_8_1.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19449_LC_15_8_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19449_LC_15_8_1.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19449_LC_15_8_1 (
            .in0(N__56185),
            .in1(N__41077),
            .in2(N__40909),
            .in3(N__48292),
            .lcout(n22082),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_3_i26_3_lut_LC_15_8_2.C_ON=1'b0;
    defparam mux_134_Mux_3_i26_3_lut_LC_15_8_2.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_3_i26_3_lut_LC_15_8_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_134_Mux_3_i26_3_lut_LC_15_8_2 (
            .in0(N__40865),
            .in1(N__56186),
            .in2(_gnd_net_),
            .in3(N__41786),
            .lcout(),
            .ltout(n26_adj_1541_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18223_4_lut_LC_15_8_3.C_ON=1'b0;
    defparam i18223_4_lut_LC_15_8_3.SEQ_MODE=4'b0000;
    defparam i18223_4_lut_LC_15_8_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18223_4_lut_LC_15_8_3 (
            .in0(N__56187),
            .in1(N__40844),
            .in2(N__40829),
            .in3(N__48294),
            .lcout(),
            .ltout(n20837_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19464_LC_15_8_4.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19464_LC_15_8_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19464_LC_15_8_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19464_LC_15_8_4 (
            .in0(N__44501),
            .in1(N__48736),
            .in2(N__40826),
            .in3(N__49053),
            .lcout(),
            .ltout(n22094_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22094_bdd_4_lut_LC_15_8_5.C_ON=1'b0;
    defparam n22094_bdd_4_lut_LC_15_8_5.SEQ_MODE=4'b0000;
    defparam n22094_bdd_4_lut_LC_15_8_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22094_bdd_4_lut_LC_15_8_5 (
            .in0(N__48737),
            .in1(N__40823),
            .in2(N__40817),
            .in3(N__40814),
            .lcout(),
            .ltout(n22097_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i3_LC_15_8_6.C_ON=1'b0;
    defparam comm_buf_0__i3_LC_15_8_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i3_LC_15_8_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_0__i3_LC_15_8_6 (
            .in0(_gnd_net_),
            .in1(N__40758),
            .in2(N__40700),
            .in3(N__53994),
            .lcout(comm_buf_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57844),
            .ce(N__42724),
            .sr(N__42852));
    defparam i6988_2_lut_LC_15_9_1.C_ON=1'b0;
    defparam i6988_2_lut_LC_15_9_1.SEQ_MODE=4'b0000;
    defparam i6988_2_lut_LC_15_9_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 i6988_2_lut_LC_15_9_1 (
            .in0(N__52390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54006),
            .lcout(n9321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_217_LC_15_9_2.C_ON=1'b0;
    defparam i1_4_lut_adj_217_LC_15_9_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_217_LC_15_9_2.LUT_INIT=16'b1000100010001100;
    LogicCell40 i1_4_lut_adj_217_LC_15_9_2 (
            .in0(N__54637),
            .in1(N__51542),
            .in2(N__51605),
            .in3(N__52393),
            .lcout(n11406),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam flagcntwd_313_LC_15_9_3.C_ON=1'b0;
    defparam flagcntwd_313_LC_15_9_3.SEQ_MODE=4'b1000;
    defparam flagcntwd_313_LC_15_9_3.LUT_INIT=16'b1100110011111111;
    LogicCell40 flagcntwd_313_LC_15_9_3 (
            .in0(_gnd_net_),
            .in1(N__54008),
            .in2(_gnd_net_),
            .in3(N__53504),
            .lcout(flagcntwd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57854),
            .ce(N__40667),
            .sr(N__51212));
    defparam i1_2_lut_3_lut_adj_301_LC_15_9_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_301_LC_15_9_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_301_LC_15_9_5.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_adj_301_LC_15_9_5 (
            .in0(N__52391),
            .in1(N__54007),
            .in2(_gnd_net_),
            .in3(N__54635),
            .lcout(n12242),
            .ltout(n12242_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_86_LC_15_9_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_86_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_86_LC_15_9_6.LUT_INIT=16'b1111000010100000;
    LogicCell40 i1_2_lut_3_lut_adj_86_LC_15_9_6 (
            .in0(N__54636),
            .in1(_gnd_net_),
            .in2(N__41108),
            .in3(N__52392),
            .lcout(n20599),
            .ltout(n20599_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_236_LC_15_9_7.C_ON=1'b0;
    defparam i1_4_lut_adj_236_LC_15_9_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_236_LC_15_9_7.LUT_INIT=16'b1011000010100000;
    LogicCell40 i1_4_lut_adj_236_LC_15_9_7 (
            .in0(N__50925),
            .in1(N__53503),
            .in2(N__41105),
            .in3(N__43238),
            .lcout(n12047),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_254_LC_15_10_0.C_ON=1'b0;
    defparam i2_3_lut_adj_254_LC_15_10_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_254_LC_15_10_0.LUT_INIT=16'b1111111101100110;
    LogicCell40 i2_3_lut_adj_254_LC_15_10_0 (
            .in0(N__47911),
            .in1(N__50552),
            .in2(_gnd_net_),
            .in3(N__47866),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i4_LC_15_10_1.C_ON=1'b0;
    defparam buf_device_acadc_i4_LC_15_10_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i4_LC_15_10_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i4_LC_15_10_1 (
            .in0(N__49449),
            .in1(N__41390),
            .in2(N__44302),
            .in3(N__41073),
            .lcout(IAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57864),
            .ce(),
            .sr(_gnd_net_));
    defparam i12241_2_lut_LC_15_10_2.C_ON=1'b0;
    defparam i12241_2_lut_LC_15_10_2.SEQ_MODE=4'b0000;
    defparam i12241_2_lut_LC_15_10_2.LUT_INIT=16'b0101010100000000;
    LogicCell40 i12241_2_lut_LC_15_10_2 (
            .in0(N__41053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41885),
            .lcout(n14663),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12360_2_lut_LC_15_10_3.C_ON=1'b0;
    defparam i12360_2_lut_LC_15_10_3.SEQ_MODE=4'b0000;
    defparam i12360_2_lut_LC_15_10_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12360_2_lut_LC_15_10_3 (
            .in0(_gnd_net_),
            .in1(N__54654),
            .in2(_gnd_net_),
            .in3(N__47029),
            .lcout(n14773),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18728_2_lut_LC_15_10_4.C_ON=1'b0;
    defparam i18728_2_lut_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam i18728_2_lut_LC_15_10_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18728_2_lut_LC_15_10_4 (
            .in0(_gnd_net_),
            .in1(N__40958),
            .in2(_gnd_net_),
            .in3(N__56324),
            .lcout(n20973),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18739_2_lut_LC_15_10_5.C_ON=1'b0;
    defparam i18739_2_lut_LC_15_10_5.SEQ_MODE=4'b0000;
    defparam i18739_2_lut_LC_15_10_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 i18739_2_lut_LC_15_10_5 (
            .in0(N__56323),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40946),
            .lcout(n20983),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i5_LC_15_10_6.C_ON=1'b0;
    defparam buf_device_acadc_i5_LC_15_10_6.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i5_LC_15_10_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_device_acadc_i5_LC_15_10_6 (
            .in0(N__41389),
            .in1(N__44127),
            .in2(N__49833),
            .in3(N__41322),
            .lcout(VAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57864),
            .ce(),
            .sr(_gnd_net_));
    defparam i18816_2_lut_LC_15_10_7.C_ON=1'b0;
    defparam i18816_2_lut_LC_15_10_7.SEQ_MODE=4'b0000;
    defparam i18816_2_lut_LC_15_10_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 i18816_2_lut_LC_15_10_7 (
            .in0(N__56322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47510),
            .lcout(n21046),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21998_bdd_4_lut_LC_15_11_0.C_ON=1'b0;
    defparam n21998_bdd_4_lut_LC_15_11_0.SEQ_MODE=4'b0000;
    defparam n21998_bdd_4_lut_LC_15_11_0.LUT_INIT=16'b1010101011100100;
    LogicCell40 n21998_bdd_4_lut_LC_15_11_0 (
            .in0(N__41204),
            .in1(N__41291),
            .in2(N__46469),
            .in3(N__49106),
            .lcout(n22001),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19385_LC_15_11_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19385_LC_15_11_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19385_LC_15_11_1.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19385_LC_15_11_1 (
            .in0(N__49105),
            .in1(N__41270),
            .in2(N__41258),
            .in3(N__48337),
            .lcout(n22004),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_0_i26_3_lut_LC_15_11_2.C_ON=1'b0;
    defparam mux_135_Mux_0_i26_3_lut_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_0_i26_3_lut_LC_15_11_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_0_i26_3_lut_LC_15_11_2 (
            .in0(N__41233),
            .in1(N__56271),
            .in2(_gnd_net_),
            .in3(N__46492),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19380_LC_15_11_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19380_LC_15_11_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19380_LC_15_11_3.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19380_LC_15_11_3 (
            .in0(N__49104),
            .in1(N__41216),
            .in2(N__41207),
            .in3(N__48336),
            .lcout(n21998),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22004_bdd_4_lut_LC_15_11_4.C_ON=1'b0;
    defparam n22004_bdd_4_lut_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam n22004_bdd_4_lut_LC_15_11_4.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22004_bdd_4_lut_LC_15_11_4 (
            .in0(N__41198),
            .in1(N__41186),
            .in2(N__52157),
            .in3(N__49107),
            .lcout(),
            .ltout(n22007_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1548473_i1_3_lut_LC_15_11_5.C_ON=1'b0;
    defparam i1548473_i1_3_lut_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam i1548473_i1_3_lut_LC_15_11_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 i1548473_i1_3_lut_LC_15_11_5 (
            .in0(_gnd_net_),
            .in1(N__48607),
            .in2(N__41180),
            .in3(N__41177),
            .lcout(),
            .ltout(n30_adj_1486_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i0_LC_15_11_6.C_ON=1'b0;
    defparam comm_buf_1__i0_LC_15_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i0_LC_15_11_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_1__i0_LC_15_11_6 (
            .in0(_gnd_net_),
            .in1(N__54051),
            .in2(N__41171),
            .in3(N__50771),
            .lcout(comm_buf_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57874),
            .ce(N__47053),
            .sr(N__46970));
    defparam n21992_bdd_4_lut_LC_15_12_0.C_ON=1'b0;
    defparam n21992_bdd_4_lut_LC_15_12_0.SEQ_MODE=4'b0000;
    defparam n21992_bdd_4_lut_LC_15_12_0.LUT_INIT=16'b1010110110101000;
    LogicCell40 n21992_bdd_4_lut_LC_15_12_0 (
            .in0(N__41591),
            .in1(N__41657),
            .in2(N__48423),
            .in3(N__49979),
            .lcout(n21995),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19390_LC_15_12_1.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19390_LC_15_12_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19390_LC_15_12_1.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19390_LC_15_12_1 (
            .in0(N__56319),
            .in1(N__41630),
            .in2(N__48365),
            .in3(N__43901),
            .lcout(n21992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18303_3_lut_LC_15_12_2.C_ON=1'b0;
    defparam i18303_3_lut_LC_15_12_2.SEQ_MODE=4'b0000;
    defparam i18303_3_lut_LC_15_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 i18303_3_lut_LC_15_12_2 (
            .in0(N__41585),
            .in1(N__56320),
            .in2(_gnd_net_),
            .in3(N__43460),
            .lcout(),
            .ltout(n20917_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18305_4_lut_LC_15_12_3.C_ON=1'b0;
    defparam i18305_4_lut_LC_15_12_3.SEQ_MODE=4'b0000;
    defparam i18305_4_lut_LC_15_12_3.LUT_INIT=16'b1110111011110000;
    LogicCell40 i18305_4_lut_LC_15_12_3 (
            .in0(N__56321),
            .in1(N__41564),
            .in2(N__41555),
            .in3(N__48408),
            .lcout(),
            .ltout(n20919_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19567_LC_15_12_4.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19567_LC_15_12_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19567_LC_15_12_4.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_2__bdd_4_lut_19567_LC_15_12_4 (
            .in0(N__49013),
            .in1(N__41552),
            .in2(N__41546),
            .in3(N__48700),
            .lcout(),
            .ltout(n22220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22220_bdd_4_lut_LC_15_12_5.C_ON=1'b0;
    defparam n22220_bdd_4_lut_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam n22220_bdd_4_lut_LC_15_12_5.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22220_bdd_4_lut_LC_15_12_5 (
            .in0(N__41543),
            .in1(N__41531),
            .in2(N__41516),
            .in3(N__48688),
            .lcout(),
            .ltout(n22223_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i0_LC_15_12_6.C_ON=1'b0;
    defparam comm_buf_0__i0_LC_15_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i0_LC_15_12_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_0__i0_LC_15_12_6 (
            .in0(_gnd_net_),
            .in1(N__54052),
            .in2(N__41513),
            .in3(N__50782),
            .lcout(comm_buf_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57887),
            .ce(N__42722),
            .sr(N__42857));
    defparam i19053_4_lut_4_lut_LC_15_12_7.C_ON=1'b0;
    defparam i19053_4_lut_4_lut_LC_15_12_7.SEQ_MODE=4'b0000;
    defparam i19053_4_lut_4_lut_LC_15_12_7.LUT_INIT=16'b1110111101101011;
    LogicCell40 i19053_4_lut_4_lut_LC_15_12_7 (
            .in0(N__56318),
            .in1(N__48687),
            .in2(N__48364),
            .in3(N__49012),
            .lcout(n21094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_cntvec_i0_i0_LC_15_13_0.C_ON=1'b1;
    defparam data_cntvec_i0_i0_LC_15_13_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i0_LC_15_13_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i0_LC_15_13_0 (
            .in0(_gnd_net_),
            .in1(N__46491),
            .in2(N__41441),
            .in3(_gnd_net_),
            .lcout(data_cntvec_0),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(n19354),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i1_LC_15_13_1.C_ON=1'b1;
    defparam data_cntvec_i0_i1_LC_15_13_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i1_LC_15_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i1_LC_15_13_1 (
            .in0(_gnd_net_),
            .in1(N__46767),
            .in2(_gnd_net_),
            .in3(N__41684),
            .lcout(data_cntvec_1),
            .ltout(),
            .carryin(n19354),
            .carryout(n19355),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i2_LC_15_13_2.C_ON=1'b1;
    defparam data_cntvec_i0_i2_LC_15_13_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i2_LC_15_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i2_LC_15_13_2 (
            .in0(_gnd_net_),
            .in1(N__46845),
            .in2(_gnd_net_),
            .in3(N__41681),
            .lcout(data_cntvec_2),
            .ltout(),
            .carryin(n19355),
            .carryout(n19356),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i3_LC_15_13_3.C_ON=1'b1;
    defparam data_cntvec_i0_i3_LC_15_13_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i3_LC_15_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i3_LC_15_13_3 (
            .in0(_gnd_net_),
            .in1(N__47730),
            .in2(_gnd_net_),
            .in3(N__41678),
            .lcout(data_cntvec_3),
            .ltout(),
            .carryin(n19356),
            .carryout(n19357),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i4_LC_15_13_4.C_ON=1'b1;
    defparam data_cntvec_i0_i4_LC_15_13_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i4_LC_15_13_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i4_LC_15_13_4 (
            .in0(_gnd_net_),
            .in1(N__46744),
            .in2(_gnd_net_),
            .in3(N__41675),
            .lcout(data_cntvec_4),
            .ltout(),
            .carryin(n19357),
            .carryout(n19358),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i5_LC_15_13_5.C_ON=1'b1;
    defparam data_cntvec_i0_i5_LC_15_13_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i5_LC_15_13_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i5_LC_15_13_5 (
            .in0(_gnd_net_),
            .in1(N__47753),
            .in2(_gnd_net_),
            .in3(N__41672),
            .lcout(data_cntvec_5),
            .ltout(),
            .carryin(n19358),
            .carryout(n19359),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i6_LC_15_13_6.C_ON=1'b1;
    defparam data_cntvec_i0_i6_LC_15_13_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i6_LC_15_13_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i6_LC_15_13_6 (
            .in0(_gnd_net_),
            .in1(N__46521),
            .in2(_gnd_net_),
            .in3(N__41669),
            .lcout(data_cntvec_6),
            .ltout(),
            .carryin(n19359),
            .carryout(n19360),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i7_LC_15_13_7.C_ON=1'b1;
    defparam data_cntvec_i0_i7_LC_15_13_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i7_LC_15_13_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i7_LC_15_13_7 (
            .in0(_gnd_net_),
            .in1(N__49225),
            .in2(_gnd_net_),
            .in3(N__41666),
            .lcout(data_cntvec_7),
            .ltout(),
            .carryin(n19360),
            .carryout(n19361),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__41887),
            .sr(N__41832));
    defparam data_cntvec_i0_i8_LC_15_14_0.C_ON=1'b1;
    defparam data_cntvec_i0_i8_LC_15_14_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i8_LC_15_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i8_LC_15_14_0 (
            .in0(_gnd_net_),
            .in1(N__43459),
            .in2(_gnd_net_),
            .in3(N__41663),
            .lcout(data_cntvec_8),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(n19362),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i9_LC_15_14_1.C_ON=1'b1;
    defparam data_cntvec_i0_i9_LC_15_14_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i9_LC_15_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i9_LC_15_14_1 (
            .in0(_gnd_net_),
            .in1(N__47530),
            .in2(_gnd_net_),
            .in3(N__41660),
            .lcout(data_cntvec_9),
            .ltout(),
            .carryin(n19362),
            .carryout(n19363),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i10_LC_15_14_2.C_ON=1'b1;
    defparam data_cntvec_i0_i10_LC_15_14_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i10_LC_15_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i10_LC_15_14_2 (
            .in0(_gnd_net_),
            .in1(N__42061),
            .in2(_gnd_net_),
            .in3(N__41906),
            .lcout(data_cntvec_10),
            .ltout(),
            .carryin(n19363),
            .carryout(n19364),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i11_LC_15_14_3.C_ON=1'b1;
    defparam data_cntvec_i0_i11_LC_15_14_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i11_LC_15_14_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i11_LC_15_14_3 (
            .in0(_gnd_net_),
            .in1(N__41785),
            .in2(_gnd_net_),
            .in3(N__41903),
            .lcout(data_cntvec_11),
            .ltout(),
            .carryin(n19364),
            .carryout(n19365),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i12_LC_15_14_4.C_ON=1'b1;
    defparam data_cntvec_i0_i12_LC_15_14_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i12_LC_15_14_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i12_LC_15_14_4 (
            .in0(_gnd_net_),
            .in1(N__42080),
            .in2(_gnd_net_),
            .in3(N__41900),
            .lcout(data_cntvec_12),
            .ltout(),
            .carryin(n19365),
            .carryout(n19366),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i13_LC_15_14_5.C_ON=1'b1;
    defparam data_cntvec_i0_i13_LC_15_14_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i13_LC_15_14_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i13_LC_15_14_5 (
            .in0(_gnd_net_),
            .in1(N__43438),
            .in2(_gnd_net_),
            .in3(N__41897),
            .lcout(data_cntvec_13),
            .ltout(),
            .carryin(n19366),
            .carryout(n19367),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i14_LC_15_14_6.C_ON=1'b1;
    defparam data_cntvec_i0_i14_LC_15_14_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i14_LC_15_14_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i14_LC_15_14_6 (
            .in0(_gnd_net_),
            .in1(N__41798),
            .in2(_gnd_net_),
            .in3(N__41894),
            .lcout(data_cntvec_14),
            .ltout(),
            .carryin(n19367),
            .carryout(n19368),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam data_cntvec_i0_i15_LC_15_14_7.C_ON=1'b0;
    defparam data_cntvec_i0_i15_LC_15_14_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i15_LC_15_14_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i15_LC_15_14_7 (
            .in0(_gnd_net_),
            .in1(N__47485),
            .in2(_gnd_net_),
            .in3(N__41891),
            .lcout(data_cntvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__41888),
            .sr(N__41828));
    defparam i7_4_lut_adj_182_LC_15_15_0.C_ON=1'b0;
    defparam i7_4_lut_adj_182_LC_15_15_0.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_182_LC_15_15_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_adj_182_LC_15_15_0 (
            .in0(N__41797),
            .in1(N__41784),
            .in2(N__44536),
            .in3(N__41763),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6414_3_lut_LC_15_15_1.C_ON=1'b0;
    defparam i6414_3_lut_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam i6414_3_lut_LC_15_15_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6414_3_lut_LC_15_15_1 (
            .in0(N__52489),
            .in1(N__41949),
            .in2(_gnd_net_),
            .in3(N__41750),
            .lcout(n8_adj_1559),
            .ltout(n8_adj_1559_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_6_i15_4_lut_LC_15_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_6_i15_4_lut_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_6_i15_4_lut_LC_15_15_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 comm_state_3__I_0_365_Mux_6_i15_4_lut_LC_15_15_2 (
            .in0(N__41983),
            .in1(N__54868),
            .in2(N__42305),
            .in3(N__49521),
            .lcout(data_index_9_N_216_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_365_Mux_1_i15_4_lut_LC_15_15_3.C_ON=1'b0;
    defparam comm_state_3__I_0_365_Mux_1_i15_4_lut_LC_15_15_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_365_Mux_1_i15_4_lut_LC_15_15_3.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_365_Mux_1_i15_4_lut_LC_15_15_3 (
            .in0(N__54867),
            .in1(N__42212),
            .in2(N__49629),
            .in3(N__42199),
            .lcout(data_index_9_N_216_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i2_LC_15_15_4.C_ON=1'b0;
    defparam acadc_skipCount_i2_LC_15_15_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i2_LC_15_15_4.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i2_LC_15_15_4 (
            .in0(N__47135),
            .in1(N__49366),
            .in2(N__46288),
            .in3(N__49522),
            .lcout(acadc_skipCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57928),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_184_LC_15_15_5.C_ON=1'b0;
    defparam i5_4_lut_adj_184_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_184_LC_15_15_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i5_4_lut_adj_184_LC_15_15_5 (
            .in0(N__42079),
            .in1(N__42060),
            .in2(N__42040),
            .in3(N__42009),
            .lcout(n21_adj_1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i6_LC_15_15_6.C_ON=1'b0;
    defparam data_index_i6_LC_15_15_6.SEQ_MODE=4'b1000;
    defparam data_index_i6_LC_15_15_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 data_index_i6_LC_15_15_6 (
            .in0(N__41993),
            .in1(N__54869),
            .in2(N__41987),
            .in3(N__49523),
            .lcout(data_index_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57928),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_15_15_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_15_15_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \comm_spi.RESET_I_0_96_2_lut_LC_15_15_7  (
            .in0(N__56852),
            .in1(N__55311),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_771 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_cnt_3772_3773__i1_LC_15_16_0.C_ON=1'b1;
    defparam clk_cnt_3772_3773__i1_LC_15_16_0.SEQ_MODE=4'b1000;
    defparam clk_cnt_3772_3773__i1_LC_15_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3772_3773__i1_LC_15_16_0 (
            .in0(_gnd_net_),
            .in1(N__42512),
            .in2(_gnd_net_),
            .in3(N__41915),
            .lcout(clk_cnt_0),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(n19505),
            .clk(N__45083),
            .ce(),
            .sr(N__43838));
    defparam clk_cnt_3772_3773__i2_LC_15_16_1.C_ON=1'b1;
    defparam clk_cnt_3772_3773__i2_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam clk_cnt_3772_3773__i2_LC_15_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3772_3773__i2_LC_15_16_1 (
            .in0(_gnd_net_),
            .in1(N__42487),
            .in2(_gnd_net_),
            .in3(N__41912),
            .lcout(clk_cnt_1),
            .ltout(),
            .carryin(n19505),
            .carryout(n19506),
            .clk(N__45083),
            .ce(),
            .sr(N__43838));
    defparam clk_cnt_3772_3773__i3_LC_15_16_2.C_ON=1'b1;
    defparam clk_cnt_3772_3773__i3_LC_15_16_2.SEQ_MODE=4'b1000;
    defparam clk_cnt_3772_3773__i3_LC_15_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3772_3773__i3_LC_15_16_2 (
            .in0(_gnd_net_),
            .in1(N__42457),
            .in2(_gnd_net_),
            .in3(N__41909),
            .lcout(clk_cnt_2),
            .ltout(),
            .carryin(n19506),
            .carryout(n19507),
            .clk(N__45083),
            .ce(),
            .sr(N__43838));
    defparam clk_cnt_3772_3773__i4_LC_15_16_3.C_ON=1'b1;
    defparam clk_cnt_3772_3773__i4_LC_15_16_3.SEQ_MODE=4'b1000;
    defparam clk_cnt_3772_3773__i4_LC_15_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3772_3773__i4_LC_15_16_3 (
            .in0(_gnd_net_),
            .in1(N__42473),
            .in2(_gnd_net_),
            .in3(N__42518),
            .lcout(clk_cnt_3),
            .ltout(),
            .carryin(n19507),
            .carryout(n19508),
            .clk(N__45083),
            .ce(),
            .sr(N__43838));
    defparam clk_cnt_3772_3773__i5_LC_15_16_4.C_ON=1'b0;
    defparam clk_cnt_3772_3773__i5_LC_15_16_4.SEQ_MODE=4'b1000;
    defparam clk_cnt_3772_3773__i5_LC_15_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_cnt_3772_3773__i5_LC_15_16_4 (
            .in0(_gnd_net_),
            .in1(N__42500),
            .in2(_gnd_net_),
            .in3(N__42515),
            .lcout(clk_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45083),
            .ce(),
            .sr(N__43838));
    defparam i1_2_lut_adj_232_LC_15_17_0.C_ON=1'b0;
    defparam i1_2_lut_adj_232_LC_15_17_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_232_LC_15_17_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_adj_232_LC_15_17_0 (
            .in0(N__42511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42499),
            .lcout(),
            .ltout(n6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_234_LC_15_17_1.C_ON=1'b0;
    defparam i4_4_lut_adj_234_LC_15_17_1.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_234_LC_15_17_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_adj_234_LC_15_17_1 (
            .in0(N__42488),
            .in1(N__42472),
            .in2(N__42461),
            .in3(N__42458),
            .lcout(n14730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_3_i23_3_lut_LC_15_17_4.C_ON=1'b0;
    defparam mux_134_Mux_3_i23_3_lut_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_3_i23_3_lut_LC_15_17_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_134_Mux_3_i23_3_lut_LC_15_17_4 (
            .in0(N__44197),
            .in1(N__56334),
            .in2(_gnd_net_),
            .in3(N__42443),
            .lcout(n23_adj_1540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_15_17_5.C_ON=1'b0;
    defparam i5_4_lut_LC_15_17_5.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_15_17_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_15_17_5 (
            .in0(N__42415),
            .in1(N__42403),
            .in2(N__42392),
            .in3(N__42376),
            .lcout(),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_165_LC_15_17_6.C_ON=1'b0;
    defparam i6_4_lut_adj_165_LC_15_17_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_165_LC_15_17_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_165_LC_15_17_6 (
            .in0(N__42364),
            .in1(N__42352),
            .in2(N__42341),
            .in3(N__42337),
            .lcout(n20543),
            .ltout(n20543_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclk_304_LC_15_17_7.C_ON=1'b0;
    defparam dds0_mclk_304_LC_15_17_7.SEQ_MODE=4'b1000;
    defparam dds0_mclk_304_LC_15_17_7.LUT_INIT=16'b1100001111001100;
    LogicCell40 dds0_mclk_304_LC_15_17_7 (
            .in0(_gnd_net_),
            .in1(N__45028),
            .in2(N__42320),
            .in3(N__42317),
            .lcout(dds0_mclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclk_304C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i3_LC_15_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i3_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i3_LC_15_18_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \SIG_DDS.bit_cnt_i3_LC_15_18_0  (
            .in0(N__44753),
            .in1(N__44845),
            .in2(N__44870),
            .in3(N__44828),
            .lcout(\SIG_DDS.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57960),
            .ce(N__50176),
            .sr(N__44765));
    defparam \SIG_DDS.bit_cnt_i1_LC_15_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i1_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i1_LC_15_18_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.bit_cnt_i1_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__44862),
            .in2(_gnd_net_),
            .in3(N__44751),
            .lcout(\SIG_DDS.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57960),
            .ce(N__50176),
            .sr(N__44765));
    defparam \SIG_DDS.bit_cnt_i2_LC_15_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i2_LC_15_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i2_LC_15_18_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \SIG_DDS.bit_cnt_i2_LC_15_18_2  (
            .in0(N__44752),
            .in1(_gnd_net_),
            .in2(N__44869),
            .in3(N__44844),
            .lcout(\SIG_DDS.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57960),
            .ce(N__50176),
            .sr(N__44765));
    defparam \SIG_DDS.dds_state_i2_LC_15_19_2 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i2_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i2_LC_15_19_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \SIG_DDS.dds_state_i2_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__50233),
            .in2(_gnd_net_),
            .in3(N__50156),
            .lcout(dds_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57964),
            .ce(),
            .sr(_gnd_net_));
    defparam i18840_2_lut_LC_16_2_2.C_ON=1'b0;
    defparam i18840_2_lut_LC_16_2_2.SEQ_MODE=4'b0000;
    defparam i18840_2_lut_LC_16_2_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18840_2_lut_LC_16_2_2 (
            .in0(_gnd_net_),
            .in1(N__42638),
            .in2(_gnd_net_),
            .in3(N__56370),
            .lcout(n21038),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.bit_cnt_3778__i3_LC_16_4_0 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3778__i3_LC_16_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3778__i3_LC_16_4_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \comm_spi.bit_cnt_3778__i3_LC_16_4_0  (
            .in0(N__42575),
            .in1(N__42610),
            .in2(N__42542),
            .in3(N__42560),
            .lcout(\comm_spi.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3778__i3C_net ),
            .ce(),
            .sr(N__56823));
    defparam \comm_spi.bit_cnt_3778__i2_LC_16_4_1 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3778__i2_LC_16_4_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3778__i2_LC_16_4_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \comm_spi.bit_cnt_3778__i2_LC_16_4_1  (
            .in0(N__42559),
            .in1(N__42538),
            .in2(_gnd_net_),
            .in3(N__42574),
            .lcout(\comm_spi.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3778__i3C_net ),
            .ce(),
            .sr(N__56823));
    defparam \comm_spi.bit_cnt_3778__i1_LC_16_4_2 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3778__i1_LC_16_4_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3778__i1_LC_16_4_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \comm_spi.bit_cnt_3778__i1_LC_16_4_2  (
            .in0(N__42537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42558),
            .lcout(\comm_spi.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3778__i3C_net ),
            .ce(),
            .sr(N__56823));
    defparam \comm_spi.bit_cnt_3778__i0_LC_16_4_3 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3778__i0_LC_16_4_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3778__i0_LC_16_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \comm_spi.bit_cnt_3778__i0_LC_16_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42536),
            .lcout(\comm_spi.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3778__i3C_net ),
            .ce(),
            .sr(N__56823));
    defparam comm_buf_0__i7_LC_16_5_0.C_ON=1'b0;
    defparam comm_buf_0__i7_LC_16_5_0.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i7_LC_16_5_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i7_LC_16_5_0 (
            .in0(N__51342),
            .in1(N__54035),
            .in2(_gnd_net_),
            .in3(N__42893),
            .lcout(comm_buf_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57826),
            .ce(N__42721),
            .sr(N__42847));
    defparam comm_buf_0__i5_LC_16_5_1.C_ON=1'b0;
    defparam comm_buf_0__i5_LC_16_5_1.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i5_LC_16_5_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i5_LC_16_5_1 (
            .in0(N__54033),
            .in1(N__50995),
            .in2(_gnd_net_),
            .in3(N__42878),
            .lcout(comm_buf_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57826),
            .ce(N__42721),
            .sr(N__42847));
    defparam comm_buf_0__i1_LC_16_5_2.C_ON=1'b0;
    defparam comm_buf_0__i1_LC_16_5_2.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i1_LC_16_5_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i1_LC_16_5_2 (
            .in0(N__45322),
            .in1(N__54034),
            .in2(_gnd_net_),
            .in3(N__44003),
            .lcout(comm_buf_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57826),
            .ce(N__42721),
            .sr(N__42847));
    defparam i18822_2_lut_LC_16_6_0.C_ON=1'b0;
    defparam i18822_2_lut_LC_16_6_0.SEQ_MODE=4'b0000;
    defparam i18822_2_lut_LC_16_6_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18822_2_lut_LC_16_6_0 (
            .in0(_gnd_net_),
            .in1(N__45742),
            .in2(_gnd_net_),
            .in3(N__53518),
            .lcout(),
            .ltout(n21199_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i3_LC_16_6_1.C_ON=1'b0;
    defparam comm_state_i3_LC_16_6_1.SEQ_MODE=4'b1000;
    defparam comm_state_i3_LC_16_6_1.LUT_INIT=16'b0011000001010101;
    LogicCell40 comm_state_i3_LC_16_6_1 (
            .in0(N__45221),
            .in1(N__49626),
            .in2(N__42791),
            .in3(N__54559),
            .lcout(comm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57835),
            .ce(N__45749),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_16_6_2.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_16_6_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_16_6_2.LUT_INIT=16'b1100110011011100;
    LogicCell40 i1_3_lut_4_lut_LC_16_6_2 (
            .in0(N__54029),
            .in1(N__50885),
            .in2(N__45205),
            .in3(N__53516),
            .lcout(n11869),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_105_LC_16_6_5.C_ON=1'b0;
    defparam i1_2_lut_adj_105_LC_16_6_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_105_LC_16_6_5.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_105_LC_16_6_5 (
            .in0(_gnd_net_),
            .in1(N__52259),
            .in2(_gnd_net_),
            .in3(N__54558),
            .lcout(n20681),
            .ltout(n20681_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_adj_129_LC_16_6_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_adj_129_LC_16_6_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_adj_129_LC_16_6_6.LUT_INIT=16'b1111110011111110;
    LogicCell40 i1_2_lut_3_lut_4_lut_adj_129_LC_16_6_6 (
            .in0(N__45201),
            .in1(N__53862),
            .in2(N__42788),
            .in3(N__53517),
            .lcout(),
            .ltout(n12108_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_233_LC_16_6_7.C_ON=1'b0;
    defparam i1_4_lut_adj_233_LC_16_6_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_233_LC_16_6_7.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_233_LC_16_6_7 (
            .in0(N__50886),
            .in1(N__42778),
            .in2(N__42734),
            .in3(N__42731),
            .lcout(n11977),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_6_i2_3_lut_LC_16_7_0.C_ON=1'b0;
    defparam mux_143_Mux_6_i2_3_lut_LC_16_7_0.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_6_i2_3_lut_LC_16_7_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_143_Mux_6_i2_3_lut_LC_16_7_0 (
            .in0(N__54344),
            .in1(N__42659),
            .in2(_gnd_net_),
            .in3(N__42647),
            .lcout(n2_adj_1584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19041_2_lut_LC_16_7_1.C_ON=1'b0;
    defparam i19041_2_lut_LC_16_7_1.SEQ_MODE=4'b0000;
    defparam i19041_2_lut_LC_16_7_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19041_2_lut_LC_16_7_1 (
            .in0(_gnd_net_),
            .in1(N__43205),
            .in2(_gnd_net_),
            .in3(N__54345),
            .lcout(),
            .ltout(n21329_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19489_LC_16_7_2.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19489_LC_16_7_2.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19489_LC_16_7_2.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_1__bdd_4_lut_19489_LC_16_7_2 (
            .in0(N__50547),
            .in1(N__54191),
            .in2(N__43187),
            .in3(N__50682),
            .lcout(),
            .ltout(n21986_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i6_LC_16_7_3.C_ON=1'b0;
    defparam comm_tx_buf_i6_LC_16_7_3.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i6_LC_16_7_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i6_LC_16_7_3 (
            .in0(N__50683),
            .in1(N__43079),
            .in2(N__43184),
            .in3(N__43181),
            .lcout(comm_tx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57845),
            .ce(N__46213),
            .sr(N__46116));
    defparam mux_143_Mux_6_i1_3_lut_LC_16_7_5.C_ON=1'b0;
    defparam mux_143_Mux_6_i1_3_lut_LC_16_7_5.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_6_i1_3_lut_LC_16_7_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_143_Mux_6_i1_3_lut_LC_16_7_5 (
            .in0(N__43136),
            .in1(N__52505),
            .in2(_gnd_net_),
            .in3(N__54343),
            .lcout(n1_adj_1583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_295_LC_16_7_6.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_295_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_295_LC_16_7_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 i2_2_lut_3_lut_adj_295_LC_16_7_6 (
            .in0(N__50546),
            .in1(N__43063),
            .in2(_gnd_net_),
            .in3(N__50681),
            .lcout(),
            .ltout(n7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_156_LC_16_7_7.C_ON=1'b0;
    defparam i1_4_lut_adj_156_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_156_LC_16_7_7.LUT_INIT=16'b1100110010000000;
    LogicCell40 i1_4_lut_adj_156_LC_16_7_7 (
            .in0(N__45764),
            .in1(N__51568),
            .in2(N__43043),
            .in3(N__54530),
            .lcout(n12244),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19419_LC_16_8_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19419_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19419_LC_16_8_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_19419_LC_16_8_0 (
            .in0(N__54270),
            .in1(N__43040),
            .in2(N__43025),
            .in3(N__50482),
            .lcout(),
            .ltout(n22046_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22046_bdd_4_lut_LC_16_8_1.C_ON=1'b0;
    defparam n22046_bdd_4_lut_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam n22046_bdd_4_lut_LC_16_8_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22046_bdd_4_lut_LC_16_8_1 (
            .in0(N__50483),
            .in1(N__42972),
            .in2(N__42896),
            .in3(N__47134),
            .lcout(n22049),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_2_i4_3_lut_LC_16_8_2.C_ON=1'b0;
    defparam mux_143_Mux_2_i4_3_lut_LC_16_8_2.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_2_i4_3_lut_LC_16_8_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_143_Mux_2_i4_3_lut_LC_16_8_2 (
            .in0(N__54271),
            .in1(N__43328),
            .in2(_gnd_net_),
            .in3(N__43316),
            .lcout(),
            .ltout(n4_adj_1593_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18187_4_lut_LC_16_8_3.C_ON=1'b0;
    defparam i18187_4_lut_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam i18187_4_lut_LC_16_8_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18187_4_lut_LC_16_8_3 (
            .in0(N__50484),
            .in1(N__43307),
            .in2(N__43283),
            .in3(N__54272),
            .lcout(),
            .ltout(n20801_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i2_LC_16_8_4.C_ON=1'b0;
    defparam comm_tx_buf_i2_LC_16_8_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i2_LC_16_8_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 comm_tx_buf_i2_LC_16_8_4 (
            .in0(_gnd_net_),
            .in1(N__43280),
            .in2(N__43274),
            .in3(N__50636),
            .lcout(comm_tx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57855),
            .ce(N__46205),
            .sr(N__46133));
    defparam i18878_3_lut_LC_16_8_5.C_ON=1'b0;
    defparam i18878_3_lut_LC_16_8_5.SEQ_MODE=4'b0000;
    defparam i18878_3_lut_LC_16_8_5.LUT_INIT=16'b0100010000000000;
    LogicCell40 i18878_3_lut_LC_16_8_5 (
            .in0(N__50481),
            .in1(N__54269),
            .in2(_gnd_net_),
            .in3(N__43264),
            .lcout(),
            .ltout(n21092_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i45_4_lut_LC_16_8_6.C_ON=1'b0;
    defparam i45_4_lut_LC_16_8_6.SEQ_MODE=4'b0000;
    defparam i45_4_lut_LC_16_8_6.LUT_INIT=16'b1111000010001000;
    LogicCell40 i45_4_lut_LC_16_8_6 (
            .in0(N__43253),
            .in1(N__45194),
            .in2(N__43241),
            .in3(N__53917),
            .lcout(n20_adj_1610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i0_LC_16_9_1.C_ON=1'b0;
    defparam comm_state_i0_LC_16_9_1.SEQ_MODE=4'b1000;
    defparam comm_state_i0_LC_16_9_1.LUT_INIT=16'b0101010111001100;
    LogicCell40 comm_state_i0_LC_16_9_1 (
            .in0(N__49448),
            .in1(N__43232),
            .in2(_gnd_net_),
            .in3(N__54705),
            .lcout(comm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57865),
            .ce(N__45671),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_308_LC_16_9_2.C_ON=1'b0;
    defparam i1_2_lut_adj_308_LC_16_9_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_308_LC_16_9_2.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_308_LC_16_9_2 (
            .in0(_gnd_net_),
            .in1(N__53770),
            .in2(_gnd_net_),
            .in3(N__53495),
            .lcout(),
            .ltout(n20695_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_292_LC_16_9_3.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_292_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_292_LC_16_9_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i2_3_lut_4_lut_adj_292_LC_16_9_3 (
            .in0(N__50906),
            .in1(N__51827),
            .in2(N__43220),
            .in3(N__51670),
            .lcout(n20697),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18267_3_lut_LC_16_9_4.C_ON=1'b0;
    defparam i18267_3_lut_LC_16_9_4.SEQ_MODE=4'b0000;
    defparam i18267_3_lut_LC_16_9_4.LUT_INIT=16'b1100110010111011;
    LogicCell40 i18267_3_lut_LC_16_9_4 (
            .in0(N__51825),
            .in1(N__53771),
            .in2(_gnd_net_),
            .in3(N__53496),
            .lcout(n20881),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_16_9_5.C_ON=1'b0;
    defparam i2_2_lut_LC_16_9_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_16_9_5.LUT_INIT=16'b1111111101010101;
    LogicCell40 i2_2_lut_LC_16_9_5 (
            .in0(N__53497),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51826),
            .lcout(n14545),
            .ltout(n14545_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_306_LC_16_9_6.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_306_LC_16_9_6.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_306_LC_16_9_6.LUT_INIT=16'b1111111111111101;
    LogicCell40 i2_3_lut_4_lut_adj_306_LC_16_9_6 (
            .in0(N__51671),
            .in1(N__53772),
            .in2(N__43424),
            .in3(N__50907),
            .lcout(n11420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i7_LC_16_10_0.C_ON=1'b0;
    defparam comm_buf_1__i7_LC_16_10_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i7_LC_16_10_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i7_LC_16_10_0 (
            .in0(N__51394),
            .in1(N__54026),
            .in2(_gnd_net_),
            .in3(N__43850),
            .lcout(comm_buf_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57875),
            .ce(N__47061),
            .sr(N__46989));
    defparam mux_135_Mux_1_i26_3_lut_LC_16_11_0.C_ON=1'b0;
    defparam mux_135_Mux_1_i26_3_lut_LC_16_11_0.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_1_i26_3_lut_LC_16_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_1_i26_3_lut_LC_16_11_0 (
            .in0(N__43420),
            .in1(N__56329),
            .in2(_gnd_net_),
            .in3(N__46768),
            .lcout(),
            .ltout(n26_adj_1522_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19547_LC_16_11_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19547_LC_16_11_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19547_LC_16_11_1.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19547_LC_16_11_1 (
            .in0(N__45839),
            .in1(N__48339),
            .in2(N__43403),
            .in3(N__49114),
            .lcout(),
            .ltout(n22190_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22190_bdd_4_lut_LC_16_11_2.C_ON=1'b0;
    defparam n22190_bdd_4_lut_LC_16_11_2.SEQ_MODE=4'b0000;
    defparam n22190_bdd_4_lut_LC_16_11_2.LUT_INIT=16'b1111001011000010;
    LogicCell40 n22190_bdd_4_lut_LC_16_11_2 (
            .in0(N__43400),
            .in1(N__49115),
            .in2(N__43376),
            .in3(N__46694),
            .lcout(),
            .ltout(n22193_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1546061_i1_3_lut_LC_16_11_3.C_ON=1'b0;
    defparam i1546061_i1_3_lut_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam i1546061_i1_3_lut_LC_16_11_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1546061_i1_3_lut_LC_16_11_3 (
            .in0(_gnd_net_),
            .in1(N__43607),
            .in2(N__43373),
            .in3(N__48727),
            .lcout(),
            .ltout(n30_adj_1523_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i1_LC_16_11_4.C_ON=1'b0;
    defparam comm_buf_1__i1_LC_16_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i1_LC_16_11_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i1_LC_16_11_4 (
            .in0(_gnd_net_),
            .in1(N__45372),
            .in2(N__43370),
            .in3(N__54053),
            .lcout(comm_buf_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57888),
            .ce(N__47070),
            .sr(N__46993));
    defparam comm_cmd_1__bdd_4_lut_19434_LC_16_11_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19434_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19434_LC_16_11_5.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19434_LC_16_11_5 (
            .in0(N__43367),
            .in1(N__48338),
            .in2(N__43352),
            .in3(N__49112),
            .lcout(),
            .ltout(n22064_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22064_bdd_4_lut_LC_16_11_6.C_ON=1'b0;
    defparam n22064_bdd_4_lut_LC_16_11_6.SEQ_MODE=4'b0000;
    defparam n22064_bdd_4_lut_LC_16_11_6.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22064_bdd_4_lut_LC_16_11_6 (
            .in0(N__49113),
            .in1(N__52609),
            .in2(N__43625),
            .in3(N__43622),
            .lcout(n22067),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19499_LC_16_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19499_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19499_LC_16_12_0.LUT_INIT=16'b1011110010110000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19499_LC_16_12_0 (
            .in0(N__43601),
            .in1(N__49109),
            .in2(N__48425),
            .in3(N__46619),
            .lcout(),
            .ltout(n22142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22142_bdd_4_lut_LC_16_12_1.C_ON=1'b0;
    defparam n22142_bdd_4_lut_LC_16_12_1.SEQ_MODE=4'b0000;
    defparam n22142_bdd_4_lut_LC_16_12_1.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22142_bdd_4_lut_LC_16_12_1 (
            .in0(N__49110),
            .in1(N__43583),
            .in2(N__43547),
            .in3(N__43544),
            .lcout(n22145),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22130_bdd_4_lut_LC_16_12_2.C_ON=1'b0;
    defparam n22130_bdd_4_lut_LC_16_12_2.SEQ_MODE=4'b0000;
    defparam n22130_bdd_4_lut_LC_16_12_2.LUT_INIT=16'b1011100110101000;
    LogicCell40 n22130_bdd_4_lut_LC_16_12_2 (
            .in0(N__43466),
            .in1(N__49111),
            .in2(N__47291),
            .in3(N__43529),
            .lcout(),
            .ltout(n22133_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1549076_i1_3_lut_LC_16_12_3.C_ON=1'b0;
    defparam i1549076_i1_3_lut_LC_16_12_3.SEQ_MODE=4'b0000;
    defparam i1549076_i1_3_lut_LC_16_12_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1549076_i1_3_lut_LC_16_12_3 (
            .in0(_gnd_net_),
            .in1(N__43502),
            .in2(N__43496),
            .in3(N__48702),
            .lcout(),
            .ltout(n30_adj_1499_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i5_LC_16_12_4.C_ON=1'b0;
    defparam comm_buf_1__i5_LC_16_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i5_LC_16_12_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i5_LC_16_12_4 (
            .in0(_gnd_net_),
            .in1(N__51054),
            .in2(N__43493),
            .in3(N__54054),
            .lcout(comm_buf_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57900),
            .ce(N__47068),
            .sr(N__46994));
    defparam mux_135_Mux_5_i26_3_lut_LC_16_12_5.C_ON=1'b0;
    defparam mux_135_Mux_5_i26_3_lut_LC_16_12_5.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_5_i26_3_lut_LC_16_12_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_5_i26_3_lut_LC_16_12_5 (
            .in0(N__43490),
            .in1(N__56325),
            .in2(_gnd_net_),
            .in3(N__47745),
            .lcout(),
            .ltout(n26_adj_1498_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19494_LC_16_12_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19494_LC_16_12_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19494_LC_16_12_6.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19494_LC_16_12_6 (
            .in0(N__52541),
            .in1(N__48295),
            .in2(N__43469),
            .in3(N__49108),
            .lcout(n22130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_189_LC_16_13_0.C_ON=1'b0;
    defparam i3_4_lut_adj_189_LC_16_13_0.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_189_LC_16_13_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i3_4_lut_adj_189_LC_16_13_0 (
            .in0(N__43458),
            .in1(N__47547),
            .in2(N__43439),
            .in3(N__43899),
            .lcout(),
            .ltout(n19_adj_1597_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_adj_194_LC_16_13_1.C_ON=1'b0;
    defparam i13_4_lut_adj_194_LC_16_13_1.SEQ_MODE=4'b0000;
    defparam i13_4_lut_adj_194_LC_16_13_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_adj_194_LC_16_13_1 (
            .in0(N__46445),
            .in1(N__47687),
            .in2(N__43931),
            .in3(N__46676),
            .lcout(),
            .ltout(n29_adj_1635_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_196_LC_16_13_2.C_ON=1'b0;
    defparam i1_3_lut_adj_196_LC_16_13_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_196_LC_16_13_2.LUT_INIT=16'b1100110011001111;
    LogicCell40 i1_3_lut_adj_196_LC_16_13_2 (
            .in0(_gnd_net_),
            .in1(N__44897),
            .in2(N__43928),
            .in3(N__44354),
            .lcout(n16_adj_1623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i8_LC_16_13_3.C_ON=1'b0;
    defparam req_data_cnt_i8_LC_16_13_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i8_LC_16_13_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 req_data_cnt_i8_LC_16_13_3 (
            .in0(N__43900),
            .in1(_gnd_net_),
            .in2(N__44489),
            .in3(N__47397),
            .lcout(req_data_cnt_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57917),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_stop_339_LC_16_13_5.C_ON=1'b0;
    defparam eis_stop_339_LC_16_13_5.SEQ_MODE=4'b1000;
    defparam eis_stop_339_LC_16_13_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 eis_stop_339_LC_16_13_5 (
            .in0(N__44898),
            .in1(N__45536),
            .in2(_gnd_net_),
            .in3(N__43886),
            .lcout(eis_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57917),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i4_LC_16_13_6.C_ON=1'b0;
    defparam req_data_cnt_i4_LC_16_13_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i4_LC_16_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i4_LC_16_13_6 (
            .in0(N__47396),
            .in1(N__51118),
            .in2(_gnd_net_),
            .in3(N__46716),
            .lcout(req_data_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57917),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i2_LC_16_13_7.C_ON=1'b0;
    defparam req_data_cnt_i2_LC_16_13_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i2_LC_16_13_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i2_LC_16_13_7 (
            .in0(N__44050),
            .in1(N__47395),
            .in2(_gnd_net_),
            .in3(N__46310),
            .lcout(req_data_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57917),
            .ce(),
            .sr(_gnd_net_));
    defparam n22058_bdd_4_lut_LC_16_14_0.C_ON=1'b0;
    defparam n22058_bdd_4_lut_LC_16_14_0.SEQ_MODE=4'b0000;
    defparam n22058_bdd_4_lut_LC_16_14_0.LUT_INIT=16'b1110111000110000;
    LogicCell40 n22058_bdd_4_lut_LC_16_14_0 (
            .in0(N__43862),
            .in1(N__48735),
            .in2(N__44921),
            .in3(N__49187),
            .lcout(n22061),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_RTD_297_LC_16_14_2.C_ON=1'b0;
    defparam clk_RTD_297_LC_16_14_2.SEQ_MODE=4'b1000;
    defparam clk_RTD_297_LC_16_14_2.LUT_INIT=16'b0101010110101010;
    LogicCell40 clk_RTD_297_LC_16_14_2 (
            .in0(N__43656),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43837),
            .lcout(clk_RTD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45080),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_181_LC_16_14_3.C_ON=1'b0;
    defparam i6_4_lut_adj_181_LC_16_14_3.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_181_LC_16_14_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i6_4_lut_adj_181_LC_16_14_3 (
            .in0(N__46849),
            .in1(N__49224),
            .in2(N__49157),
            .in3(N__46308),
            .lcout(),
            .ltout(n22_adj_1568_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_192_LC_16_14_4.C_ON=1'b0;
    defparam i14_4_lut_adj_192_LC_16_14_4.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_192_LC_16_14_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_192_LC_16_14_4 (
            .in0(N__44369),
            .in1(N__44363),
            .in2(N__44357),
            .in3(N__47468),
            .lcout(n30_adj_1641),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18198_3_lut_LC_16_14_5.C_ON=1'b0;
    defparam i18198_3_lut_LC_16_14_5.SEQ_MODE=4'b0000;
    defparam i18198_3_lut_LC_16_14_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18198_3_lut_LC_16_14_5 (
            .in0(N__56335),
            .in1(N__44348),
            .in2(_gnd_net_),
            .in3(N__47526),
            .lcout(),
            .ltout(n20812_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18200_4_lut_LC_16_14_6.C_ON=1'b0;
    defparam i18200_4_lut_LC_16_14_6.SEQ_MODE=4'b0000;
    defparam i18200_4_lut_LC_16_14_6.LUT_INIT=16'b1111110010111000;
    LogicCell40 i18200_4_lut_LC_16_14_6 (
            .in0(N__44327),
            .in1(N__48285),
            .in2(N__44312),
            .in3(N__56336),
            .lcout(n20814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i3_LC_16_15_0.C_ON=1'b0;
    defparam buf_control_i3_LC_16_15_0.SEQ_MODE=4'b1000;
    defparam buf_control_i3_LC_16_15_0.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i3_LC_16_15_0 (
            .in0(N__49739),
            .in1(N__44441),
            .in2(N__44303),
            .in3(N__44193),
            .lcout(SELIRNG1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57941),
            .ce(),
            .sr(_gnd_net_));
    defparam i15254_2_lut_3_lut_LC_16_15_1.C_ON=1'b0;
    defparam i15254_2_lut_3_lut_LC_16_15_1.SEQ_MODE=4'b0000;
    defparam i15254_2_lut_3_lut_LC_16_15_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15254_2_lut_3_lut_LC_16_15_1 (
            .in0(N__54129),
            .in1(N__44139),
            .in2(_gnd_net_),
            .in3(N__52409),
            .lcout(n14_adj_1571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15261_2_lut_3_lut_LC_16_15_2.C_ON=1'b0;
    defparam i15261_2_lut_3_lut_LC_16_15_2.SEQ_MODE=4'b0000;
    defparam i15261_2_lut_3_lut_LC_16_15_2.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15261_2_lut_3_lut_LC_16_15_2 (
            .in0(N__52408),
            .in1(N__47133),
            .in2(_gnd_net_),
            .in3(N__54128),
            .lcout(n14_adj_1549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_LC_16_15_3.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_LC_16_15_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_LC_16_15_3.LUT_INIT=16'b1110101001001010;
    LogicCell40 comm_cmd_2__bdd_4_lut_LC_16_15_3 (
            .in0(N__49124),
            .in1(N__44594),
            .in2(N__48743),
            .in3(N__44024),
            .lcout(),
            .ltout(n22232_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22232_bdd_4_lut_LC_16_15_4.C_ON=1'b0;
    defparam n22232_bdd_4_lut_LC_16_15_4.SEQ_MODE=4'b0000;
    defparam n22232_bdd_4_lut_LC_16_15_4.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22232_bdd_4_lut_LC_16_15_4 (
            .in0(N__44018),
            .in1(N__44666),
            .in2(N__44006),
            .in3(N__48734),
            .lcout(n22235),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22226_bdd_4_lut_LC_16_15_5.C_ON=1'b0;
    defparam n22226_bdd_4_lut_LC_16_15_5.SEQ_MODE=4'b0000;
    defparam n22226_bdd_4_lut_LC_16_15_5.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22226_bdd_4_lut_LC_16_15_5 (
            .in0(N__48384),
            .in1(N__43991),
            .in2(N__43960),
            .in3(N__44681),
            .lcout(n22229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22034_bdd_4_lut_LC_16_16_0.C_ON=1'b0;
    defparam n22034_bdd_4_lut_LC_16_16_0.SEQ_MODE=4'b0000;
    defparam n22034_bdd_4_lut_LC_16_16_0.LUT_INIT=16'b1011101010011000;
    LogicCell40 n22034_bdd_4_lut_LC_16_16_0 (
            .in0(N__44879),
            .in1(N__48370),
            .in2(N__44653),
            .in3(N__44615),
            .lcout(n22037),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_7_i16_3_lut_LC_16_16_1.C_ON=1'b0;
    defparam mux_135_Mux_7_i16_3_lut_LC_16_16_1.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_7_i16_3_lut_LC_16_16_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_7_i16_3_lut_LC_16_16_1 (
            .in0(N__44587),
            .in1(N__44563),
            .in2(_gnd_net_),
            .in3(N__56331),
            .lcout(n16_adj_1503),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18222_4_lut_LC_16_16_2.C_ON=1'b0;
    defparam i18222_4_lut_LC_16_16_2.SEQ_MODE=4'b0000;
    defparam i18222_4_lut_LC_16_16_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 i18222_4_lut_LC_16_16_2 (
            .in0(N__56332),
            .in1(N__48371),
            .in2(N__44540),
            .in3(N__44507),
            .lcout(n20836),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i0_LC_16_16_3.C_ON=1'b0;
    defparam buf_control_i0_LC_16_16_3.SEQ_MODE=4'b1000;
    defparam buf_control_i0_LC_16_16_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_control_i0_LC_16_16_3 (
            .in0(N__44488),
            .in1(N__44438),
            .in2(_gnd_net_),
            .in3(N__49971),
            .lcout(buf_control_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57952),
            .ce(),
            .sr(_gnd_net_));
    defparam i18970_2_lut_LC_16_16_4.C_ON=1'b0;
    defparam i18970_2_lut_LC_16_16_4.SEQ_MODE=4'b0000;
    defparam i18970_2_lut_LC_16_16_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 i18970_2_lut_LC_16_16_4 (
            .in0(N__52410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48372),
            .lcout(),
            .ltout(n21073_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18852_4_lut_LC_16_16_5.C_ON=1'b0;
    defparam i18852_4_lut_LC_16_16_5.SEQ_MODE=4'b0000;
    defparam i18852_4_lut_LC_16_16_5.LUT_INIT=16'b0010000000000000;
    LogicCell40 i18852_4_lut_LC_16_16_5 (
            .in0(N__49125),
            .in1(N__54736),
            .in2(N__44375),
            .in3(N__48740),
            .lcout(),
            .ltout(n21072_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i2_LC_16_16_6.C_ON=1'b0;
    defparam comm_length_i2_LC_16_16_6.SEQ_MODE=4'b1000;
    defparam comm_length_i2_LC_16_16_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_length_i2_LC_16_16_6 (
            .in0(N__56333),
            .in1(N__51442),
            .in2(N__44372),
            .in3(N__47888),
            .lcout(comm_length_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57952),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19135_4_lut_LC_16_17_3 .C_ON=1'b0;
    defparam \SIG_DDS.i19135_4_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19135_4_lut_LC_16_17_3 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \SIG_DDS.i19135_4_lut_LC_16_17_3  (
            .in0(N__50083),
            .in1(N__44816),
            .in2(N__50362),
            .in3(N__50261),
            .lcout(\SIG_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i12483_3_lut_LC_16_17_4 .C_ON=1'b0;
    defparam \SIG_DDS.i12483_3_lut_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i12483_3_lut_LC_16_17_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \SIG_DDS.i12483_3_lut_LC_16_17_4  (
            .in0(N__50260),
            .in1(N__50349),
            .in2(_gnd_net_),
            .in3(N__50082),
            .lcout(n14900),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_16MHz_I_0_3_lut_LC_16_17_5.C_ON=1'b0;
    defparam clk_16MHz_I_0_3_lut_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam clk_16MHz_I_0_3_lut_LC_16_17_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 clk_16MHz_I_0_3_lut_LC_16_17_5 (
            .in0(N__45098),
            .in1(N__45032),
            .in2(_gnd_net_),
            .in3(N__45016),
            .lcout(DDS_MCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18183_3_lut_LC_16_17_6.C_ON=1'b0;
    defparam i18183_3_lut_LC_16_17_6.SEQ_MODE=4'b0000;
    defparam i18183_3_lut_LC_16_17_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18183_3_lut_LC_16_17_6 (
            .in0(N__44963),
            .in1(N__44927),
            .in2(_gnd_net_),
            .in3(N__48369),
            .lcout(n20797),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19410_LC_16_17_7.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19410_LC_16_17_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19410_LC_16_17_7.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19410_LC_16_17_7 (
            .in0(N__56330),
            .in1(N__44906),
            .in2(N__48409),
            .in3(N__47432),
            .lcout(n22034),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i4_4_lut_LC_16_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.i4_4_lut_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i4_4_lut_LC_16_18_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \SIG_DDS.i4_4_lut_LC_16_18_1  (
            .in0(N__44861),
            .in1(N__44749),
            .in2(N__44846),
            .in3(N__50353),
            .lcout(\SIG_DDS.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i18809_2_lut_LC_16_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.i18809_2_lut_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i18809_2_lut_LC_16_18_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \SIG_DDS.i18809_2_lut_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__44827),
            .in2(_gnd_net_),
            .in3(N__50223),
            .lcout(\SIG_DDS.n21331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i23_4_lut_LC_16_18_4 .C_ON=1'b0;
    defparam \SIG_DDS.i23_4_lut_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i23_4_lut_LC_16_18_4 .LUT_INIT=16'b1100110010011011;
    LogicCell40 \SIG_DDS.i23_4_lut_LC_16_18_4  (
            .in0(N__50354),
            .in1(N__50224),
            .in2(N__44815),
            .in3(N__50084),
            .lcout(\SIG_DDS.n9_adj_1394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i0_LC_16_18_5 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i0_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i0_LC_16_18_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \SIG_DDS.bit_cnt_i0_LC_16_18_5  (
            .in0(N__50086),
            .in1(N__44750),
            .in2(_gnd_net_),
            .in3(N__44764),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57965),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.MOSI_31_LC_16_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.MOSI_31_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.MOSI_31_LC_16_18_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \SIG_DDS.MOSI_31_LC_16_18_7  (
            .in0(N__50085),
            .in1(N__44732),
            .in2(_gnd_net_),
            .in3(N__44692),
            .lcout(DDS_MOSI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57965),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.CS_28_LC_16_19_4 .C_ON=1'b0;
    defparam \SIG_DDS.CS_28_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.CS_28_LC_16_19_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \SIG_DDS.CS_28_LC_16_19_4  (
            .in0(N__50254),
            .in1(N__50360),
            .in2(_gnd_net_),
            .in3(N__50130),
            .lcout(DDS_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57973),
            .ce(N__45260),
            .sr(_gnd_net_));
    defparam i18846_2_lut_LC_17_3_5.C_ON=1'b0;
    defparam i18846_2_lut_LC_17_3_5.SEQ_MODE=4'b0000;
    defparam i18846_2_lut_LC_17_3_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18846_2_lut_LC_17_3_5 (
            .in0(_gnd_net_),
            .in1(N__45245),
            .in2(_gnd_net_),
            .in3(N__56369),
            .lcout(n20984),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_353_Mux_3_i7_4_lut_LC_17_5_0.C_ON=1'b0;
    defparam comm_state_3__I_0_353_Mux_3_i7_4_lut_LC_17_5_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_353_Mux_3_i7_4_lut_LC_17_5_0.LUT_INIT=16'b1110111011110000;
    LogicCell40 comm_state_3__I_0_353_Mux_3_i7_4_lut_LC_17_5_0 (
            .in0(N__45643),
            .in1(N__45799),
            .in2(N__45215),
            .in3(N__52305),
            .lcout(n17738),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11728_2_lut_LC_17_5_1.C_ON=1'b0;
    defparam i11728_2_lut_LC_17_5_1.SEQ_MODE=4'b0000;
    defparam i11728_2_lut_LC_17_5_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 i11728_2_lut_LC_17_5_1 (
            .in0(N__53957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53563),
            .lcout(n14146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i32_4_lut_LC_17_5_2.C_ON=1'b0;
    defparam i32_4_lut_LC_17_5_2.SEQ_MODE=4'b0000;
    defparam i32_4_lut_LC_17_5_2.LUT_INIT=16'b1011100010001000;
    LogicCell40 i32_4_lut_LC_17_5_2 (
            .in0(N__50855),
            .in1(N__53959),
            .in2(N__45206),
            .in3(N__52306),
            .lcout(),
            .ltout(n15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i2_LC_17_5_3.C_ON=1'b0;
    defparam comm_state_i2_LC_17_5_3.SEQ_MODE=4'b1000;
    defparam comm_state_i2_LC_17_5_3.LUT_INIT=16'b1000100011111000;
    LogicCell40 comm_state_i2_LC_17_5_3 (
            .in0(N__49934),
            .in1(N__45134),
            .in2(N__45137),
            .in3(N__53565),
            .lcout(comm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57836),
            .ce(N__50813),
            .sr(N__54836));
    defparam i33_3_lut_LC_17_5_4.C_ON=1'b0;
    defparam i33_3_lut_LC_17_5_4.SEQ_MODE=4'b0000;
    defparam i33_3_lut_LC_17_5_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 i33_3_lut_LC_17_5_4 (
            .in0(N__53564),
            .in1(N__45800),
            .in2(_gnd_net_),
            .in3(N__53958),
            .lcout(n12_adj_1649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_1_i4_3_lut_LC_17_6_0.C_ON=1'b0;
    defparam mux_143_Mux_1_i4_3_lut_LC_17_6_0.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_1_i4_3_lut_LC_17_6_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_143_Mux_1_i4_3_lut_LC_17_6_0 (
            .in0(N__45128),
            .in1(N__45116),
            .in2(_gnd_net_),
            .in3(N__54346),
            .lcout(),
            .ltout(n4_adj_1595_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18193_4_lut_LC_17_6_1.C_ON=1'b0;
    defparam i18193_4_lut_LC_17_6_1.SEQ_MODE=4'b0000;
    defparam i18193_4_lut_LC_17_6_1.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18193_4_lut_LC_17_6_1 (
            .in0(N__54347),
            .in1(N__45289),
            .in2(N__45101),
            .in3(N__50534),
            .lcout(n20807),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_LC_17_6_2.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_LC_17_6_2.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_LC_17_6_2.LUT_INIT=16'b1111100000111000;
    LogicCell40 comm_index_0__bdd_4_lut_LC_17_6_2 (
            .in0(N__45605),
            .in1(N__50535),
            .in2(N__54374),
            .in3(N__45593),
            .lcout(),
            .ltout(n22052_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22052_bdd_4_lut_LC_17_6_3.C_ON=1'b0;
    defparam n22052_bdd_4_lut_LC_17_6_3.SEQ_MODE=4'b0000;
    defparam n22052_bdd_4_lut_LC_17_6_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22052_bdd_4_lut_LC_17_6_3 (
            .in0(N__50536),
            .in1(N__45537),
            .in2(N__45470),
            .in3(N__45453),
            .lcout(),
            .ltout(n22055_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i1_LC_17_6_4.C_ON=1'b0;
    defparam comm_tx_buf_i1_LC_17_6_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i1_LC_17_6_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_tx_buf_i1_LC_17_6_4 (
            .in0(_gnd_net_),
            .in1(N__45413),
            .in2(N__45407),
            .in3(N__50665),
            .lcout(comm_tx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57846),
            .ce(N__46214),
            .sr(N__46132));
    defparam i15005_3_lut_LC_17_6_5.C_ON=1'b0;
    defparam i15005_3_lut_LC_17_6_5.SEQ_MODE=4'b0000;
    defparam i15005_3_lut_LC_17_6_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 i15005_3_lut_LC_17_6_5 (
            .in0(N__50663),
            .in1(N__45404),
            .in2(_gnd_net_),
            .in3(N__45912),
            .lcout(),
            .ltout(n17404_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18337_4_lut_LC_17_6_6.C_ON=1'b0;
    defparam i18337_4_lut_LC_17_6_6.SEQ_MODE=4'b0000;
    defparam i18337_4_lut_LC_17_6_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 i18337_4_lut_LC_17_6_6 (
            .in0(N__45392),
            .in1(N__50537),
            .in2(N__45383),
            .in3(N__50664),
            .lcout(),
            .ltout(n20951_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i5_LC_17_6_7.C_ON=1'b0;
    defparam comm_tx_buf_i5_LC_17_6_7.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i5_LC_17_6_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 comm_tx_buf_i5_LC_17_6_7 (
            .in0(_gnd_net_),
            .in1(N__54351),
            .in2(N__45380),
            .in3(N__45704),
            .lcout(comm_tx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57846),
            .ce(N__46214),
            .sr(N__46132));
    defparam comm_buf_6__i1_LC_17_7_0.C_ON=1'b0;
    defparam comm_buf_6__i1_LC_17_7_0.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i1_LC_17_7_0.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_buf_6__i1_LC_17_7_0 (
            .in0(N__51284),
            .in1(N__45290),
            .in2(N__45376),
            .in3(N__54537),
            .lcout(comm_buf_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57856),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_307_LC_17_7_1.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_307_LC_17_7_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_307_LC_17_7_1.LUT_INIT=16'b0111011111110101;
    LogicCell40 i1_4_lut_4_lut_adj_307_LC_17_7_1 (
            .in0(N__53812),
            .in1(N__53537),
            .in2(N__51782),
            .in3(N__51673),
            .lcout(),
            .ltout(n4_adj_1598_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_84_LC_17_7_2.C_ON=1'b0;
    defparam i1_4_lut_adj_84_LC_17_7_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_84_LC_17_7_2.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_84_LC_17_7_2 (
            .in0(N__51482),
            .in1(N__50834),
            .in2(N__45752),
            .in3(N__45698),
            .lcout(n20573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i235_2_lut_LC_17_7_3.C_ON=1'b0;
    defparam i235_2_lut_LC_17_7_3.SEQ_MODE=4'b0000;
    defparam i235_2_lut_LC_17_7_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 i235_2_lut_LC_17_7_3 (
            .in0(N__51766),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51672),
            .lcout(n1272),
            .ltout(n1272_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_353_Mux_1_i8_3_lut_4_lut_LC_17_7_4.C_ON=1'b0;
    defparam comm_state_3__I_0_353_Mux_1_i8_3_lut_4_lut_LC_17_7_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_353_Mux_1_i8_3_lut_4_lut_LC_17_7_4.LUT_INIT=16'b0001101100010001;
    LogicCell40 comm_state_3__I_0_353_Mux_1_i8_3_lut_4_lut_LC_17_7_4 (
            .in0(N__53538),
            .in1(N__45743),
            .in2(N__45719),
            .in3(N__53813),
            .lcout(n8_adj_1576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22172_bdd_4_lut_LC_17_7_5.C_ON=1'b0;
    defparam n22172_bdd_4_lut_LC_17_7_5.SEQ_MODE=4'b0000;
    defparam n22172_bdd_4_lut_LC_17_7_5.LUT_INIT=16'b1010110110101000;
    LogicCell40 n22172_bdd_4_lut_LC_17_7_5 (
            .in0(N__50414),
            .in1(N__45716),
            .in2(N__50555),
            .in3(N__46355),
            .lcout(n22175),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_299_LC_17_7_6.C_ON=1'b0;
    defparam i2_4_lut_adj_299_LC_17_7_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_299_LC_17_7_6.LUT_INIT=16'b1110111100000000;
    LogicCell40 i2_4_lut_adj_299_LC_17_7_6 (
            .in0(N__50942),
            .in1(N__51476),
            .in2(N__51838),
            .in3(N__45806),
            .lcout(n20551),
            .ltout(n20551_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_17_7_7.C_ON=1'b0;
    defparam i1_4_lut_LC_17_7_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_17_7_7.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_LC_17_7_7 (
            .in0(N__51477),
            .in1(N__45692),
            .in2(N__45683),
            .in3(N__45680),
            .lcout(n20575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_1__bdd_4_lut_LC_17_8_0.C_ON=1'b0;
    defparam comm_state_1__bdd_4_lut_LC_17_8_0.SEQ_MODE=4'b0000;
    defparam comm_state_1__bdd_4_lut_LC_17_8_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_state_1__bdd_4_lut_LC_17_8_0 (
            .in0(N__45659),
            .in1(N__53921),
            .in2(N__45636),
            .in3(N__52376),
            .lcout(n22238),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_353_Mux_1_i2_3_lut_4_lut_LC_17_8_1.C_ON=1'b0;
    defparam comm_state_3__I_0_353_Mux_1_i2_3_lut_4_lut_LC_17_8_1.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_353_Mux_1_i2_3_lut_4_lut_LC_17_8_1.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_state_3__I_0_353_Mux_1_i2_3_lut_4_lut_LC_17_8_1 (
            .in0(N__53466),
            .in1(N__51839),
            .in2(N__54056),
            .in3(N__45821),
            .lcout(),
            .ltout(n2_adj_1575_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22238_bdd_4_lut_LC_17_8_2.C_ON=1'b0;
    defparam n22238_bdd_4_lut_LC_17_8_2.SEQ_MODE=4'b0000;
    defparam n22238_bdd_4_lut_LC_17_8_2.LUT_INIT=16'b1011100110101000;
    LogicCell40 n22238_bdd_4_lut_LC_17_8_2 (
            .in0(N__45614),
            .in1(N__52377),
            .in2(N__45608),
            .in3(N__53467),
            .lcout(),
            .ltout(n22241_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i1_LC_17_8_3.C_ON=1'b0;
    defparam comm_state_i1_LC_17_8_3.SEQ_MODE=4'b1000;
    defparam comm_state_i1_LC_17_8_3.LUT_INIT=16'b0111010000110000;
    LogicCell40 comm_state_i1_LC_17_8_3 (
            .in0(N__49627),
            .in1(N__54722),
            .in2(N__45830),
            .in3(N__45827),
            .lcout(comm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57866),
            .ce(N__50951),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_296_LC_17_8_7.C_ON=1'b0;
    defparam i1_4_lut_adj_296_LC_17_8_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_296_LC_17_8_7.LUT_INIT=16'b1111110100000000;
    LogicCell40 i1_4_lut_adj_296_LC_17_8_7 (
            .in0(N__53465),
            .in1(N__45820),
            .in2(N__51573),
            .in3(N__45812),
            .lcout(n4_adj_1614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_309_LC_17_9_0.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_309_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_309_LC_17_9_0.LUT_INIT=16'b1101111011111111;
    LogicCell40 i1_2_lut_4_lut_adj_309_LC_17_9_0 (
            .in0(N__50493),
            .in1(N__47867),
            .in2(N__47915),
            .in3(N__53774),
            .lcout(n20668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i1_LC_17_9_1.C_ON=1'b0;
    defparam comm_index_i1_LC_17_9_1.SEQ_MODE=4'b1000;
    defparam comm_index_i1_LC_17_9_1.LUT_INIT=16'b1101111100100000;
    LogicCell40 comm_index_i1_LC_17_9_1 (
            .in0(N__51692),
            .in1(N__51842),
            .in2(N__54367),
            .in3(N__50495),
            .lcout(comm_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57876),
            .ce(N__45788),
            .sr(N__45770));
    defparam comm_index_i0_LC_17_9_2.C_ON=1'b0;
    defparam comm_index_i0_LC_17_9_2.SEQ_MODE=4'b1000;
    defparam comm_index_i0_LC_17_9_2.LUT_INIT=16'b1001100111001100;
    LogicCell40 comm_index_i0_LC_17_9_2 (
            .in0(N__51841),
            .in1(N__54320),
            .in2(_gnd_net_),
            .in3(N__51691),
            .lcout(comm_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57876),
            .ce(N__45788),
            .sr(N__45770));
    defparam i1_4_lut_adj_226_LC_17_9_4.C_ON=1'b0;
    defparam i1_4_lut_adj_226_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_226_LC_17_9_4.LUT_INIT=16'b1010111000000000;
    LogicCell40 i1_4_lut_adj_226_LC_17_9_4 (
            .in0(N__54707),
            .in1(N__53350),
            .in2(N__52406),
            .in3(N__51550),
            .lcout(n14753),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i2_LC_17_9_5.C_ON=1'b0;
    defparam comm_index_i2_LC_17_9_5.SEQ_MODE=4'b1000;
    defparam comm_index_i2_LC_17_9_5.LUT_INIT=16'b0111100011110000;
    LogicCell40 comm_index_i2_LC_17_9_5 (
            .in0(N__54319),
            .in1(N__50494),
            .in2(N__50668),
            .in3(N__50854),
            .lcout(comm_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57876),
            .ce(N__45788),
            .sr(N__45770));
    defparam i3_3_lut_LC_17_9_6.C_ON=1'b0;
    defparam i3_3_lut_LC_17_9_6.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_17_9_6.LUT_INIT=16'b0010001000000000;
    LogicCell40 i3_3_lut_LC_17_9_6 (
            .in0(N__52349),
            .in1(N__54318),
            .in2(_gnd_net_),
            .in3(N__53773),
            .lcout(n8_adj_1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_252_LC_17_9_7.C_ON=1'b0;
    defparam i1_4_lut_adj_252_LC_17_9_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_252_LC_17_9_7.LUT_INIT=16'b1010101010000000;
    LogicCell40 i1_4_lut_adj_252_LC_17_9_7 (
            .in0(N__51549),
            .in1(N__52348),
            .in2(N__53351),
            .in3(N__54706),
            .lcout(n11503),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_7_i2_3_lut_LC_17_10_0.C_ON=1'b0;
    defparam mux_143_Mux_7_i2_3_lut_LC_17_10_0.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_7_i2_3_lut_LC_17_10_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_143_Mux_7_i2_3_lut_LC_17_10_0 (
            .in0(N__46253),
            .in1(N__46241),
            .in2(_gnd_net_),
            .in3(N__54290),
            .lcout(),
            .ltout(n2_adj_1581_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i7_LC_17_10_1.C_ON=1'b0;
    defparam comm_tx_buf_i7_LC_17_10_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i7_LC_17_10_1.LUT_INIT=16'b1010101011100100;
    LogicCell40 comm_tx_buf_i7_LC_17_10_1 (
            .in0(N__45923),
            .in1(N__45965),
            .in2(N__46226),
            .in3(N__50632),
            .lcout(comm_tx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57889),
            .ce(N__46198),
            .sr(N__46142));
    defparam i18720_2_lut_LC_17_10_2.C_ON=1'b0;
    defparam i18720_2_lut_LC_17_10_2.SEQ_MODE=4'b0000;
    defparam i18720_2_lut_LC_17_10_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18720_2_lut_LC_17_10_2 (
            .in0(_gnd_net_),
            .in1(N__51265),
            .in2(_gnd_net_),
            .in3(N__54287),
            .lcout(n20966),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_7_i1_3_lut_LC_17_10_3.C_ON=1'b0;
    defparam mux_143_Mux_7_i1_3_lut_LC_17_10_3.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_7_i1_3_lut_LC_17_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_143_Mux_7_i1_3_lut_LC_17_10_3 (
            .in0(N__54289),
            .in1(N__47630),
            .in2(_gnd_net_),
            .in3(N__46041),
            .lcout(n1_adj_1580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_143_Mux_7_i4_3_lut_LC_17_10_4.C_ON=1'b0;
    defparam mux_143_Mux_7_i4_3_lut_LC_17_10_4.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_7_i4_3_lut_LC_17_10_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_143_Mux_7_i4_3_lut_LC_17_10_4 (
            .in0(N__45959),
            .in1(N__45944),
            .in2(_gnd_net_),
            .in3(N__54288),
            .lcout(),
            .ltout(n4_adj_1582_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19361_LC_17_10_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19361_LC_17_10_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19361_LC_17_10_5.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_index_1__bdd_4_lut_19361_LC_17_10_5 (
            .in0(N__45932),
            .in1(N__50506),
            .in2(N__45926),
            .in3(N__50631),
            .lcout(n21968),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19194_4_lut_3_lut_LC_17_10_6 .C_ON=1'b0;
    defparam \comm_spi.i19194_4_lut_3_lut_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19194_4_lut_3_lut_LC_17_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19194_4_lut_3_lut_LC_17_10_6  (
            .in0(N__55450),
            .in1(N__56505),
            .in2(_gnd_net_),
            .in3(N__56807),
            .lcout(\comm_spi.n14619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15244_2_lut_3_lut_LC_17_11_0.C_ON=1'b0;
    defparam i15244_2_lut_3_lut_LC_17_11_0.SEQ_MODE=4'b0000;
    defparam i15244_2_lut_3_lut_LC_17_11_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15244_2_lut_3_lut_LC_17_11_0 (
            .in0(N__53951),
            .in1(N__45886),
            .in2(_gnd_net_),
            .in3(N__52365),
            .lcout(n14_adj_1578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19029_2_lut_LC_17_11_1.C_ON=1'b0;
    defparam i19029_2_lut_LC_17_11_1.SEQ_MODE=4'b0000;
    defparam i19029_2_lut_LC_17_11_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19029_2_lut_LC_17_11_1 (
            .in0(_gnd_net_),
            .in1(N__45854),
            .in2(_gnd_net_),
            .in3(N__56357),
            .lcout(n21270),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_238_LC_17_11_2.C_ON=1'b0;
    defparam i1_4_lut_adj_238_LC_17_11_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_238_LC_17_11_2.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_238_LC_17_11_2 (
            .in0(N__46613),
            .in1(N__54824),
            .in2(N__49701),
            .in3(N__46586),
            .lcout(n12467),
            .ltout(n12467_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i0_LC_17_11_3.C_ON=1'b0;
    defparam req_data_cnt_i0_LC_17_11_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i0_LC_17_11_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 req_data_cnt_i0_LC_17_11_3 (
            .in0(_gnd_net_),
            .in1(N__46461),
            .in2(N__46550),
            .in3(N__46543),
            .lcout(req_data_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57901),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_191_LC_17_11_4.C_ON=1'b0;
    defparam i1_4_lut_adj_191_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_191_LC_17_11_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_191_LC_17_11_4 (
            .in0(N__46523),
            .in1(N__46496),
            .in2(N__46465),
            .in3(N__46323),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21956_bdd_4_lut_LC_17_11_5.C_ON=1'b0;
    defparam n21956_bdd_4_lut_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam n21956_bdd_4_lut_LC_17_11_5.LUT_INIT=16'b1010101011100100;
    LogicCell40 n21956_bdd_4_lut_LC_17_11_5 (
            .in0(N__46880),
            .in1(N__46436),
            .in2(N__51873),
            .in3(N__49126),
            .lcout(n21959),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_102_LC_17_11_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_102_LC_17_11_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_102_LC_17_11_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i1_2_lut_3_lut_adj_102_LC_17_11_6 (
            .in0(N__53950),
            .in1(N__46367),
            .in2(_gnd_net_),
            .in3(N__52364),
            .lcout(n14_adj_1577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i6_LC_17_11_7.C_ON=1'b0;
    defparam req_data_cnt_i6_LC_17_11_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i6_LC_17_11_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i6_LC_17_11_7 (
            .in0(N__46324),
            .in1(N__52174),
            .in2(_gnd_net_),
            .in3(N__47350),
            .lcout(req_data_cnt_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57901),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_LC_17_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_LC_17_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_LC_17_12_0.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_1__bdd_4_lut_LC_17_12_0 (
            .in0(N__48418),
            .in1(N__49102),
            .in2(N__55700),
            .in3(N__46823),
            .lcout(),
            .ltout(n22208_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22208_bdd_4_lut_LC_17_12_1.C_ON=1'b0;
    defparam n22208_bdd_4_lut_LC_17_12_1.SEQ_MODE=4'b0000;
    defparam n22208_bdd_4_lut_LC_17_12_1.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22208_bdd_4_lut_LC_17_12_1 (
            .in0(N__49103),
            .in1(N__46309),
            .in2(N__46292),
            .in3(N__46289),
            .lcout(),
            .ltout(n22211_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1546664_i1_3_lut_LC_17_12_2.C_ON=1'b0;
    defparam i1546664_i1_3_lut_LC_17_12_2.SEQ_MODE=4'b0000;
    defparam i1546664_i1_3_lut_LC_17_12_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1546664_i1_3_lut_LC_17_12_2 (
            .in0(_gnd_net_),
            .in1(N__46262),
            .in2(N__47255),
            .in3(N__48676),
            .lcout(),
            .ltout(n30_adj_1518_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i2_LC_17_12_3.C_ON=1'b0;
    defparam comm_buf_1__i2_LC_17_12_3.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i2_LC_17_12_3.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_1__i2_LC_17_12_3 (
            .in0(N__54027),
            .in1(N__47246),
            .in2(N__47153),
            .in3(_gnd_net_),
            .lcout(comm_buf_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57918),
            .ce(N__47075),
            .sr(N__46996));
    defparam comm_cmd_1__bdd_4_lut_19375_LC_17_12_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19375_LC_17_12_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19375_LC_17_12_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19375_LC_17_12_4 (
            .in0(N__46916),
            .in1(N__48414),
            .in2(N__46901),
            .in3(N__49101),
            .lcout(n21956),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_2_i26_3_lut_LC_17_12_6.C_ON=1'b0;
    defparam mux_135_Mux_2_i26_3_lut_LC_17_12_6.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_2_i26_3_lut_LC_17_12_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_2_i26_3_lut_LC_17_12_6 (
            .in0(N__46874),
            .in1(N__56362),
            .in2(_gnd_net_),
            .in3(N__46850),
            .lcout(n26_adj_1517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i1_LC_17_13_1.C_ON=1'b0;
    defparam req_data_cnt_i1_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i1_LC_17_13_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i1_LC_17_13_1 (
            .in0(N__47376),
            .in1(N__46817),
            .in2(_gnd_net_),
            .in3(N__46690),
            .lcout(req_data_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57929),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i15_LC_17_13_2.C_ON=1'b0;
    defparam req_data_cnt_i15_LC_17_13_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i15_LC_17_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i15_LC_17_13_2 (
            .in0(N__46796),
            .in1(N__47375),
            .in2(_gnd_net_),
            .in3(N__47506),
            .lcout(req_data_cnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57929),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_188_LC_17_13_3.C_ON=1'b0;
    defparam i2_4_lut_adj_188_LC_17_13_3.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_188_LC_17_13_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_188_LC_17_13_3 (
            .in0(N__46772),
            .in1(N__46745),
            .in2(N__46723),
            .in3(N__46689),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_5_i19_3_lut_LC_17_13_4.C_ON=1'b0;
    defparam mux_135_Mux_5_i19_3_lut_LC_17_13_4.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_5_i19_3_lut_LC_17_13_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_135_Mux_5_i19_3_lut_LC_17_13_4 (
            .in0(N__46670),
            .in1(N__46642),
            .in2(_gnd_net_),
            .in3(N__56338),
            .lcout(n19_adj_1497),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i3_LC_17_13_5.C_ON=1'b0;
    defparam req_data_cnt_i3_LC_17_13_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i3_LC_17_13_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i3_LC_17_13_5 (
            .in0(N__47377),
            .in1(N__47842),
            .in2(_gnd_net_),
            .in3(N__47701),
            .lcout(req_data_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57929),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_134_Mux_7_i23_3_lut_LC_17_13_6.C_ON=1'b0;
    defparam mux_134_Mux_7_i23_3_lut_LC_17_13_6.SEQ_MODE=4'b0000;
    defparam mux_134_Mux_7_i23_3_lut_LC_17_13_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_134_Mux_7_i23_3_lut_LC_17_13_6 (
            .in0(N__51233),
            .in1(N__56337),
            .in2(_gnd_net_),
            .in3(N__47794),
            .lcout(n23_adj_1527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_185_LC_17_13_7.C_ON=1'b0;
    defparam i4_4_lut_adj_185_LC_17_13_7.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_185_LC_17_13_7.LUT_INIT=16'b0111101111011110;
    LogicCell40 i4_4_lut_adj_185_LC_17_13_7 (
            .in0(N__47752),
            .in1(N__47732),
            .in2(N__47284),
            .in3(N__47700),
            .lcout(n20_adj_1596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15258_2_lut_3_lut_LC_17_14_1.C_ON=1'b0;
    defparam i15258_2_lut_3_lut_LC_17_14_1.SEQ_MODE=4'b0000;
    defparam i15258_2_lut_3_lut_LC_17_14_1.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15258_2_lut_3_lut_LC_17_14_1 (
            .in0(N__47656),
            .in1(N__54076),
            .in2(_gnd_net_),
            .in3(N__52366),
            .lcout(n14_adj_1546),
            .ltout(n14_adj_1546_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i7_LC_17_14_2.C_ON=1'b0;
    defparam req_data_cnt_i7_LC_17_14_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i7_LC_17_14_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 req_data_cnt_i7_LC_17_14_2 (
            .in0(N__47380),
            .in1(_gnd_net_),
            .in2(N__47594),
            .in3(N__49153),
            .lcout(req_data_cnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57942),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i13_LC_17_14_3.C_ON=1'b0;
    defparam req_data_cnt_i13_LC_17_14_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i13_LC_17_14_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i13_LC_17_14_3 (
            .in0(N__47575),
            .in1(N__47378),
            .in2(_gnd_net_),
            .in3(N__47551),
            .lcout(req_data_cnt_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57942),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_180_LC_17_14_4.C_ON=1'b0;
    defparam i8_4_lut_adj_180_LC_17_14_4.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_180_LC_17_14_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i8_4_lut_adj_180_LC_17_14_4 (
            .in0(N__47531),
            .in1(N__47502),
            .in2(N__47486),
            .in3(N__47427),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i9_LC_17_14_5.C_ON=1'b0;
    defparam req_data_cnt_i9_LC_17_14_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i9_LC_17_14_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i9_LC_17_14_5 (
            .in0(N__47428),
            .in1(N__47461),
            .in2(_gnd_net_),
            .in3(N__47381),
            .lcout(req_data_cnt_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57942),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i5_LC_17_14_6.C_ON=1'b0;
    defparam req_data_cnt_i5_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i5_LC_17_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i5_LC_17_14_6 (
            .in0(N__47379),
            .in1(N__47326),
            .in2(_gnd_net_),
            .in3(N__47283),
            .lcout(req_data_cnt_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57942),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i4_LC_17_14_7.C_ON=1'b0;
    defparam acadc_skipCount_i4_LC_17_14_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i4_LC_17_14_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i4_LC_17_14_7 (
            .in0(N__49834),
            .in1(N__49372),
            .in2(N__51187),
            .in3(N__49275),
            .lcout(acadc_skipCount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57942),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_135_Mux_7_i26_3_lut_LC_17_15_0.C_ON=1'b0;
    defparam mux_135_Mux_7_i26_3_lut_LC_17_15_0.SEQ_MODE=4'b0000;
    defparam mux_135_Mux_7_i26_3_lut_LC_17_15_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_135_Mux_7_i26_3_lut_LC_17_15_0 (
            .in0(N__49253),
            .in1(N__56371),
            .in2(_gnd_net_),
            .in3(N__49229),
            .lcout(),
            .ltout(n26_adj_1500_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18196_4_lut_LC_17_15_1.C_ON=1'b0;
    defparam i18196_4_lut_LC_17_15_1.SEQ_MODE=4'b0000;
    defparam i18196_4_lut_LC_17_15_1.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18196_4_lut_LC_17_15_1 (
            .in0(N__56372),
            .in1(N__49205),
            .in2(N__49193),
            .in3(N__48415),
            .lcout(),
            .ltout(n20810_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19454_LC_17_15_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19454_LC_17_15_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19454_LC_17_15_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19454_LC_17_15_2 (
            .in0(N__49133),
            .in1(N__48730),
            .in2(N__49190),
            .in3(N__49121),
            .lcout(n22058),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18195_3_lut_LC_17_15_3.C_ON=1'b0;
    defparam i18195_3_lut_LC_17_15_3.SEQ_MODE=4'b0000;
    defparam i18195_3_lut_LC_17_15_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18195_3_lut_LC_17_15_3 (
            .in0(N__48410),
            .in1(N__49180),
            .in2(_gnd_net_),
            .in3(N__49152),
            .lcout(n20809),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i0_LC_17_15_4.C_ON=1'b0;
    defparam comm_length_i0_LC_17_15_4.SEQ_MODE=4'b1000;
    defparam comm_length_i0_LC_17_15_4.LUT_INIT=16'b0000011110011010;
    LogicCell40 comm_length_i0_LC_17_15_4 (
            .in0(N__48416),
            .in1(N__56373),
            .in2(N__48728),
            .in3(N__49123),
            .lcout(comm_length_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57953),
            .ce(N__51443),
            .sr(N__50405));
    defparam comm_length_i1_LC_17_15_5.C_ON=1'b0;
    defparam comm_length_i1_LC_17_15_5.SEQ_MODE=4'b1000;
    defparam comm_length_i1_LC_17_15_5.LUT_INIT=16'b1011110011111011;
    LogicCell40 comm_length_i1_LC_17_15_5 (
            .in0(N__49122),
            .in1(N__48677),
            .in2(N__56378),
            .in3(N__48417),
            .lcout(comm_length_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57953),
            .ce(N__51443),
            .sr(N__50405));
    defparam i1_4_lut_adj_244_LC_17_15_6.C_ON=1'b0;
    defparam i1_4_lut_adj_244_LC_17_15_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_244_LC_17_15_6.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_244_LC_17_15_6 (
            .in0(N__47887),
            .in1(N__54308),
            .in2(N__47876),
            .in3(N__50684),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_17_16_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_17_16_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_94_2_lut_LC_17_16_3  (
            .in0(N__56751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55237),
            .lcout(\comm_spi.data_tx_7__N_769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12253_3_lut_LC_17_16_4.C_ON=1'b0;
    defparam i12253_3_lut_LC_17_16_4.SEQ_MODE=4'b0000;
    defparam i12253_3_lut_LC_17_16_4.LUT_INIT=16'b1010101000100010;
    LogicCell40 i12253_3_lut_LC_17_16_4 (
            .in0(N__51435),
            .in1(N__52367),
            .in2(_gnd_net_),
            .in3(N__54912),
            .lcout(n14671),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i1_LC_17_17_7 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i1_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i1_LC_17_17_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.dds_state_i1_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(N__50262),
            .in2(_gnd_net_),
            .in3(N__50359),
            .lcout(dds_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57966),
            .ce(N__50381),
            .sr(N__50186));
    defparam \SIG_DDS.dds_state_i0_LC_17_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i0_LC_17_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i0_LC_17_18_2 .LUT_INIT=16'b1010000000110011;
    LogicCell40 \SIG_DDS.dds_state_i0_LC_17_18_2  (
            .in0(N__50396),
            .in1(N__50358),
            .in2(N__50390),
            .in3(N__50098),
            .lcout(dds_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57974),
            .ce(N__50380),
            .sr(_gnd_net_));
    defparam \SIG_DDS.SCLK_27_LC_17_19_1 .C_ON=1'b0;
    defparam \SIG_DDS.SCLK_27_LC_17_19_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.SCLK_27_LC_17_19_1 .LUT_INIT=16'b0011001010110001;
    LogicCell40 \SIG_DDS.SCLK_27_LC_17_19_1  (
            .in0(N__50361),
            .in1(N__50250),
            .in2(N__50026),
            .in3(N__50131),
            .lcout(DDS_SCK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57976),
            .ce(),
            .sr(_gnd_net_));
    defparam i15030_2_lut_2_lut_LC_17_19_7.C_ON=1'b0;
    defparam i15030_2_lut_2_lut_LC_17_19_7.SEQ_MODE=4'b0000;
    defparam i15030_2_lut_2_lut_LC_17_19_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 i15030_2_lut_2_lut_LC_17_19_7 (
            .in0(N__50009),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49978),
            .lcout(CONT_SD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15087_2_lut_LC_18_5_1.C_ON=1'b0;
    defparam i15087_2_lut_LC_18_5_1.SEQ_MODE=4'b0000;
    defparam i15087_2_lut_LC_18_5_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 i15087_2_lut_LC_18_5_1 (
            .in0(_gnd_net_),
            .in1(N__54655),
            .in2(_gnd_net_),
            .in3(N__53562),
            .lcout(n17485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_224_LC_18_5_3.C_ON=1'b0;
    defparam i1_2_lut_adj_224_LC_18_5_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_224_LC_18_5_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 i1_2_lut_adj_224_LC_18_5_3 (
            .in0(N__51741),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52304),
            .lcout(n20608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i46_2_lut_LC_18_5_4.C_ON=1'b0;
    defparam i46_2_lut_LC_18_5_4.SEQ_MODE=4'b0000;
    defparam i46_2_lut_LC_18_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 i46_2_lut_LC_18_5_4 (
            .in0(_gnd_net_),
            .in1(N__51745),
            .in2(_gnd_net_),
            .in3(N__53955),
            .lcout(n23_adj_1501),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_18_5_5.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_18_5_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_18_5_5.LUT_INIT=16'b0010011000000000;
    LogicCell40 i1_4_lut_4_lut_LC_18_5_5 (
            .in0(N__53956),
            .in1(N__52302),
            .in2(N__51762),
            .in3(N__51690),
            .lcout(),
            .ltout(n21_adj_1600_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19152_4_lut_LC_18_5_6.C_ON=1'b0;
    defparam i19152_4_lut_LC_18_5_6.SEQ_MODE=4'b0000;
    defparam i19152_4_lut_LC_18_5_6.LUT_INIT=16'b0000101111111111;
    LogicCell40 i19152_4_lut_LC_18_5_6 (
            .in0(N__52303),
            .in1(N__50828),
            .in2(N__50822),
            .in3(N__50819),
            .lcout(n18_adj_1633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12212_12213_set_LC_18_6_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12212_12213_set_LC_18_6_6 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_rx_i0_12212_12213_set_LC_18_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_rx_i0_12212_12213_set_LC_18_6_6  (
            .in0(N__53327),
            .in1(N__53300),
            .in2(_gnd_net_),
            .in3(N__53279),
            .lcout(\comm_spi.n14630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57062),
            .ce(),
            .sr(N__52526));
    defparam \comm_spi.i12200_3_lut_LC_18_7_0 .C_ON=1'b0;
    defparam \comm_spi.i12200_3_lut_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12200_3_lut_LC_18_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i12200_3_lut_LC_18_7_0  (
            .in0(N__53295),
            .in1(N__53277),
            .in2(_gnd_net_),
            .in3(N__53324),
            .lcout(\comm_spi.imosi ),
            .ltout(\comm_spi.imosi_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19204_4_lut_3_lut_LC_18_7_1 .C_ON=1'b0;
    defparam \comm_spi.i19204_4_lut_3_lut_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19204_4_lut_3_lut_LC_18_7_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \comm_spi.i19204_4_lut_3_lut_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(N__50801),
            .in2(N__50804),
            .in3(N__56777),
            .lcout(\comm_spi.n22667 ),
            .ltout(\comm_spi.n22667_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12214_3_lut_LC_18_7_2 .C_ON=1'b0;
    defparam \comm_spi.i12214_3_lut_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12214_3_lut_LC_18_7_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.i12214_3_lut_LC_18_7_2  (
            .in0(_gnd_net_),
            .in1(N__50795),
            .in2(N__50786),
            .in3(N__53306),
            .lcout(comm_rx_buf_0),
            .ltout(comm_rx_buf_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i0_LC_18_7_3.C_ON=1'b0;
    defparam comm_buf_6__i0_LC_18_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i0_LC_18_7_3.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i0_LC_18_7_3 (
            .in0(N__50701),
            .in1(N__54723),
            .in2(N__50705),
            .in3(N__51298),
            .lcout(comm_buf_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57867),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_2__bdd_4_lut_LC_18_7_5.C_ON=1'b0;
    defparam comm_index_2__bdd_4_lut_LC_18_7_5.SEQ_MODE=4'b0000;
    defparam comm_index_2__bdd_4_lut_LC_18_7_5.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_2__bdd_4_lut_LC_18_7_5 (
            .in0(N__50662),
            .in1(N__50567),
            .in2(N__50969),
            .in3(N__50548),
            .lcout(n22172),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i5_LC_18_7_6.C_ON=1'b0;
    defparam comm_buf_6__i5_LC_18_7_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i5_LC_18_7_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_buf_6__i5_LC_18_7_6 (
            .in0(N__51299),
            .in1(N__51042),
            .in2(N__54837),
            .in3(N__50968),
            .lcout(comm_buf_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57867),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19189_4_lut_3_lut_LC_18_7_7 .C_ON=1'b0;
    defparam \comm_spi.i19189_4_lut_3_lut_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19189_4_lut_3_lut_LC_18_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19189_4_lut_3_lut_LC_18_7_7  (
            .in0(N__53325),
            .in1(N__58135),
            .in2(_gnd_net_),
            .in3(N__56776),
            .lcout(\comm_spi.n22670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_290_LC_18_8_0.C_ON=1'b0;
    defparam i1_2_lut_adj_290_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_290_LC_18_8_0.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_290_LC_18_8_0 (
            .in0(N__54708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52368),
            .lcout(n12235),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_130_LC_18_8_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_130_LC_18_8_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_130_LC_18_8_1.LUT_INIT=16'b1110111000000000;
    LogicCell40 i1_2_lut_3_lut_adj_130_LC_18_8_1 (
            .in0(N__53787),
            .in1(N__52369),
            .in2(_gnd_net_),
            .in3(N__54709),
            .lcout(n19904),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i469_2_lut_LC_18_8_3.C_ON=1'b0;
    defparam i469_2_lut_LC_18_8_3.SEQ_MODE=4'b0000;
    defparam i469_2_lut_LC_18_8_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 i469_2_lut_LC_18_8_3 (
            .in0(N__51747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51688),
            .lcout(n2369),
            .ltout(n2369_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19055_4_lut_LC_18_8_4.C_ON=1'b0;
    defparam i19055_4_lut_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam i19055_4_lut_LC_18_8_4.LUT_INIT=16'b0011000100100000;
    LogicCell40 i19055_4_lut_LC_18_8_4 (
            .in0(N__52370),
            .in1(N__53788),
            .in2(N__50957),
            .in3(N__51746),
            .lcout(),
            .ltout(n21130_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19149_4_lut_LC_18_8_5.C_ON=1'b0;
    defparam i19149_4_lut_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam i19149_4_lut_LC_18_8_5.LUT_INIT=16'b1111111100011011;
    LogicCell40 i19149_4_lut_LC_18_8_5 (
            .in0(N__53554),
            .in1(N__51611),
            .in2(N__50954),
            .in3(N__54710),
            .lcout(n14_adj_1506),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15091_2_lut_LC_18_8_6.C_ON=1'b0;
    defparam i15091_2_lut_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam i15091_2_lut_LC_18_8_6.LUT_INIT=16'b1100110011111111;
    LogicCell40 i15091_2_lut_LC_18_8_6 (
            .in0(_gnd_net_),
            .in1(N__53786),
            .in2(_gnd_net_),
            .in3(N__53553),
            .lcout(n3),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_18_8_7.C_ON=1'b0;
    defparam i2_3_lut_LC_18_8_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_18_8_7.LUT_INIT=16'b1111110011111111;
    LogicCell40 i2_3_lut_LC_18_8_7 (
            .in0(_gnd_net_),
            .in1(N__50932),
            .in2(N__50858),
            .in3(N__50850),
            .lcout(n19655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18885_2_lut_3_lut_LC_18_9_0.C_ON=1'b0;
    defparam i18885_2_lut_3_lut_LC_18_9_0.SEQ_MODE=4'b0000;
    defparam i18885_2_lut_3_lut_LC_18_9_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 i18885_2_lut_3_lut_LC_18_9_0 (
            .in0(N__51840),
            .in1(N__51689),
            .in2(_gnd_net_),
            .in3(N__53804),
            .lcout(n21129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18127_2_lut_LC_18_9_2.C_ON=1'b0;
    defparam i18127_2_lut_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam i18127_2_lut_LC_18_9_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 i18127_2_lut_LC_18_9_2 (
            .in0(_gnd_net_),
            .in1(N__53805),
            .in2(_gnd_net_),
            .in3(N__53505),
            .lcout(n20740),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_178_LC_18_9_4.C_ON=1'b0;
    defparam i1_2_lut_adj_178_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_178_LC_18_9_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_178_LC_18_9_4 (
            .in0(_gnd_net_),
            .in1(N__52420),
            .in2(_gnd_net_),
            .in3(N__53506),
            .lcout(),
            .ltout(n11363_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_229_LC_18_9_5.C_ON=1'b0;
    defparam i1_4_lut_adj_229_LC_18_9_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_229_LC_18_9_5.LUT_INIT=16'b1100110000001000;
    LogicCell40 i1_4_lut_adj_229_LC_18_9_5 (
            .in0(N__53806),
            .in1(N__51552),
            .in2(N__51593),
            .in3(N__54717),
            .lcout(n11935),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_88_LC_18_9_6.C_ON=1'b0;
    defparam i1_4_lut_adj_88_LC_18_9_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_88_LC_18_9_6.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_88_LC_18_9_6 (
            .in0(N__53346),
            .in1(N__51551),
            .in2(N__51481),
            .in3(N__51455),
            .lcout(n11876),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i7_LC_18_9_7.C_ON=1'b0;
    defparam comm_buf_6__i7_LC_18_9_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i7_LC_18_9_7.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i7_LC_18_9_7 (
            .in0(N__51266),
            .in1(N__54718),
            .in2(N__51407),
            .in3(N__51311),
            .lcout(comm_buf_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57890),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i7_LC_18_10_2.C_ON=1'b0;
    defparam buf_control_i7_LC_18_10_2.SEQ_MODE=4'b1000;
    defparam buf_control_i7_LC_18_10_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 buf_control_i7_LC_18_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51254),
            .lcout(buf_control_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57902),
            .ce(N__51224),
            .sr(N__51208));
    defparam i15260_2_lut_3_lut_LC_18_11_0.C_ON=1'b0;
    defparam i15260_2_lut_3_lut_LC_18_11_0.SEQ_MODE=4'b0000;
    defparam i15260_2_lut_3_lut_LC_18_11_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15260_2_lut_3_lut_LC_18_11_0 (
            .in0(N__51181),
            .in1(N__53964),
            .in2(_gnd_net_),
            .in3(N__52412),
            .lcout(n14_adj_1548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_18_11_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_18_11_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i20_LC_18_11_1  (
            .in0(N__53012),
            .in1(N__53254),
            .in2(N__51076),
            .in3(N__52088),
            .lcout(cmd_rdadctmp_20_adj_1430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57919),
            .ce(),
            .sr(_gnd_net_));
    defparam i15259_2_lut_3_lut_LC_18_11_2.C_ON=1'b0;
    defparam i15259_2_lut_3_lut_LC_18_11_2.SEQ_MODE=4'b0000;
    defparam i15259_2_lut_3_lut_LC_18_11_2.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15259_2_lut_3_lut_LC_18_11_2 (
            .in0(N__52493),
            .in1(N__53963),
            .in2(_gnd_net_),
            .in3(N__52411),
            .lcout(n14_adj_1547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19184_4_lut_3_lut_LC_18_11_6 .C_ON=1'b0;
    defparam \comm_spi.i19184_4_lut_3_lut_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19184_4_lut_3_lut_LC_18_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i19184_4_lut_3_lut_LC_18_11_6  (
            .in0(N__56809),
            .in1(N__58055),
            .in2(_gnd_net_),
            .in3(N__56425),
            .lcout(\comm_spi.n22664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_18_11_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_18_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_92_2_lut_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__56506),
            .in2(_gnd_net_),
            .in3(N__56808),
            .lcout(\comm_spi.data_tx_7__N_767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i8_LC_18_12_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i8_LC_18_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i8_LC_18_12_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i8_LC_18_12_0  (
            .in0(N__53002),
            .in1(N__53179),
            .in2(N__52121),
            .in3(N__52143),
            .lcout(buf_adcdata_iac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57930),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19199_4_lut_3_lut_LC_18_12_1 .C_ON=1'b0;
    defparam \comm_spi.i19199_4_lut_3_lut_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19199_4_lut_3_lut_LC_18_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i19199_4_lut_3_lut_LC_18_12_1  (
            .in0(N__56816),
            .in1(N__55020),
            .in2(_gnd_net_),
            .in3(N__55068),
            .lcout(\comm_spi.n22685 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_18_12_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_18_12_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i17_LC_18_12_2  (
            .in0(N__53003),
            .in1(N__52626),
            .in2(N__52120),
            .in3(N__52086),
            .lcout(cmd_rdadctmp_17_adj_1433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57930),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_18_12_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_18_12_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i18_LC_18_12_3  (
            .in0(N__52085),
            .in1(N__51885),
            .in2(N__52633),
            .in3(N__53007),
            .lcout(cmd_rdadctmp_18_adj_1432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57930),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_18_12_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_18_12_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i19_LC_18_12_4  (
            .in0(N__53004),
            .in1(N__53250),
            .in2(N__51890),
            .in3(N__52087),
            .lcout(cmd_rdadctmp_19_adj_1431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57930),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i10_LC_18_12_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i10_LC_18_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i10_LC_18_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i10_LC_18_12_5  (
            .in0(N__53177),
            .in1(N__53005),
            .in2(N__51874),
            .in3(N__51889),
            .lcout(buf_adcdata_iac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57930),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19219_4_lut_3_lut_LC_18_12_6 .C_ON=1'b0;
    defparam \comm_spi.i19219_4_lut_3_lut_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19219_4_lut_3_lut_LC_18_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19219_4_lut_3_lut_LC_18_12_6  (
            .in0(N__58224),
            .in1(N__55272),
            .in2(_gnd_net_),
            .in3(N__56817),
            .lcout(\comm_spi.n22676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i11_LC_18_12_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i11_LC_18_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i11_LC_18_12_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i11_LC_18_12_7  (
            .in0(N__53178),
            .in1(N__53006),
            .in2(N__53255),
            .in3(N__53229),
            .lcout(buf_adcdata_iac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57930),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i9_LC_18_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i9_LC_18_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i9_LC_18_13_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i9_LC_18_13_0  (
            .in0(N__53176),
            .in1(N__53011),
            .in2(N__52634),
            .in3(N__52602),
            .lcout(buf_adcdata_iac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57943),
            .ce(),
            .sr(_gnd_net_));
    defparam i18953_2_lut_LC_18_13_2.C_ON=1'b0;
    defparam i18953_2_lut_LC_18_13_2.SEQ_MODE=4'b0000;
    defparam i18953_2_lut_LC_18_13_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18953_2_lut_LC_18_13_2 (
            .in0(_gnd_net_),
            .in1(N__52583),
            .in2(_gnd_net_),
            .in3(N__56317),
            .lcout(n21230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_18_13_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_18_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_106_2_lut_LC_18_13_3  (
            .in0(N__55027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56775),
            .lcout(\comm_spi.data_tx_7__N_793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19021_2_lut_LC_18_14_3.C_ON=1'b0;
    defparam i19021_2_lut_LC_18_14_3.SEQ_MODE=4'b0000;
    defparam i19021_2_lut_LC_18_14_3.LUT_INIT=16'b1110111011101110;
    LogicCell40 i19021_2_lut_LC_18_14_3 (
            .in0(N__56313),
            .in1(N__52553),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n21297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_18_14_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_18_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_86_2_lut_LC_18_14_5  (
            .in0(N__56760),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55127),
            .lcout(\comm_spi.DOUT_7__N_747 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19209_4_lut_3_lut_LC_18_15_0 .C_ON=1'b0;
    defparam \comm_spi.i19209_4_lut_3_lut_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19209_4_lut_3_lut_LC_18_15_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19209_4_lut_3_lut_LC_18_15_0  (
            .in0(N__55386),
            .in1(N__55160),
            .in2(_gnd_net_),
            .in3(N__56745),
            .lcout(\comm_spi.n22682 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_18_15_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_18_15_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_104_2_lut_LC_18_15_4  (
            .in0(N__55318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56743),
            .lcout(\comm_spi.data_tx_7__N_787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_18_15_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_18_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_95_2_lut_LC_18_15_6  (
            .in0(N__55279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56744),
            .lcout(\comm_spi.data_tx_7__N_770 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_18_15_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_18_15_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_101_2_lut_LC_18_15_7  (
            .in0(N__56742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55510),
            .lcout(\comm_spi.data_tx_7__N_778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_clear_311_LC_18_16_0.C_ON=1'b0;
    defparam comm_clear_311_LC_18_16_0.SEQ_MODE=4'b1000;
    defparam comm_clear_311_LC_18_16_0.LUT_INIT=16'b0111011101010101;
    LogicCell40 comm_clear_311_LC_18_16_0 (
            .in0(N__54170),
            .in1(N__54913),
            .in2(_gnd_net_),
            .in3(N__53582),
            .lcout(comm_clear),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57967),
            .ce(N__54431),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i4_12228_12229_set_LC_18_17_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12228_12229_set_LC_18_17_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i4_12228_12229_set_LC_18_17_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i4_12228_12229_set_LC_18_17_0  (
            .in0(N__55187),
            .in1(N__55220),
            .in2(_gnd_net_),
            .in3(N__55201),
            .lcout(\comm_spi.n14646 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57049),
            .ce(),
            .sr(N__54416));
    defparam mux_143_Mux_6_i4_3_lut_LC_19_6_2.C_ON=1'b0;
    defparam mux_143_Mux_6_i4_3_lut_LC_19_6_2.SEQ_MODE=4'b0000;
    defparam mux_143_Mux_6_i4_3_lut_LC_19_6_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_143_Mux_6_i4_3_lut_LC_19_6_2 (
            .in0(N__54407),
            .in1(N__54395),
            .in2(_gnd_net_),
            .in3(N__54368),
            .lcout(n4_adj_1585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6849_2_lut_LC_19_6_7.C_ON=1'b0;
    defparam i6849_2_lut_LC_19_6_7.SEQ_MODE=4'b0000;
    defparam i6849_2_lut_LC_19_6_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 i6849_2_lut_LC_19_6_7 (
            .in0(_gnd_net_),
            .in1(N__54028),
            .in2(_gnd_net_),
            .in3(N__53548),
            .lcout(n9270),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12212_12213_reset_LC_19_7_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12212_12213_reset_LC_19_7_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i0_12212_12213_reset_LC_19_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_rx_i0_12212_12213_reset_LC_19_7_2  (
            .in0(N__53326),
            .in1(N__53296),
            .in2(_gnd_net_),
            .in3(N__53278),
            .lcout(\comm_spi.n14631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57058),
            .ce(),
            .sr(N__55106));
    defparam \comm_spi.imosi_44_12198_12199_set_LC_19_8_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12198_12199_set_LC_19_8_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imosi_44_12198_12199_set_LC_19_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.imosi_44_12198_12199_set_LC_19_8_0  (
            .in0(N__58152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57891),
            .ce(),
            .sr(N__55094));
    defparam \comm_spi.imosi_44_12198_12199_reset_LC_19_9_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12198_12199_reset_LC_19_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imosi_44_12198_12199_reset_LC_19_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_12198_12199_reset_LC_19_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58153),
            .lcout(\comm_spi.n14617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57903),
            .ce(),
            .sr(N__58097));
    defparam \comm_spi.imiso_83_12208_12209_set_LC_19_10_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12208_12209_set_LC_19_10_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imiso_83_12208_12209_set_LC_19_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_12208_12209_set_LC_19_10_0  (
            .in0(N__56563),
            .in1(N__55412),
            .in2(_gnd_net_),
            .in3(N__55465),
            .lcout(\comm_spi.n14626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12208_12209_setC_net ),
            .ce(),
            .sr(N__56549));
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_19_10_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_19_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_105_2_lut_LC_19_10_1  (
            .in0(_gnd_net_),
            .in1(N__55152),
            .in2(_gnd_net_),
            .in3(N__56836),
            .lcout(\comm_spi.data_tx_7__N_790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_19_10_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_19_10_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_97_2_lut_LC_19_10_2  (
            .in0(N__55153),
            .in1(_gnd_net_),
            .in2(N__56853),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_19_10_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_19_10_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_87_2_lut_LC_19_10_6  (
            .in0(N__56837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55123),
            .lcout(\comm_spi.DOUT_7__N_748 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_19_10_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_19_10_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_19_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_88_2_lut_LC_19_10_7  (
            .in0(_gnd_net_),
            .in1(N__58154),
            .in2(_gnd_net_),
            .in3(N__56835),
            .lcout(\comm_spi.imosi_N_753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i2_12220_12221_reset_LC_19_11_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12220_12221_reset_LC_19_11_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i2_12220_12221_reset_LC_19_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12220_12221_reset_LC_19_11_0  (
            .in0(N__55070),
            .in1(N__55043),
            .in2(_gnd_net_),
            .in3(N__56459),
            .lcout(\comm_spi.n14639 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57012),
            .ce(),
            .sr(N__55082));
    defparam \comm_spi.data_tx_i2_12220_12221_set_LC_19_12_5 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12220_12221_set_LC_19_12_5 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i2_12220_12221_set_LC_19_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12220_12221_set_LC_19_12_5  (
            .in0(N__55069),
            .in1(N__55039),
            .in2(_gnd_net_),
            .in3(N__56455),
            .lcout(\comm_spi.n14638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57017),
            .ce(),
            .sr(N__55052));
    defparam \comm_spi.data_tx_i1_12216_12217_set_LC_19_13_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12216_12217_set_LC_19_13_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i1_12216_12217_set_LC_19_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12216_12217_set_LC_19_13_0  (
            .in0(N__56396),
            .in1(N__58085),
            .in2(_gnd_net_),
            .in3(N__57080),
            .lcout(\comm_spi.n14634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56917),
            .ce(),
            .sr(N__54992));
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_19_13_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_19_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_98_2_lut_LC_19_13_2  (
            .in0(N__55028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56841),
            .lcout(\comm_spi.data_tx_7__N_773 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12194_12195_set_LC_19_14_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12194_12195_set_LC_19_14_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.iclk_40_12194_12195_set_LC_19_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12194_12195_set_LC_19_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58041),
            .lcout(\comm_spi.n14612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57961),
            .ce(),
            .sr(N__56408));
    defparam \comm_spi.data_tx_i3_12224_12225_reset_LC_19_15_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12224_12225_reset_LC_19_15_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i3_12224_12225_reset_LC_19_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12224_12225_reset_LC_19_15_0  (
            .in0(N__55393),
            .in1(N__55366),
            .in2(_gnd_net_),
            .in3(N__55339),
            .lcout(\comm_spi.n14643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56918),
            .ce(),
            .sr(N__55325));
    defparam \comm_spi.i19214_4_lut_3_lut_LC_19_16_0 .C_ON=1'b0;
    defparam \comm_spi.i19214_4_lut_3_lut_LC_19_16_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19214_4_lut_3_lut_LC_19_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19214_4_lut_3_lut_LC_19_16_0  (
            .in0(N__55218),
            .in1(N__55319),
            .in2(_gnd_net_),
            .in3(N__56749),
            .lcout(\comm_spi.n22679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_19_16_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_19_16_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_19_16_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_103_2_lut_LC_19_16_2  (
            .in0(_gnd_net_),
            .in1(N__55280),
            .in2(_gnd_net_),
            .in3(N__56747),
            .lcout(\comm_spi.data_tx_7__N_784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_19_16_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_19_16_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_19_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_93_2_lut_LC_19_16_4  (
            .in0(_gnd_net_),
            .in1(N__55511),
            .in2(_gnd_net_),
            .in3(N__56748),
            .lcout(\comm_spi.data_tx_7__N_768 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_19_16_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_19_16_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_19_16_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_102_2_lut_LC_19_16_5  (
            .in0(N__56746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55246),
            .lcout(\comm_spi.data_tx_7__N_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19224_4_lut_3_lut_LC_19_16_6 .C_ON=1'b0;
    defparam \comm_spi.i19224_4_lut_3_lut_LC_19_16_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19224_4_lut_3_lut_LC_19_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19224_4_lut_3_lut_LC_19_16_6  (
            .in0(N__55247),
            .in1(N__55653),
            .in2(_gnd_net_),
            .in3(N__56750),
            .lcout(\comm_spi.n22673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i4_12228_12229_reset_LC_19_17_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12228_12229_reset_LC_19_17_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i4_12228_12229_reset_LC_19_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12228_12229_reset_LC_19_17_0  (
            .in0(N__55219),
            .in1(N__55202),
            .in2(_gnd_net_),
            .in3(N__55186),
            .lcout(\comm_spi.n14647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56997),
            .ce(),
            .sr(N__55172));
    defparam \comm_spi.data_tx_i5_12232_12233_reset_LC_19_18_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12232_12233_reset_LC_19_18_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i5_12232_12233_reset_LC_19_18_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12232_12233_reset_LC_19_18_0  (
            .in0(N__58237),
            .in1(N__58207),
            .in2(_gnd_net_),
            .in3(N__58192),
            .lcout(\comm_spi.n14651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57016),
            .ce(),
            .sr(N__55604));
    defparam i18943_2_lut_LC_20_2_0.C_ON=1'b0;
    defparam i18943_2_lut_LC_20_2_0.SEQ_MODE=4'b0000;
    defparam i18943_2_lut_LC_20_2_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18943_2_lut_LC_20_2_0 (
            .in0(_gnd_net_),
            .in1(N__55592),
            .in2(_gnd_net_),
            .in3(N__56377),
            .lcout(n21204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12204_3_lut_LC_20_6_6 .C_ON=1'b0;
    defparam \comm_spi.i12204_3_lut_LC_20_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12204_3_lut_LC_20_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i12204_3_lut_LC_20_6_6  (
            .in0(N__55478),
            .in1(N__55544),
            .in2(_gnd_net_),
            .in3(N__55520),
            .lcout(ICE_SPI_MISO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.MISO_48_12202_12203_reset_LC_20_7_1 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12202_12203_reset_LC_20_7_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.MISO_48_12202_12203_reset_LC_20_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.MISO_48_12202_12203_reset_LC_20_7_1  (
            .in0(N__55538),
            .in1(N__55427),
            .in2(_gnd_net_),
            .in3(N__55477),
            .lcout(\comm_spi.n14621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12202_12203_resetC_net ),
            .ce(),
            .sr(N__56487));
    defparam \comm_spi.MISO_48_12202_12203_set_LC_20_8_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12202_12203_set_LC_20_8_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.MISO_48_12202_12203_set_LC_20_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.MISO_48_12202_12203_set_LC_20_8_0  (
            .in0(N__55423),
            .in1(N__55534),
            .in2(_gnd_net_),
            .in3(N__55469),
            .lcout(\comm_spi.n14620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12202_12203_setC_net ),
            .ce(),
            .sr(N__56535));
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_20_8_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_20_8_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_91_2_lut_LC_20_8_2  (
            .in0(N__58030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56844),
            .lcout(\comm_spi.iclk_N_764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19229_4_lut_3_lut_LC_20_8_4 .C_ON=1'b0;
    defparam \comm_spi.i19229_4_lut_3_lut_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19229_4_lut_3_lut_LC_20_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19229_4_lut_3_lut_LC_20_8_4  (
            .in0(N__56577),
            .in1(N__55497),
            .in2(_gnd_net_),
            .in3(N__56845),
            .lcout(\comm_spi.n22661 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imiso_83_12208_12209_reset_LC_20_9_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12208_12209_reset_LC_20_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imiso_83_12208_12209_reset_LC_20_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_12208_12209_reset_LC_20_9_0  (
            .in0(N__56564),
            .in1(N__55411),
            .in2(_gnd_net_),
            .in3(N__55476),
            .lcout(\comm_spi.n14627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12208_12209_resetC_net ),
            .ce(),
            .sr(N__56488));
    defparam \comm_spi.data_tx_i7_12205_12206_reset_LC_20_10_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12205_12206_reset_LC_20_10_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i7_12205_12206_reset_LC_20_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12205_12206_reset_LC_20_10_0  (
            .in0(N__56584),
            .in1(N__55619),
            .in2(_gnd_net_),
            .in3(N__55685),
            .lcout(\comm_spi.n14624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56983),
            .ce(),
            .sr(N__56489));
    defparam \comm_spi.data_tx_i7_12205_12206_set_LC_20_11_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12205_12206_set_LC_20_11_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i7_12205_12206_set_LC_20_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12205_12206_set_LC_20_11_0  (
            .in0(N__56585),
            .in1(N__55618),
            .in2(_gnd_net_),
            .in3(N__55684),
            .lcout(\comm_spi.n14623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56991),
            .ce(),
            .sr(N__56542));
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_20_12_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_20_12_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_20_12_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_100_2_lut_LC_20_12_7  (
            .in0(_gnd_net_),
            .in1(N__56513),
            .in2(_gnd_net_),
            .in3(N__56810),
            .lcout(\comm_spi.data_tx_7__N_775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_12216_12217_reset_LC_20_13_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12216_12217_reset_LC_20_13_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i1_12216_12217_reset_LC_20_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12216_12217_reset_LC_20_13_0  (
            .in0(N__56395),
            .in1(N__58084),
            .in2(_gnd_net_),
            .in3(N__57079),
            .lcout(\comm_spi.n14635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56910),
            .ce(),
            .sr(N__56444));
    defparam \comm_spi.i12196_3_lut_LC_20_14_0 .C_ON=1'b0;
    defparam \comm_spi.i12196_3_lut_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12196_3_lut_LC_20_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.i12196_3_lut_LC_20_14_0  (
            .in0(N__57995),
            .in1(N__56432),
            .in2(_gnd_net_),
            .in3(N__56414),
            .lcout(\comm_spi.iclk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_20_14_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_20_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_90_2_lut_LC_20_14_1  (
            .in0(_gnd_net_),
            .in1(N__58031),
            .in2(_gnd_net_),
            .in3(N__56832),
            .lcout(\comm_spi.iclk_N_763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19234_4_lut_3_lut_LC_20_14_3 .C_ON=1'b0;
    defparam \comm_spi.i19234_4_lut_3_lut_LC_20_14_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19234_4_lut_3_lut_LC_20_14_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19234_4_lut_3_lut_LC_20_14_3  (
            .in0(N__56632),
            .in1(N__56394),
            .in2(_gnd_net_),
            .in3(N__56833),
            .lcout(\comm_spi.n22688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19080_2_lut_LC_20_14_4.C_ON=1'b0;
    defparam i19080_2_lut_LC_20_14_4.SEQ_MODE=4'b0000;
    defparam i19080_2_lut_LC_20_14_4.LUT_INIT=16'b0100010001000100;
    LogicCell40 i19080_2_lut_LC_20_14_4 (
            .in0(N__56367),
            .in1(N__55712),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n21320),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12236_12237_reset_LC_20_15_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12236_12237_reset_LC_20_15_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i6_12236_12237_reset_LC_20_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12236_12237_reset_LC_20_15_0  (
            .in0(N__55655),
            .in1(N__58181),
            .in2(_gnd_net_),
            .in3(N__55637),
            .lcout(\comm_spi.n14655 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56911),
            .ce(),
            .sr(N__55670));
    defparam \comm_spi.data_tx_i6_12236_12237_set_LC_20_16_5 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12236_12237_set_LC_20_16_5 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i6_12236_12237_set_LC_20_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12236_12237_set_LC_20_16_5  (
            .in0(N__55654),
            .in1(N__58177),
            .in2(_gnd_net_),
            .in3(N__55636),
            .lcout(\comm_spi.n14654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56987),
            .ce(),
            .sr(N__58247));
    defparam \comm_spi.data_tx_i5_12232_12233_set_LC_20_17_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12232_12233_set_LC_20_17_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i5_12232_12233_set_LC_20_17_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12232_12233_set_LC_20_17_0  (
            .in0(N__58241),
            .in1(N__58208),
            .in2(_gnd_net_),
            .in3(N__58193),
            .lcout(\comm_spi.n14650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56996),
            .ce(),
            .sr(N__58166));
    defparam CONSTANT_ONE_LUT4_LC_22_3_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_3_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_3_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_22_9_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_22_9_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_22_9_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_89_2_lut_LC_22_9_0  (
            .in0(N__58128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56842),
            .lcout(\comm_spi.imosi_N_754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_22_9_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_22_9_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_22_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_99_2_lut_LC_22_9_6  (
            .in0(_gnd_net_),
            .in1(N__56628),
            .in2(_gnd_net_),
            .in3(N__56843),
            .lcout(\comm_spi.data_tx_7__N_774 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12190_12191_set_LC_22_10_7 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12190_12191_set_LC_22_10_7 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i0_12190_12191_set_LC_22_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_12190_12191_set_LC_22_10_7  (
            .in0(N__57186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57051),
            .ce(),
            .sr(N__58067));
    defparam \comm_spi.iclk_40_12194_12195_reset_LC_22_12_5 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12194_12195_reset_LC_22_12_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.iclk_40_12194_12195_reset_LC_22_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.iclk_40_12194_12195_reset_LC_22_12_5  (
            .in0(N__58054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57970),
            .ce(),
            .sr(N__57440));
    defparam \comm_spi.data_tx_i0_12190_12191_reset_LC_22_13_1 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12190_12191_reset_LC_22_13_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i0_12190_12191_reset_LC_22_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_12190_12191_reset_LC_22_13_1  (
            .in0(N__57237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__57040),
            .ce(),
            .sr(N__56597));
    defparam \comm_spi.RESET_I_0_2_lut_LC_22_14_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_2_lut_LC_22_14_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_2_lut_LC_22_14_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_2_lut_LC_22_14_7  (
            .in0(N__56834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56633),
            .lcout(\comm_spi.data_tx_7__N_796 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // zim
